
module pri_encoder( clk );
  input wire clk;

  integer ctr = 0;

  reg [6:0] state = 0;
  reg [6:0] diff_shif;
  reg [54:0] diff = 0;

  //integer i, width;
  //reg[55:0] part;
  
  
  always @(posedge clk) begin
    state <= (state + 1) % 56;
    ctr <= ctr + 1;

    if (ctr >= 1000) $finish();


    casex(state)  
      0: diff <= 55'b1111111111111111111111111111111111111111111111111111111; // : diff_shift <=  0;
      1: diff <= 55'b0111111111111111111111111111111111111111111111111111111; // : diff_shift <=  1;
      2: diff <= 55'b0011111111111111111111111111111111111111111111111111111; // : diff_shift <=  2;
      3: diff <= 55'b0001111111111111111111111111111111111111111111111111111; // : diff_shift <=  3;
      4: diff <= 55'b0000111111111111111111111111111111111111111111111111111; // : diff_shift <=  4;
      5: diff <= 55'b0000011111111111111111111111111111111111111111111111111; // : diff_shift <=  5;
      6: diff <= 55'b0000001111111111111111111111111111111111111111111111111; // : diff_shift <=  6;
      7: diff <= 55'b0000000111111111111111111111111111111111111111111111111; // : diff_shift <=  7;
      8: diff <= 55'b0000000011111111111111111111111111111111111111111111111; // : diff_shift <=  8;
      9: diff <= 55'b0000000001111111111111111111111111111111111111111111111; // : diff_shift <=  9;
      10: diff <= 55'b0000000000111111111111111111111111111111111111111111111; // : diff_shift <=  10;
      11: diff <= 55'b0000000000011111111111111111111111111111111111111111111; // : diff_shift <=  11;
      12: diff <= 55'b0000000000001111111111111111111111111111111111111111111; // : diff_shift <=  12;
      13: diff <= 55'b0000000000000111111111111111111111111111111111111111111; // : diff_shift <=  13;
      14: diff <= 55'b0000000000000011111111111111111111111111111111111111111; // : diff_shift <=  14;
      15: diff <= 55'b0000000000000001111111111111111111111111111111111111111; // : diff_shift <=  15;
      16: diff <= 55'b0000000000000000111111111111111111111111111111111111111; // : diff_shift <=  16;
      17: diff <= 55'b0000000000000000011111111111111111111111111111111111111; // : diff_shift <=  17;
      18: diff <= 55'b0000000000000000001111111111111111111111111111111111111; // : diff_shift <=  18;
      19: diff <= 55'b0000000000000000000111111111111111111111111111111111111; // : diff_shift <=  19;
      20: diff <= 55'b0000000000000000000011111111111111111111111111111111111; // : diff_shift <=  20;
      21: diff <= 55'b0000000000000000000001111111111111111111111111111111111; // : diff_shift <=  21;
      22: diff <= 55'b0000000000000000000000111111111111111111111111111111111; // : diff_shift <=  22;
      23: diff <= 55'b0000000000000000000000011111111111111111111111111111111; // : diff_shift <=  23;
      24: diff <= 55'b0000000000000000000000001111111111111111111111111111111; // : diff_shift <=  24;
      25: diff <= 55'b0000000000000000000000000111111111111111111111111111111; // : diff_shift <=  25;
      26: diff <= 55'b0000000000000000000000000011111111111111111111111111111; // : diff_shift <=  26;
      27: diff <= 55'b0000000000000000000000000001111111111111111111111111111; // : diff_shift <=  27;
      28: diff <= 55'b0000000000000000000000000000111111111111111111111111111; // : diff_shift <=  28;
      29: diff <= 55'b0000000000000000000000000000011111111111111111111111111; // : diff_shift <=  29;
      30: diff <= 55'b0000000000000000000000000000001111111111111111111111111; // : diff_shift <=  30;
      31: diff <= 55'b0000000000000000000000000000000111111111111111111111111; // : diff_shift <=  31;
      32: diff <= 55'b0000000000000000000000000000000011111111111111111111111; // : diff_shift <=  32;
      33: diff <= 55'b0000000000000000000000000000000001111111111111111111111; // : diff_shift <=  33;
      34: diff <= 55'b0000000000000000000000000000000000111111111111111111111; // : diff_shift <=  34;
      35: diff <= 55'b0000000000000000000000000000000000011111111111111111111; // : diff_shift <=  35;
      36: diff <= 55'b0000000000000000000000000000000000001111111111111111111; // : diff_shift <=  36;
      37: diff <= 55'b0000000000000000000000000000000000000111111111111111111; // : diff_shift <=  37;
      38: diff <= 55'b0000000000000000000000000000000000000011111111111111111; // : diff_shift <=  38;
      39: diff <= 55'b0000000000000000000000000000000000000001111111111111111; // : diff_shift <=  39;
      40: diff <= 55'b0000000000000000000000000000000000000000111111111111111; // : diff_shift <=  40;
      41: diff <= 55'b0000000000000000000000000000000000000000011111111111111; // : diff_shift <=  41;
      42: diff <= 55'b0000000000000000000000000000000000000000001111111111111; // : diff_shift <=  42;
      43: diff <= 55'b0000000000000000000000000000000000000000000111111111111; // : diff_shift <=  43;
      44: diff <= 55'b0000000000000000000000000000000000000000000011111111111; // : diff_shift <=  44;
      45: diff <= 55'b0000000000000000000000000000000000000000000001111111111; // : diff_shift <=  45;
      46: diff <= 55'b0000000000000000000000000000000000000000000000111111111; // : diff_shift <=  46;
      47: diff <= 55'b0000000000000000000000000000000000000000000000011111111; // : diff_shift <=  47;
      48: diff <= 55'b0000000000000000000000000000000000000000000000001111111; // : diff_shift <=  48;
      49: diff <= 55'b0000000000000000000000000000000000000000000000000111111; // : diff_shift <=  49;
      50: diff <= 55'b0000000000000000000000000000000000000000000000000011111; // : diff_shift <=  50;
      51: diff <= 55'b0000000000000000000000000000000000000000000000000001111; // : diff_shift <=  51;
      52: diff <= 55'b0000000000000000000000000000000000000000000000000000111; // : diff_shift <=  52;
      53: diff <= 55'b0000000000000000000000000000000000000000000000000000011; // : diff_shift <=  53;
      54: diff <= 55'b0000000000000000000000000000000000000000000000000000001; // : diff_shift <=  54;
      55: diff <= 55'b0000000000000000000000000000000000000000000000000000000; // : diff_shift <=  55;
    endcase    

    $display("state: %d, diff: %d", state, diff);
    $display("msb: %d", msb);

  end // always @ (posedge clk)


  parameter WIDTH = 56;
  parameter WIDTH_LOG = 6;

  wire [WIDTH_LOG - 1:0] msb;
  
  wire [(WIDTH_LOG * WIDTH) - 1:0] ors;

  assign ors[WIDTH_LOG * WIDTH - 1:(WIDTH_LOG - 1) * WIDTH ] = diff;

  genvar w;

  for (w = WIDTH_LOG - 1; w >= 0; w = w - 1) begin
    assign msb[w] = |ors[w * WIDTH + 2 * (1 << w) - 1: w * WIDTH + (1 << w)];
    if (w > 0) begin
      assign ors[(w - 1) * WIDTH + (1 << w) - 1:(w - 1) * WIDTH] = msb[w] ? ors[w*WIDTH + 2*(1 << w) - 1:w*WIDTH + (1 << w)] : ors[w*WIDTH + (1 << w) - 1:w*WIDTH];
    end
  end

endmodule


//pri_encoder pe(clock.val);
