include fpu_pri_encoder.v;

module pri_encoder( clk );
  input wire clk;

  integer ctr = 0;

  reg [6:0] state = 0;
  reg [6:0] diff_shift;
  reg [105:0] diff = 0;
  
  always @(posedge clk) begin
    state <= (state + 1) % 56;
    ctr <= ctr + 1;

    if (ctr >= 57) $finish();


    case(state)  // uses prev state (before this cycle)
      //1: diff <= 55'b1000000000000000000000000000000000000000000000000000000;
      //0: diff <= 55'b0000000000000000000000000000000000000000000000000000001;
      //1: diff <= 55'b0000000000000000000000000000000000000000000000000000010;
      //2: diff <= 55'b0000000000000000000000000000000000000000000000000100000;
      //3: diff <= 55'b0000111111111111111111111111111111111111111111111111111;
      //0: diff <= 106'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      //default: diff <= 55'b0000000000000000000000000000000000000000000000000001000;
      
      0: diff <= 55'b1111111111111111111111111111111111111111111111111111111;
      1: diff <= 55'b0111111111111111111111111111111111111111111111111111111; 
      2: diff <= 55'b0011111111111111111111111111111111111111111111111111111; 
      3: diff <= 55'b0001111111111111111111111111111111111111111111111111111; 
      4: diff <= 55'b0000111111111111111111111111111111111111111111111111111; 
      5: diff <= 55'b0000011111111111111111111111111111111111111111111111111; 
      6: diff <= 55'b0000001111111111111111111111111111111111111111111111111; 
      7: diff <= 55'b0000000111111111111111111111111111111111111111111111111; 
      8: diff <= 55'b0000000011111111111111111111111111111111111111111111111; 
      9: diff <= 55'b0000000001111111111111111111111111111111111111111111111; 
      10: diff <= 55'b0000000000111111111111111111111111111111111111111111111;
      11: diff <= 55'b0000000000011111111111111111111111111111111111111111111;
      12: diff <= 55'b0000000000001111111111111111111111111111111111111111111;
      13: diff <= 55'b0000000000000111111111111111111111111111111111111111111;
      14: diff <= 55'b0000000000000011111111111111111111111111111111111111111;
      15: diff <= 55'b0000000000000001111111111111111111111111111111111111111;
      16: diff <= 55'b0000000000000000111111111111111111111111111111111111111;
      17: diff <= 55'b0000000000000000011111111111111111111111111111111111111;
      18: diff <= 55'b0000000000000000001111111111111111111111111111111111111;
      19: diff <= 55'b0000000000000000000111111111111111111111111111111111111;
      20: diff <= 55'b0000000000000000000011111111111111111111111111111111111;
      21: diff <= 55'b0000000000000000000001111111111111111111111111111111111;
      22: diff <= 55'b0000000000000000000000111111111111111111111111111111111;
      23: diff <= 55'b0000000000000000000000011111111111111111111111111111111;
      24: diff <= 55'b0000000000000000000000001111111111111111111111111111111;
      25: diff <= 55'b0000000000000000000000000111111111111111111111111111111;
      26: diff <= 55'b0000000000000000000000000011111111111111111111111111111;
      27: diff <= 55'b0000000000000000000000000001111111111111111111111111111;
      28: diff <= 55'b0000000000000000000000000000111111111111111111111111111;
      29: diff <= 55'b0000000000000000000000000000011111111111111111111111111;
      30: diff <= 55'b0000000000000000000000000000001111111111111111111111111;
      31: diff <= 55'b0000000000000000000000000000000111111111111111111111111;
      32: diff <= 55'b0000000000000000000000000000000011111111111111111111111;
      33: diff <= 55'b0000000000000000000000000000000001111111111111111111111;
      34: diff <= 55'b0000000000000000000000000000000000111111111111111111111;
      35: diff <= 55'b0000000000000000000000000000000000011111111111111111111;
      36: diff <= 55'b0000000000000000000000000000000000001111111111111111111;
      37: diff <= 55'b0000000000000000000000000000000000000111111111111111111;
      38: diff <= 55'b0000000000000000000000000000000000000011111111111111111;
      39: diff <= 55'b0000000000000000000000000000000000000001111111111111111;
      40: diff <= 55'b0000000000000000000000000000000000000000111111111111111;
      41: diff <= 55'b0000000000000000000000000000000000000000011111111111111;
      42: diff <= 55'b0000000000000000000000000000000000000000001111111111111;
      43: diff <= 55'b0000000000000000000000000000000000000000000111111111111;
      44: diff <= 55'b0000000000000000000000000000000000000000000011111111111;
      45: diff <= 55'b0000000000000000000000000000000000000000000001111111111;
      46: diff <= 55'b0000000000000000000000000000000000000000000000111111111;
      47: diff <= 55'b0000000000000000000000000000000000000000000000011111111;
      48: diff <= 55'b0000000000000000000000000000000000000000000000001111111;
      49: diff <= 55'b0000000000000000000000000000000000000000000000000111111;
      50: diff <= 55'b0000000000000000000000000000000000000000000000000011111;
      51: diff <= 55'b0000000000000000000000000000000000000000000000000001111;
      52: diff <= 55'b0000000000000000000000000000000000000000000000000000111;
      53: diff <= 55'b0000000000000000000000000000000000000000000000000000011;
      54: diff <= 55'b0000000000000000000000000000000000000000000000000000001;
      55: diff <= 55'b0000000000000000000000000000000000000000000000000000000;
 
    endcase    

    $display("state: %d, diff: %d, msb: %d, diff_shift: %d", state, diff, msb, diff_shift);
    

  end // always @ (posedge clk)

  always @(*) begin
    diff_shift <= msb ? (54 - msb) : (diff ? 54 : 55);
  end

  fpu_pri_encoder pri_en(diff, msb);



  //parameter WIDTH = 106;
  parameter WIDTH_LOG = 7;
  //
  wire [WIDTH_LOG - 1:0] msb;
  //
  //genvar i;
  //
  //for (i = 0; i < WIDTH_LOG; i = i + 1) begin : ORS
  //  wire [WIDTH - 1:0] oi;
  //  wire msbi;
  //
  //  if (i == 0)
  //    assign oi = diff;
  //  else
  //    assign oi[(1 << ((WIDTH_LOG - 1 - i) + 1)) - 1:0] = ORS[i - 1].msbi ? ORS[i - 1].oi[2 * (1 << ((WIDTH_LOG - 1 - i) + 1)) - 1:(1 << ((WIDTH_LOG - 1 - i) + 1))] : ORS[i - 1].oi[(1 << ((WIDTH_LOG - 1 - i) + 1)) - 1 : 0];
  //
  //  assign msbi = |oi[2 * (1 << (WIDTH_LOG - 1 - i)) - 1: (1 << (WIDTH_LOG - 1 - i))];
  //  assign msb[WIDTH_LOG - 1 - i] = |oi[2 * (1 << (WIDTH_LOG - 1 - i)) - 1: (1 << (WIDTH_LOG - 1 - i))];
  //  
  //end

endmodule // pri_encoder



pri_encoder pe(clock.val);
