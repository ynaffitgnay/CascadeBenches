//---------------------------------------------------------------------------------------
//  Project:  ADPCM Encoder / Decoder
//
//  Filename:  tb_ima_adpcm.v      (April 26, 2010 )
//
//  Author(s):  Moti Litochevski
//
//  Description:
//    This file implements the ADPCM encoder & decoder test bench. The input samples
//    to be encoded are read from a binary input file. The encoder stream output and
//    decoded samples are also compared with binary files generated by the Scilab
//    simulation.
//
//---------------------------------------------------------------------------------------
//
//  To Do:
//  -
//
//---------------------------------------------------------------------------------------
//
//  Copyright (C) 2010 Moti Litochevski
//
//  This source file may be used and distributed without restriction provided that this
//  copyright statement is not removed from the file and that any derivative work
//  contains the original copyright notice and the associated disclaimer.
//
//  THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES,
//  INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND
//  FITNESS FOR A PARTICULAR PURPOSE.
//
//---------------------------------------------------------------------------------------
// Refactored to run on Cascade in April 2019 by Tiffany Yang

`include "ima_adpcm_enc.v"
`include "ima_adpcm_dec.v"

module test(clk);
  parameter BUFFER_BYTES = 32;

  // Truncated for development
  parameter TOTAL_IN_BYTES = 87040;
  parameter TOTAL_ENC_BYTES = 43520;
  parameter TOTAL_DEC_BYTES = 87040;

  parameter MAIN0 = 0;
  parameter MAIN1 = 1;
  parameter MAIN2 = 2;

  parameter IN0 = 0;
  parameter IN1 = 1;
  parameter IN2 = 2;
  parameter IN3 = 3;
  parameter IN4 = 4;
  parameter IN5 = 5;

  parameter ENC0 = 0;
  parameter ENC1 = 1;
  parameter ENC2 = 2;
  parameter ENC3 = 3;
  parameter ENC4 = 4;

  parameter DEC0 = 0;
  parameter DEC1 = 1;
  parameter DEC2 = 2;
  parameter DEC3 = 3;
  parameter DEC4 = 4;

  parameter TESTS_TO_RUN = 1;

  
  input wire clk;

  //---------------------------------------------------------------------------------------
  // internal signal
  reg rst;        // global reset
  reg [15:0] inSamp;    // encoder input sample
  reg inValid;      // encoder input valid flag
  wire inReady;      // encoder input ready indication
  wire [3:0] encPcm;    // encoder encoded output value
  wire encValid;      // encoder output valid flag
  wire decReady;     // decoder ready for input indication
  wire [15:0] decSamp;  // decoder output sample value
  wire decValid;      // decoder output valid flag
  integer sampCount, encCount, decCount;

  reg [7:0] intmp, enctmp, dectmp;
  reg [3:0] encExpVal;
  reg [15:0] decExpVal;
  reg [31:0] dispCount;

  reg inDone, encDone, decDone;

  reg[31:0] testCount;

  reg[7:0] inReg, decReg;

  // Variables to read file input into before copying to in-mem buffer
  reg[(BUFFER_BYTES << 3) - 1:0] inVal;
  reg[(BUFFER_BYTES << 3) - 1:0] encVal;
  reg[(BUFFER_BYTES << 3) - 1:0] decVal;

  reg[15:0] inIdx, encIdx, decIdx;

  // Buffers to hold file content
  reg[(BUFFER_BYTES << 3) - 1:0] inBuf [(TOTAL_IN_BYTES / BUFFER_BYTES) - 1:0];
  reg[(BUFFER_BYTES << 3) - 1:0] encBuf [(TOTAL_ENC_BYTES / BUFFER_BYTES) - 1:0];
  reg[(BUFFER_BYTES << 3) - 1:0] decBuf [(TOTAL_DEC_BYTES / BUFFER_BYTES) - 1:0];
  reg[31:0] inBytesRead, encBytesRead, decBytesRead;


  reg[3:0] mainState;
  reg[3:0] inState;
  reg[3:0] encState;
  reg[3:0] decState;

  reg[31:0] mCtr;
  reg[31:0] iCtr;
  reg[31:0] eCtr;
  reg[31:0] dCtr;

  initial begin
    $display("Initializing");

    testCount = 0;

    mCtr = 0;
    mainState = 0;

    iCtr = 0;
    inState = 0;

    eCtr = 0;
    encState = 0;

    dCtr = 0;
    decState = 0;

    
    inBuf[0] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[1] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[2] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[3] = 256'h0000000000000000000000000000000000000000000000000000000000000000;    
    inBuf[4] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[5] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[6] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[7] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[8] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[9] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[10] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[11] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[12] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[13] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[14] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[15] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[16] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[17] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[18] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[19] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[20] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[21] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[22] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[23] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[24] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[25] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[26] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[27] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[28] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[29] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[30] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[31] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[32] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[33] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[34] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[35] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[36] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[37] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[38] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[39] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[40] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[41] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[42] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[43] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[44] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[45] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[46] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[47] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[48] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[49] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[50] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[51] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[52] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[53] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[54] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[55] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[56] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[57] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[58] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[59] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[60] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[61] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[62] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[63] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[64] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[65] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[66] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[67] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[68] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[69] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[70] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[71] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[72] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[73] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[74] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[75] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[76] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[77] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[78] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[79] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[80] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[81] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[82] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[83] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[84] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[85] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[86] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[87] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[88] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[89] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[90] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[91] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[92] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[93] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[94] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[95] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[96] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[97] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[98] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[99] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[100] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[101] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[102] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[103] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[104] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[105] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[106] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[107] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[108] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[109] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[110] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[111] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[112] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[113] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[114] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[115] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[116] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[117] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[118] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[119] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[120] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[121] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[122] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[123] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[124] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[125] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[126] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[127] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[128] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[129] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[130] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[131] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[132] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[133] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[134] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[135] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[136] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[137] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[138] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[139] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[140] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[141] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[142] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[143] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[144] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[145] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[146] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[147] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[148] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[149] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[150] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[151] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[152] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[153] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[154] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[155] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[156] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[157] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[158] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[159] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[160] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[161] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[162] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[163] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[164] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[165] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[166] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[167] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[168] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[169] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[170] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[171] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[172] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[173] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[174] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[175] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[176] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[177] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[178] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[179] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[180] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[181] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[182] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[183] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[184] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[185] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[186] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[187] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[188] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[189] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[190] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[191] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[192] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[193] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[194] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[195] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[196] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[197] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[198] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[199] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[200] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[201] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[202] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[203] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[204] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[205] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[206] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[207] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[208] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[209] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[210] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[211] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[212] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[213] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[214] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[215] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[216] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[217] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[218] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[219] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[220] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[221] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[222] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[223] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[224] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[225] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[226] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[227] = 256'h000000000000ffff000000000000000000000000000000000000000000000000;
    inBuf[228] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[229] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[230] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[231] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[232] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[233] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[234] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[235] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[236] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[237] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[238] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[239] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[240] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[241] = 256'h0000000000000000ffff00000000000000000000000000000000000000000000;
    inBuf[242] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[243] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[244] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[245] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[246] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[247] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[248] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[249] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[250] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[251] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[252] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[253] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[254] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[255] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[256] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[257] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[258] = 256'h0000000000000000000000000000010001000000000000000000ffff00000000;
    inBuf[259] = 256'h0000000000000000ffff00000000000000000000ffffffff0000000000000000;
    inBuf[260] = 256'h00000000000000000000ffff000000000000000000000000000000000000ffff;
    inBuf[261] = 256'h0000000000000000000000000000ffff00000000ffffffff0000000000000000;
    inBuf[262] = 256'h0000ffff00000000000000000000000000000000010000000000000000000000;
    inBuf[263] = 256'h0000000000000100010000000000010000000000000000000000000001000000;
    inBuf[264] = 256'h0000000000000000000000000000000000000000ffffffff0000010000000000;
    inBuf[265] = 256'h00000000ffff0000010001000000000000000000ffff00000000000000000000;
    inBuf[266] = 256'h00000000000000000000000000000000ffff0000000000000000000000000000;
    inBuf[267] = 256'h00000000ffff0000000000000000010000000000000000000000000000000000;
    inBuf[268] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[269] = 256'h000000000000000000000000ffffffff000001000100ffffffff000000000000;
    inBuf[270] = 256'h000000000000ffff0000000000000000010000000000ffff0000010001000000;
    inBuf[271] = 256'h0000000000000000000000000000000001000000000000000000000000000100;
    inBuf[272] = 256'h0000ffff00000000ffff00000000000000000000000000000000000000000000;
    inBuf[273] = 256'h0000ffff0000010001000000000000000000ffff0000010001000000ffff0100;
    inBuf[274] = 256'h0100000000000000000000000000010000000000000000000000000000000000;
    inBuf[275] = 256'h0000000001000000000000000000000000000000000000000100010000000000;
    inBuf[276] = 256'h00000000010000000000000000000000000000000000000000000000ffff0000;
    inBuf[277] = 256'h00000000000000000000ffffffff000001000000000000000000000000000000;
    inBuf[278] = 256'h0000000000000000ffff00000100000000000000000000000100010000000000;
    inBuf[279] = 256'h00000000000000000000000001000100ffffffff00000000ffffffff00000000;
    inBuf[280] = 256'h00000000000000000000ffff0000010000000000000000000000000000000000;
    inBuf[281] = 256'h0000000000000000010000000000000000000000000000000000000000000000;
    inBuf[282] = 256'h00000000000000000000ffff0000000000000000000000000000000000000000;
    inBuf[283] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[284] = 256'h00000000000000000000000000000000ffff0000000000000000000000000000;
    inBuf[285] = 256'h0000000000000000000000000000000000000000000001000100000000000000;
    inBuf[286] = 256'h00000000000000000000010000000000000001000000ffff0000000000000000;
    inBuf[287] = 256'h000000000000000000000000ffffffff00000000000000000000000000000000;
    inBuf[288] = 256'h0000000000000100010000000000000000000000000000000000000000000000;
    inBuf[289] = 256'h00000000000000000000ffff000000000000ffff000000000000ffff00000000;
    inBuf[290] = 256'h0000000000000000000000000000ffff0000010001000000ffff000000000000;
    inBuf[291] = 256'h00000000000001000000000000000000ffff000001000100000001000000ffff;
    inBuf[292] = 256'h00000000010000000000000000000000ffff0000000000000000000000000000;
    inBuf[293] = 256'h0000ffffffff00000000000000000000000000000000000000000000ffffffff;
    inBuf[294] = 256'h00000100000000000000000000000000ffffffff00000100000000000000ffff;
    inBuf[295] = 256'hffff000001000000000000000000000000000000000000000000000001000000;
    inBuf[296] = 256'h000000000000ffff000000000000000000000000000000000000000001000100;
    inBuf[297] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[298] = 256'hffff000000000000000001000100000000000000000000000000000000000100;
    inBuf[299] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[300] = 256'h000000000000000000000000ffffffff000001000000ffffffffffff00000000;
    inBuf[301] = 256'h0000000000000000000000000000000000000000000000000000000001000000;
    inBuf[302] = 256'h0000000000000000010000000000000000000000000000000000000000000000;
    inBuf[303] = 256'h000000000000ffffffff000000000000ffff0000000000000000000000000000;
    inBuf[304] = 256'h0000000000000000000000000000000000000000000000000100000000000000;
    inBuf[305] = 256'h0000ffff00000100010000000000000000000000000000000000000000000100;
    inBuf[306] = 256'h0100000000000000000000000000000000000000000000000000000000000000;
    inBuf[307] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[308] = 256'h000000000000010001000000ffff000000000000000000000000000000000000;
    inBuf[309] = 256'h0000000000000000000000000000000000000000000000000000000001000000;
    inBuf[310] = 256'h0000000000000000000000000000000000000100000000000000000000000000;
    inBuf[311] = 256'h00000000000000000000000000000000000000000000ffffffff00000000ffff;
    inBuf[312] = 256'hffff00000000000000000000000000000000ffff000000000000000000000100;
    inBuf[313] = 256'h010000000000000001000000000000000000000001000100000000000000ffff;
    inBuf[314] = 256'hffff000000000000000000000000000000000000000000000000000000000000;
    inBuf[315] = 256'h0000000000000000000000000000ffff00000000ffffffff010001000000ffff;
    inBuf[316] = 256'h000000000000000000000000000000000000000000000000000001000000ffff;
    inBuf[317] = 256'hffff000000000000010000000000ffffffff0000000000000000010000000000;
    inBuf[318] = 256'h000000000000000000000000000000000000000000000000000000000000ffff;
    inBuf[319] = 256'h0000000000000000010000000000000000000000000000000000000000000000;
    inBuf[320] = 256'h0000010000000000000000000000000000000000000000000000000000000000;
    inBuf[321] = 256'h000000000000010000000000000000000000000000000100000000000000ffff;
    inBuf[322] = 256'h00000000000000000000000000000000ffffffff0000ffff0000010000000000;
    inBuf[323] = 256'h00000000ffffffffffffffffffff000000000000000001000000ffff00000100;
    inBuf[324] = 256'hffffffff00000000000000000000000001000100ffffffff0000000000000000;
    inBuf[325] = 256'h01000000000000000000ffffffff00000000000001000100010000000000ffff;
    inBuf[326] = 256'h00000000ffff000000000000010000000000ffff000001000000000000000100;
    inBuf[327] = 256'h01000000ffff000001000100000000000000ffffffff00000000000000000000;
    inBuf[328] = 256'h000000000000000000000000000000000000ffff000001000000ffff00000000;
    inBuf[329] = 256'h0000000001000000000000000000000000000100000000000000000000000000;
    inBuf[330] = 256'h00000000000000000100000000000000000000000000ffffffff000001000000;
    inBuf[331] = 256'h00000000ffffffff000000000000ffffffff0000000000000000000000000000;
    inBuf[332] = 256'h0000000000000100fffffffffffffefffbfffbff00000d0019001200f7ffe9ff;
    inBuf[333] = 256'hf8ff0000ecffdfffedfffcff02000f0019000a00f4ffeffff9ff03000b000f00;
    inBuf[334] = 256'h0c0009000a000c000f001a0027002e002a001600ffff0a002e002800f0ffd1ff;
    inBuf[335] = 256'he2ffedffe3fff8ff250032002200240033002d0015000600040009000e000700;
    inBuf[336] = 256'hf8fff2fff7fffcfff9ffe7ffcbffc3ffd5ffd5ffbeffceff0b0028001c002d00;
    inBuf[337] = 256'h48001900c1ffb6fff0ff0300d9ffb2ffaaffb4ffcaffe0ffe8ffeaffebffe2ff;
    inBuf[338] = 256'hdaffe4fff9ff140031002400e0ffb1ffcefff9ff0e0047008300580003002300;
    inBuf[339] = 256'h7600370091ff58ffaaff020025002a00190008000f0012000400fdfff0ffc4ff;
    inBuf[340] = 256'h9fff9aff8cff95ff00005900280007005b004400a2ffc0ff6000d1ff46ff2202;
    inBuf[341] = 256'h87078d0aec093e09120a4e0a6b093609bb099e094909b709220abd0949092909;
    inBuf[342] = 256'hb6080108ba079a072f070507590771072b072d075207ee064506eb05a5054605;
    inBuf[343] = 256'h5805f0056706770664063f0610062006680688068406a406cb06d20608079b07;
    inBuf[344] = 256'h4e080209bb092d0a270afa09ec09e209e609390ac50a4d0bc80b260c3b0c360c;
    inBuf[345] = 256'h5f0c790c3b0cea0bc30b880b3a0b450b9b0bc30bb60bba0ba90b540bfb0abe0a;
    inBuf[346] = 256'h640afb09c409a1095e092f0938092d09ee08b5087808ff0773072207ff06e906;
    inBuf[347] = 256'hf6061b072b07340754076d076b0776078c078207640767077d079407cf073a08;
    inBuf[348] = 256'ha108f8085d09bb09ee09090a1e0a1d0a0a0a0f0a3c0a800ad50a330b780b960b;
    inBuf[349] = 256'h9a0b810b430b030be30ad70ad00ad50adf0ad00aa50a740a420a0b0ada09b809;
    inBuf[350] = 256'h920963093a091409e708bc0894085e081008bc076e07330723073e0761077007;
    inBuf[351] = 256'h6c0757072907f006cd06ca06dc06ff062d075607720786079807a807bd07d707;
    inBuf[352] = 256'hed07fe070f081f082f08410854085e08620864086308630870088b089f089e08;
    inBuf[353] = 256'h86084c08eb0778071607d706b806af06ad069b066f062606c4055405ee049b04;
    inBuf[354] = 256'h5f043b042b04220413040204f403e203cc03b6039c037403470326031c032b03;
    inBuf[355] = 256'h50038103ab03be03b903a6039803a103c603ff0344048704b804d204e004ec04;
    inBuf[356] = 256'h09053c057605ae05d805ed05ee05e305d305c105ad058e0559051005b8046404;
    inBuf[357] = 256'h2104f303d103ac036e03100398021602a10146010901df00ba008d0052000e00;
    inBuf[358] = 256'hc5ff81ff45ff0dffd5fe9efe6afe3ffe20fe0efe04fef8fddffdb6fd86fd58fd;
    inBuf[359] = 256'h3bfd39fd59fd95fde0fd2cfe73feaffeddfe05ff32ff6bffb0ffffff51009e00;
    inBuf[360] = 256'hd700f600ff00f800e700d400c600bd00b2009b00760048001100daffabff87ff;
    inBuf[361] = 256'h69ff4dff2cff0affecfecdfeaefe88fe4ffefefd9bfd32fdd8fc98fc6dfc4efc;
    inBuf[362] = 256'h2dfcf9fbb2fb65fb1cfbe1fab6fa90fa69fa3efa0cfae0f9c8f9c4f9dbf908fa;
    inBuf[363] = 256'h39fa68fa8cfa9dfa9efa9afa94fa9cfab9fae5fa22fb6efbb6fbf7fb29fc3efc;
    inBuf[364] = 256'h35fc12fcd9fba3fb81fb73fb7efb9afbacfbabfb94fb63fb2cfbf9facafaaffa;
    inBuf[365] = 256'ha6fa9dfa94fa86fa64fa30faf1f9abf973f954f946f94df95ff95cf93ff906f9;
    inBuf[366] = 256'hacf849f8eff7a9f791f7adf7e7f739f88df8bdf8c1f896f840f8e5f7a4f78cf7;
    inBuf[367] = 256'hb5f71bf897f815f978f9a0f998f96ef92ff900f9f4f802f933f97cf9c0f9fef9;
    inBuf[368] = 256'h2efa3bfa34fa1bfae6f9adf97df952f93df93cf932f920f9fbf8b1f85cf811f8;
    inBuf[369] = 256'hd3f7b7f7b7f7b2f7a3f77df72df7cff67bf62ef6fff5f3f5f6f50df62ff642f6;
    inBuf[370] = 256'h4df648f61cf6e0f5a8f573f560f57af5abf5f4f541f671f692f6a9f6a7f6a7f6;
    inBuf[371] = 256'hb7f6c6f6e7f61bf750f795f7e5f720f856f887f89bf8acf8c8f8e3f810f94bf9;
    inBuf[372] = 256'h74f992f99ef982f95bf93cf91af909f907f9f9f8e9f8daf8b6f896f87bf848f8;
    inBuf[373] = 256'h0cf8ccf779f737f715f701f708f71af70ef7f0f6c3f67ef645f625f608f6fcf5;
    inBuf[374] = 256'hfbf5e6f5cef5bef5a5f5a0f5b1f5bef5d7f5fbf512f630f65ef684f6b1f6e5f6;
    inBuf[375] = 256'h05f729f757f77ef7b8f709f84ff891f8ccf8e5f8f1f8f7f8e7f8ddf8dff8d6f8;
    inBuf[376] = 256'hddf8fcf81af945f978f991f99ef99ef981f96af966f95ff966f977f96ff958f9;
    inBuf[377] = 256'h36f9fbf8c7f8a3f875f850f830f8f8f7c2f799f771f762f769f767f767f769f7;
    inBuf[378] = 256'h5af759f773f793f7c6f703f82cf851f879f895f8bdf8f5f81ff947f96cf97bf9;
    inBuf[379] = 256'h91f9b9f9e1f916fa52fa74fa89fa96fa8ffa92faa5faaffabbfac6fabafab0fa;
    inBuf[380] = 256'hb5fac0fae3fa15fb33fb42fb43fb24fb05fbf3fae0fad5facafaa6fa7afa4ffa;
    inBuf[381] = 256'h1bfaf8f9eaf9d6f9c2f9acf984f95ff946f932f936f950f966f986f9b0f9d6f9;
    inBuf[382] = 256'h07fa42fa76faabfadffa02fb2cfb65fb9ffbe3fb29fc56fc71fc80fc81fc91fc;
    inBuf[383] = 256'hbbfcf1fc37fd82fdb6fdd8fdecfde8fde2fddefdd0fdc7fdc1fdb2fda9fdaafd;
    inBuf[384] = 256'ha9fdb0fdb9fdb0fd98fd71fd34fdf6fcc5fc9dfc8ffc91fc8ffc88fc78fc54fc;
    inBuf[385] = 256'h2dfc0afceafbd8fbd2fbccfbcefbd4fbd2fbd3fbd9fbdefbeefb0efc37fc71fc;
    inBuf[386] = 256'hb5fcf6fc3afd7dfdb8fdf3fd2efe65fe9efed3fefffe29ff4eff6cff8effbaff;
    inBuf[387] = 256'hedff280066009a00c000d200cc00bb00a5008b0076006400530046003a003300;
    inBuf[388] = 256'h340039003b00380028000300cdff8aff43ff06ffddfecefeddfe00ff2dff58ff;
    inBuf[389] = 256'h72ff74ff5eff31fff5feb7fe81fe5dfe58fe70fea5fef3fe4affa0ffe9ff1c00;
    inBuf[390] = 256'h3800440045004b0062008d00d10029018401d80119023a024302390227022002;
    inBuf[391] = 256'h2a023f025d027a02870289028102740271027a028902a302be02cf02d902d702;
    inBuf[392] = 256'hc502af0296027d027302780283029502a2029902800256022202fc01eb01f101;
    inBuf[393] = 256'h180250028602b702d702df02dc02d002be02b802c002d40208035403ad030f04;
    inBuf[394] = 256'h6104890489045c040e04c50392037f039a03d30310044d0476047e0476045a04;
    inBuf[395] = 256'h2c040204da03b503a603a503aa03c203e003f803170431043d04480446043004;
    inBuf[396] = 256'h1904fd03de03d403da03e8030a042d044204580463046504750488049b04b904;
    inBuf[397] = 256'hd404e9040c0538056b05b50501063e0672068d068e0692069806a406ca06f606;
    inBuf[398] = 256'h1b07400753074c0740072307f506cc06a3067e0676067e068c06a706b2069e06;
    inBuf[399] = 256'h79063e06f305b805890561055105430531052c0527051d051f051805ff04e604;
    inBuf[400] = 256'hbf049004750466045d04660469045e045b04560456047604a104cd04fe041605;
    inBuf[401] = 256'h11050605f004dc04ea040d0544059a05f40548069c06d306e606e606c7069806;
    inBuf[402] = 256'h7c0672067e06b006e5060e07310739072c0727071e07140715070907ee06d806;
    inBuf[403] = 256'hbd06a606a806ad06af06b406a4068006600637060e06f705da05b8059e057d05;
    inBuf[404] = 256'h5d05570556055a05690565054a052905f804c404a6048e047d047d0474046304;
    inBuf[405] = 256'h5b044d043c043704290412040404f103e203e903f203fa030b040d0403040104;
    inBuf[406] = 256'hfb03f503fe03fb03ec03dc03be039f039a03a503c403fe033204540469045b04;
    inBuf[407] = 256'h36041404f103dc03e803ff031e044904650472047b04740464045d0454044f04;
    inBuf[408] = 256'h5a0464046d04800489048d0499049e04a404b604c104c604cb04be04a1047f04;
    inBuf[409] = 256'h4d041304e403ba039f03a103ae03c003d003c0038c033e03d6026a021902e301;
    inBuf[410] = 256'hd201e801080226023a022f020502cc0180013401fd00d700ca00d800ed00fe00;
    inBuf[411] = 256'h0801f900d500aa00790051003f003b0043005700660071007f008b009b00b800;
    inBuf[412] = 256'hd600f5001701310146015d01710185019d01b001c201d701e901fd0113022202;
    inBuf[413] = 256'h270223021002f701e001cb01bf01bc01bc01bb01bc01b501aa019e018b017501;
    inBuf[414] = 256'h60014901330120010901ef00d200af008e007300600054004d0040002600fdff;
    inBuf[415] = 256'hc4ff85ff4dff25ff13ff15ff22ff30ff33ff26ff0affe5febffe9dfe86fe7afe;
    inBuf[416] = 256'h7afe83fe92fea5feb3febafeb4fea1fe88fe72fe67fe6dfe83fe9dfeb3febbfe;
    inBuf[417] = 256'hb0fe98fe7cfe65fe5bfe5ffe6bfe7efe8ffe98fe9afe93fe85fe74fe66fe5cfe;
    inBuf[418] = 256'h61fe76fe98fec7fef8fe1eff36ff39ff27ff0ffffbfef5fe08ff30ff5eff8aff;
    inBuf[419] = 256'ha3ffa1ff8bff6aff49ff3bff42ff57ff76ff92ff9fffa1ff97ff85ff78ff70ff;
    inBuf[420] = 256'h68ff64ff5dff4cff3bff25ff08ffecfecbfea0fe76fe4cfe25fe11fe0efe11fe;
    inBuf[421] = 256'h16fe0bfee1fda0fd4ffdfdfcc7fcb5fcc0fce6fc10fd28fd2dfd1cfdf5fccffc;
    inBuf[422] = 256'hadfc92fc8bfc94fca9fcd1fc03fd30fd5cfd78fd7dfd79fd6ffd65fd70fd8efd;
    inBuf[423] = 256'hb8fdeffd27fe52fe78fe97feaffecffef2fe11ff32ff4cff58ff62ff68ff69ff;
    inBuf[424] = 256'h72ff7cff81ff88ff8bff85ff7eff72ff56ff37ff10ffe0febcfea6fe9dfeabfe;
    inBuf[425] = 256'hc2fed2fedbfed1feadfe7efe4afe15fef5fdeafdedfd05fe20fe2efe2efe17fe;
    inBuf[426] = 256'he6fdaefd77fd46fd30fd31fd40fd62fd85fd9cfdacfdaefd9efd8efd7ffd73fd;
    inBuf[427] = 256'h79fd8bfda0fdbffddcfdedfdfbfd02fefcfdf8fdf4fdecfdecfdf0fdeefdf0fd;
    inBuf[428] = 256'hedfddffdd1fdc1fdacfda3fda1fd9ffda5fda9fda1fd97fd87fd71fd68fd6dfd;
    inBuf[429] = 256'h7ffda7fdd9fd04fe28fe39fe31fe21fe0efefffd04fe1bfe3bfe66fe8ffea9fe;
    inBuf[430] = 256'hb8feb7fea4fe8ffe7ffe79fe8bfeb4fee5fe1fff50ff6bff75ff6eff59ff45ff;
    inBuf[431] = 256'h36ff28ff25ff28ff27ff28ff24ff13fffbfed8fea9fe7efe5bfe43fe41fe4bfe;
    inBuf[432] = 256'h53fe53fe41fe13fedafd9ffd6cfd52fd4ffd56fd60fd60fd49fd27fdfefcd5fc;
    inBuf[433] = 256'hb9fcadfca9fcb3fcc6fcddfcfffc28fd4cfd6bfd7dfd7efd7dfd82fd95fdbffd;
    inBuf[434] = 256'hfdfd3ffe7ffeb0feccfedafee2fee4feecfef7fe00ff0aff16ff22ff36ff54ff;
    inBuf[435] = 256'h71ff8fffa4ffa7ff9eff8dff78ff6dff71ff7eff95ffadffbfffcbffd1ffcdff;
    inBuf[436] = 256'hc3ffb0ff8dff61ff2ffffafecffeb5fea6fea4fea8fea5fe9dfe8dfe74fe5afe;
    inBuf[437] = 256'h43fe2cfe1cfe16fe16fe23fe3cfe5bfe7efea2febbfecbfed1fecbfec0feb4fe;
    inBuf[438] = 256'ha5fe9bfe97fe99fea3feb7fecffeeafe04ff11ff11ff05ffebfecffebcfeb5fe;
    inBuf[439] = 256'hc2fee0fe04ff29ff47ff54ff51ff3fff1efff8fed5feb7feaafeb1fec7fee9fe;
    inBuf[440] = 256'h0eff29ff36ff35ff23ff0bfff3fee1feddfeeafe06ff32ff67ff9affc5ffdfff;
    inBuf[441] = 256'he6ffdeffcfffbfffb9ffc2ffd6fff2ff11002b003f004c005300590063007000;
    inBuf[442] = 256'h7f008e0098009d0099008f00820079007300730078007c007c00710053002300;
    inBuf[443] = 256'he3ff99ff50ff13ffeafedbfee4fefafe14ff26ff25ff0fffe5feaffe7afe54fe;
    inBuf[444] = 256'h43fe4ffe72fea2fed5fefbfe0cff0bfffbfee6fed6fed4fee3fe05ff33ff65ff;
    inBuf[445] = 256'h94ffb7ffcbffd1ffd0ffd4ffe7ff0f0048008e00d00003012001280123012001;
    inBuf[446] = 256'h2a0145017001a101c901de01d901bd019501690145012e0122011f0120011c01;
    inBuf[447] = 256'h11010001e600c2009a006f004b00390039004d006f008d009a008d0064002b00;
    inBuf[448] = 256'hf4ffccffbdffcaffe8ff09002100260018000100e5ffd3ffd6ffedff1b005700;
    inBuf[449] = 256'h9400ca00f10001010001f700ef00f4000e0136016b01a201cb01e001dd01c401;
    inBuf[450] = 256'h9e0177015501410141014f0166017f018e01900186016e015101390128012201;
    inBuf[451] = 256'h23012501250125011f011c01200129013701480153015a015e015b0153014901;
    inBuf[452] = 256'h39012a01230126013f016e01a801e301110224021d020402e501d301dc01fd01;
    inBuf[453] = 256'h34027302a802ce02e102dd02cc02b7029e028802760266025d025d025f026502;
    inBuf[454] = 256'h6a0262024d022902f801c5019a0179016801620160015e015601460132012001;
    inBuf[455] = 256'h0d01ff00f500ed00eb00ec00ef00f9000a0120013a01580174019001a901bb01;
    inBuf[456] = 256'hc901d501dd01e401ec01f101f90104021002240240025e027c0294029d029d02;
    inBuf[457] = 256'h95028a0287029202aa02cf02f8021c0339034a034a033b031c03eb02b0027102;
    inBuf[458] = 256'h3702120207020e021e0223020c02d80189012d01de00a7008c008b009500a100;
    inBuf[459] = 256'had00b900c600dc00f5000a01150112010301f500f000f8000c01240136013d01;
    inBuf[460] = 256'h38012e012e013b0152016f0185018e018c01840182019301ba01ef012b025d02;
    inBuf[461] = 256'h7e028c028702760266025b02560259025e02620264025e0249022802f701b901;
    inBuf[462] = 256'h770138010501e700da00d500d300c700ac008600560029000a00fafff9ff0500;
    inBuf[463] = 256'h15002400310039003d0044004b0055006200720083009900ad00bd00ce00da00;
    inBuf[464] = 256'he200eb00f6000801250147016c019301b301c801d201ce01c301b901b201b201;
    inBuf[465] = 256'hba01c401c701c201ab01870161013b011c010901fb00ef00e000c600a5008200;
    inBuf[466] = 256'h5f00400027001000fcffeaffd7ffc6ffbcffb4ffafffacffa7ffa2ffa2ffa4ff;
    inBuf[467] = 256'hacffbeffd3ffedff090021003800510066007b009200a700bb00cf00dd00ea00;
    inBuf[468] = 256'hf9000401110122013201450157016201650162015401400129011001f900e800;
    inBuf[469] = 256'hd800cc00c300b600a3008800600031000000cfffa6ff88ff71ff5fff4fff3bff;
    inBuf[470] = 256'h29ff1bff0fff08ff07ff03fffefef6feeafee4fee9fef7fe10ff30ff4dff66ff;
    inBuf[471] = 256'h7aff87ff96ffa9ffbdffd2ffe7fff5ff02000f001c003200520075009900b800;
    inBuf[472] = 256'hcc00da00e100e300e600ef00f700000105010201fa00f000df00cd00b8009a00;
    inBuf[473] = 256'h750047000f00d8ffa6ff78ff53ff35ff17fff9fedafeb6fe97fe7efe67fe57fe;
    inBuf[474] = 256'h4cfe45fe47fe52fe65fe84fea9fecdfeecfe02ff0aff0cff08fffffefafefbfe;
    inBuf[475] = 256'hfefe08ff16ff26ff3bff51ff63ff74ff80ff86ff88ff86ff80ff81ff88ff96ff;
    inBuf[476] = 256'hb1ffd4fff9ff1d00370043004300380021000500e3ffbcff95ff6dff47ff2bff;
    inBuf[477] = 256'h1aff0fff0bff07fffcfeeffeddfeccfec6fecefee0fefcfe19ff2fff3dff40ff;
    inBuf[478] = 256'h39ff2fff25ff1cff17ff12ff0dff0cff0aff05ff02fffafeebfed4feb3fe8afe;
    inBuf[479] = 256'h61fe3cfe21fe17fe1cfe2ffe4afe66fe7efe92fe9ffea5fea9fea8fea4fe9efe;
    inBuf[480] = 256'h95fe8bfe85fe84fe8bfe9cfeb5fed3fef8fe1aff36ff4eff5dff65ff6aff6dff;
    inBuf[481] = 256'h72ff7fff91ffa6ffbcffcfffddffe7ffe9ffe4ffddffceffb7ff9aff76ff4dff;
    inBuf[482] = 256'h23fff5fec6fe98fe68fe38fe0dfee8fdcafdb5fda5fd98fd8dfd82fd7afd78fd;
    inBuf[483] = 256'h7cfd87fd99fda8fdb3fdb6fdb2fda8fd9efd96fd93fd9afda8fdbffde0fd09fe;
    inBuf[484] = 256'h39fe6cfe99febdfed2fed7fecefebffeb0feabfeb2fec4fedffefefe18ff2aff;
    inBuf[485] = 256'h32ff2eff20ff08ffe5feb8fe82fe45fe03fec2fd86fd52fd28fd06fdecfcd8fc;
    inBuf[486] = 256'hc7fcb8fca8fc95fc81fc69fc4efc32fc16fcfefbedfbeafbf7fb18fc4efc95fc;
    inBuf[487] = 256'he9fc45fda1fdf9fd49fe8dfec5feeffe09ff12ff0dfffffeeefee4fee8fe00ff;
    inBuf[488] = 256'h28ff5aff89ffa8ffb0ff9dff72ff36fff0fea7fe60fe1ffee7fdb9fd97fd80fd;
    inBuf[489] = 256'h72fd66fd54fd37fd0bfdd3fc94fc59fc27fc03fceafbd5fbbdfb9bfb6efb3bfb;
    inBuf[490] = 256'h0afbe4fad3fadafafafa2efb6ffbb5fbf8fb33fc63fc89fca6fcc2fce3fc10fd;
    inBuf[491] = 256'h4ffda0fdfffd63fec2fe10ff44ff5aff52ff32ff01ffc7fe8bfe51fe1efef4fd;
    inBuf[492] = 256'hcefdacfd94fd83fd76fd66fd50fd32fd0cfde6fcc7fcb6fcbafcd1fcf5fc1dfd;
    inBuf[493] = 256'h3dfd4cfd46fd2bfd00fdccfc96fc66fc3ffc26fc1bfc1ffc31fc4ffc70fc8cfc;
    inBuf[494] = 256'h9afc94fc79fc50fc26fc0bfc0bfc2efc71fcc9fc28fd7ffdc6fdf8fd18fe2bfe;
    inBuf[495] = 256'h35fe3afe3afe34fe2bfe1ffe15fe12fe17fe25fe3afe51fe68fe7ffe96feaefe;
    inBuf[496] = 256'hc9fee3fef7fe00fffcfeebfed5fec2febcfec7fee1fe03ff21ff33ff36ff30ff;
    inBuf[497] = 256'h2bff36ff59ff97ffe7ff3c008600bc00de00f600130140018301d6012a027002;
    inBuf[498] = 256'h9902a1028f026d024b022f021e0213020802fa01ec01e201e401f3010d022902;
    inBuf[499] = 256'h3e0246024102380236024a027802c2021f038203db031e0440043c041304cc03;
    inBuf[500] = 256'h6e030b03b3026c0239021602f901d801b101810151012c011201ff00e900bb00;
    inBuf[501] = 256'h6a00faff72ffedfe8cfe59fe5afe83feb5fed9fee0fec9fea1fe76fe5bfe55fe;
    inBuf[502] = 256'h55fe55fe4cfe31fe18fe11fe27fe71feedfe83ff2b00ca004701ae01fd013902;
    inBuf[503] = 256'h7a02b702e60206030403dc029d024e020e02f40102024202a50207035a038803;
    inBuf[504] = 256'h840361032603e402b5029002740268025a0251025c027e02c8023a03bd034a04;
    inBuf[505] = 256'hbd04f104f104b6044404ca034f03db028f025c023d02450262028f02dd023403;
    inBuf[506] = 256'h8e03ec03300451045b044e043804260425043d04560475049e04b104bc04d304;
    inBuf[507] = 256'hd904dc04e804d704b90491043704c40342039002d6012f018d00280025005f00;
    inBuf[508] = 256'hf900e101e502f103d1046d05c405d105b505830541051805fd04e004e8040705;
    inBuf[509] = 256'h2d058405fb0580062607c4074108a908e208e908d708ae0877083c08fc07b307;
    inBuf[510] = 256'h5a070607c1068f06a106f5066e071708b40808092909e9084108740767063405;
    inBuf[511] = 256'h2a041c033902d001a001cd0171021a03c4034b043d04c703c7020f012eff16fd;
    inBuf[512] = 256'hb8fac6f817f77df576f48af380f2c8f1eaf011f004f075f0aaf126f4fdf6c5f9;
    inBuf[513] = 256'h73fc14fea7feddfed9fe59ff1b0109043308550dc3123918671d042212264829;
    inBuf[514] = 256'h822ba52c6f2c3f2b9c29ec273c273e28ee2a8f2fcd358e3c1d43c248764cd34d;
    inBuf[515] = 256'hd14c49496343bf3bd9321e297b1f9816790eb0075f0288fdeff834f4d9ed95e5;
    inBuf[516] = 256'hdddb22d056c33cb7e4ab80a2419c9098a0978399189d5fa240a9b9b0ccb840c1;
    inBuf[517] = 256'h30c984d017d7b5dcc3e191e6cbeb07f23af9dc01d40b10167f20a12a2a33533a;
    inBuf[518] = 256'hfe3f4443b8446c44ab413c3d6e37fe2f1d287820f1187412430d94083a04d4ff;
    inBuf[519] = 256'h65fa8ef36bebeae148d734cc22c148b645ac8da33b9c03975394d493aa958d99;
    inBuf[520] = 256'h389e10a39ea7e3aaccacc9adf5ade0ad5faed8af85b2a0b632bcdcc250ca7ed2;
    inBuf[521] = 256'hc7dab8e26fea3bf19ff616fb2cfeb7ffd500780191016602d10346057107ca09;
    inBuf[522] = 256'h620b970c080d1d0c560a9507700349fefaf735f086e730de42d48fcac5c102ba;
    inBuf[523] = 256'hcab384afcaac61ab17ab12abe6aa87aa91a951a856a795a6bfa655a8efaa51af;
    inBuf[524] = 256'h87b5efbce0c51ed091da04e50fef7bf75afec80369071d0a5d0c060ed70f9c11;
    inBuf[525] = 256'h96122813e5123c110d0f5a0cd8085a059601e5fcb8f79ef110eacde1f1d871cf;
    inBuf[526] = 256'h53c6fdbd62b631b0aeab88a8dea6c9a6cfa76da974ab69ad7daec0ae95aeb5ad;
    inBuf[527] = 256'hb0acbeacc3adb3af69b333b8d0bc6bc161c56cc725c800c88ec61dc5c5c4f3c4;
    inBuf[528] = 256'h7cc60bca15ceebd225da37e275e987f06bf72dfe1806680f021a9126b6347b43;
    inBuf[529] = 256'h72529560906cc075bf7b587efc7d9e7b27784c74e970476eab6b9b687c64cf5d;
    inBuf[530] = 256'hfb532647c13642231c0ee6f7c8e19acdfabb7fad0fa3419c7e987d972798a799;
    inBuf[531] = 256'hcd9b349e40a1e4a54daca9b46abf30cc71daede9fef9160a371a1b2a5939f747;
    inBuf[532] = 256'h6f555261b26bf673d8798e7d127f6a7e257cab781474c46e0e69d5620b5cc654;
    inBuf[533] = 256'hdd4c2644bd3aae30e825a71a500f080437f996ef63e7c8e04bdcd7d9f9d8ced9;
    inBuf[534] = 256'hf6db94dea6e113e522e8feeaf7ed83f0c3f226f536f702f90bfbeefca8feb400;
    inBuf[535] = 256'ha2023c04e7053407bb07d20739079d057e030a011dfe39fbcff8e0f6bef5bbf5;
    inBuf[536] = 256'hcaf6d3f8e5fbc1ffe7031e08170c5a0fd811b713f114d615e6162b18c319ed1b;
    inBuf[537] = 256'h651ed4202e23162525265b268f2574231020721b81156d0e92063cfedef5ebed;
    inBuf[538] = 256'h9fe638e0dada55d68bd278cfe6ccc2ca31c928c8b7c71ec854c947cb22ceded1;
    inBuf[539] = 256'h71d602dc82e2c4e9bbf116fa7602ac0a67126619a01fef243b29ba2c772f6831;
    inBuf[540] = 256'hbc3274336833b5328331c42f8d2d0e2b46282225ab21d91d8d19d014c00f740a;
    inBuf[541] = 256'h3205520001fc60f897f594f32ff25ef100f1e4f01af199f117f288f2edf20ff3;
    inBuf[542] = 256'h01f31bf370f328f49af5b7f750fa61fd97009e037b0615095b0b990df70f6612;
    inBuf[543] = 256'hf814a5172d1a721c681ef11f13210022d4228f234b241525ba2516261b268125;
    inBuf[544] = 256'h2b243522821f0f1c2418c513fb0e240a5905ac007dfcd2f879f580f2aeefa9ec;
    inBuf[545] = 256'h6de9f6e54ae2c6deaddb2ed99cd70ad755d764d801daf1db21de85e020e305e6;
    inBuf[546] = 256'h29e978ecd5ef11f313f6cef839fb75fd92ff8a017e036105020761086309da09;
    inBuf[547] = 256'hf309c40925093908fc062505d1021e00ecfc9bf992f6bff363f1afef3fee02ed;
    inBuf[548] = 256'h00ecc7ea51e9d4e716e62ee467e2a2e0f5de8cdd34dc06db35da9cd95cd998d9;
    inBuf[549] = 256'h0fdabbda87db1ddc84dcbfdcb6dcb6dce1dc24ddd0dddede0de08ae137e3d1e4;
    inBuf[550] = 256'ha3e6b0e8bbea13eda5ef0ef26ff4a8f65af8b9f9d0fa62fbb4fbddfba5fb45fb;
    inBuf[551] = 256'hcffa15fa4bf97ff870f738f6d4f4f4f2a2f0dfed7deab7e6cbe2c4de07dbd4d7;
    inBuf[552] = 256'h1bd51dd3e1d119d1e9d046d1d3d1bdd208d45bd5ebd6b6d85eda24dc24de17e0;
    inBuf[553] = 256'h67e242e55ae8ecebe7efb6f36ef7fafae0fd5e008002ed03dd044005be04a503;
    inBuf[554] = 256'hfc0198fffafc3ffa41f769f4a7f1a9eebbebb6e842e5ade1fcdd01da2fd6bad2;
    inBuf[555] = 256'h8fcf07cd44cb1fcabec92bca2ccba4cc76ce63d033d2d5d34fd58cd6a9d7f6d8;
    inBuf[556] = 256'h5bdad0db9bdd75dfe9e02ae209e312e3abe20fe2f1e0d1df2cdfc3defbde40e0;
    inBuf[557] = 256'h07e24ae43fe716ea81ecf2eefdf09ff2e0f410f87dfc3a038d0c281809266135;
    inBuf[558] = 256'hc8443b53985fc4685a6e7c709c6f7a6c12685e63d65ebf5a39579f53394fa649;
    inBuf[559] = 256'hf0416f37692acc1af8086bf60ae4cdd277c4aab97bb260afaaaf4fb2e0b654bc;
    inBuf[560] = 256'hfbc114c84aceb1d412dc56e4a1ed86f85b048310271dd82961360743414fac5a;
    inBuf[561] = 256'h5a65986edc75457b6a7e007f7e7d157ad2744b6e0767415f5957c24f9a48cf41;
    inBuf[562] = 256'h713b5d35232f9528b921611ab612430b400406fe43f90bf62ef4e6f3e9f491f6;
    inBuf[563] = 256'hfbf8fbfbc9fe81013f043f068e078d089e08d107ca062e051d035f01b7ff23fe;
    inBuf[564] = 256'h40fdb8fc49fc55fc81fc7cfc9afc9dfc38fcb8fb20fb65fae0f9eaf9bffa96fc;
    inBuf[565] = 256'h91ffba03c7085f0e3e14d319a61ea5229325562748287f280d28562770266125;
    inBuf[566] = 256'h7424a323c022d621af20df1e431cbc1811144c0eb407820009f9cdf12aeb4ce5;
    inBuf[567] = 256'h71e0b1dcfcd960d8ced726d872d988db32de6fe106e5c1e8b7ecc9f0e1f43cf9;
    inBuf[568] = 256'hcbfd84029e07e80c3712a917e61c9f21e4256129bf2b1f2d582d432c322a5027;
    inBuf[569] = 256'hb823d81f031c581809153912e70ffc0d660c0c0bb9094c08d0063a05a6036102;
    inBuf[570] = 256'h860126017d01830211043206cf08920b5f0e1a115c13f714fc154116c815ed14;
    inBuf[571] = 256'hb9132a1299100f0f5f0dc30b4b0ada08ba070e07b506ca063807b6074308d908;
    inBuf[572] = 256'h6909140aef0a0a0c6d0d040fd810e312fa1436179619d61b031efe1f5321f421;
    inBuf[573] = 256'hc5216d20121ef11a1317e312b40e9a0ad0065a030b00ebfcdef9bcf69cf36ef0;
    inBuf[574] = 256'h34ed27ea4ee7d3e412e311e2eee1d6e28be4dfe6bae9b7ec9cef67f2ecf42cf7;
    inBuf[575] = 256'h56f969fb6cfd64ff3001b602df039304e204d3045f04a903c502af017a0018ff;
    inBuf[576] = 256'h6cfd82fb50f9c6f61bf472f1c5ee47ec11eaf4e70de67fe424e31fe29ee16de1;
    inBuf[577] = 256'h89e100e27ee2ede267e3b1e3e0e336e492e402e5a5e539e6afe607e710e7f2e6;
    inBuf[578] = 256'hcce67ce63ee60ee69de507e535e4eee29ae165e047dfbfdedcde59df67e0c4e1;
    inBuf[579] = 256'hf7e23ee48be5a4e6fce7a2e957eb5eed8fef7ef149f3d9f4faf5f5f6d3f764f8;
    inBuf[580] = 256'hd6f815f9e7f86ff8b2f78df630f5aaf3def1efefebedb2eb60e910e7b8e492e2;
    inBuf[581] = 256'hbfe022dfe5dd13dd63dcf7dbeddb0cdc93dcb1dd1adff0e050e3c6e554e8f9ea;
    inBuf[582] = 256'h41ed43ef14f173f2c1f33bf5a2f63bf80afa9cfb12fd54fef3fe2cfff9fe14fe;
    inBuf[583] = 256'hd5fc2cfbd6f844f67ff367f09fed4beb39e9cce7e5e602e642e58fe496e3a1e2;
    inBuf[584] = 256'he2e143e1f0e0f8e020e158e1aae104e273e233e351e49fe51fe7afe8c3e93dea;
    inBuf[585] = 256'h3bea73e9ede72de62ce4dfe1c0dfd8dde6db3bda09d918d8a9d7fcd7bed8e6d9;
    inBuf[586] = 256'h8edb2bdd8fde04e039e12ce2a3e3c5e5c0e88fed81f471fdbd082216b724e733;
    inBuf[587] = 256'hd04232503b5b3e63bf67da68fd66e4627d5da1571452264dc048a144f73fd139;
    inBuf[588] = 256'hb531f9265e199f0962f881e699d5b7c699ba36b2b1adb5ac05afc1b302ba37c1;
    inBuf[589] = 256'h75c85bcf0bd648dc6fe243e9c4f033f90203b40df918d624a830123c20474951;
    inBuf[590] = 256'h2d5ac4617467c06abf6b556a7266a6609c59b9519149da41c93a5a34d42e202a;
    inBuf[591] = 256'hc125a321aa1d5619a514d90fdb0aed05ab0127fe7bfb23fa0efae1fab8fc4aff;
    inBuf[592] = 256'hd6015704b1062208bf08c808b3079505e90263ff26fbd4f659f2dced0feafee6;
    inBuf[593] = 256'hb5e49be389e33de4b6e59ce793e985eb4cedcfee2df0acf199f322f68ef915fe;
    inBuf[594] = 256'h7c0395094510f816391dda225327522adf2bcd2b2a2a5c279e235b1f101bdd16;
    inBuf[595] = 256'heb124f0fd60b6a08e8041301dafc33f810f389edb0e7bee107dcc2d645d2e3ce;
    inBuf[596] = 256'habccc3cb40ccf6cdd2d0a4d413d9f5ddfee2d1e771ecb5f065f4c1f7d1fa79fd;
    inBuf[597] = 256'h0f00b40267058a084a0c95108c15eb1a2020cf2475287c2ace2a8529c2260023;
    inBuf[598] = 256'he01eba1ad7168a13ef10ec0e810d990cea0b410b790a3f095807c5049001eefd;
    inBuf[599] = 256'h65fa78f78df500f5f1f512f8fffa55fe7f0126044e06c7078508d608a808cb07;
    inBuf[600] = 256'h8c060005230383018100440037015f035906ef09b70d30114414e416fe18c81a;
    inBuf[601] = 256'h631cd41d211f47204c212b22e822c223c224d5251d275928fb28d0288027b124;
    inBuf[602] = 256'h9d20801b9b158e0fb70939045fff1bfb45f704f444f1f9ee51ed27ec3deb7cea;
    inBuf[603] = 256'h94e953e8e6e674e552e410e4ece4f4e628ea2bee89f2faf631fbfafe69029105;
    inBuf[604] = 256'h6808dd0ad80c270ea10e4c0e540df10b6b0a16091a086207cd061e06f6042903;
    inBuf[605] = 256'hbf00c1fd7afa40f71bf42ff19aee14eca3e992e7c5e571e408e45ce446e5cee6;
    inBuf[606] = 256'h63e896e960ea77eadee901e9f9e7fce64fe6bde539e5cbe442e4bde370e352e3;
    inBuf[607] = 256'h97e33ee4f3e49de5ece578e577e418e388e176e042e0eee0aee23ae5fae7c9ea;
    inBuf[608] = 256'h6ced9eef89f130f382f4a9f586f6e1f6d9f673f6c2f52cf5daf4c5f40ff589f5;
    inBuf[609] = 256'hc4f59df5f3f496f3c2f1b0ef70ed4ceb64e98fe7e6e569e4dce27de18ee0f9df;
    inBuf[610] = 256'h05e0e4e045e227e472e6abe8d4eaefecacee42f0d9f130f37df4d3f5e9f6f8f7;
    inBuf[611] = 256'h0ef9f0f9e8faf8fbd4fca5fd3bfe36feccfde3fc58fba2f9d9f7fef596f495f3;
    inBuf[612] = 256'hbcf249f2f9f172f1f3f066f0abef1fefc5ee6cee40ee27eee2ed82ed0ded70ec;
    inBuf[613] = 256'hd0eb58eb09ebe6ea08eb69ebe2eb82ec3fedc6ed16ee36eebceda3ec38eb4be9;
    inBuf[614] = 256'hefe6ace47ce24be093de52dd3ddc90db4adb02dbddda04db28db8bdb91dcf7dd;
    inBuf[615] = 256'hdfdfa7e2d6e52de903ed21f187f507fb1502f40a3616cc230c332443db52cb60;
    inBuf[616] = 256'hd36b21736676ca75ef71ee6bbd64435d69566750204b8546b641bc3b27341e2a;
    inBuf[617] = 256'h231dd20da2fc7bea37d926ca59be09b751b4beb5d9ba47c2d7cad5d335dcb6e3;
    inBuf[618] = 256'hbfea1cf135f7eefd1f05e70ccb15561f4c29ef33a73e17496353d25cd4646d6b;
    inBuf[619] = 256'hf96ff371a4710e6f2e6ab663425c2454e94b2e443c3d39376832d62e282c0c2a;
    inBuf[620] = 256'h402828264f23da1fd91b73177a137510690ebf0d750ec20f79116513a8144d15;
    inBuf[621] = 256'hac152e15ee136f120b109c0cb508ee0340fe8af8dff27bed45e956e6aae4aee4;
    inBuf[622] = 256'h1ce69ee847ecadf06cf573fa5dffdf03e807570b5a0e4a116a143318da1c3622;
    inBuf[623] = 256'h3328532ec7331e38df3a8f3b553a7d373d33142e7d28b722021d7e173612350d;
    inBuf[624] = 256'h7508fa03ceffe0fb24f890f403f166edc1e927e6c0e2c1df58dd9bdb9fda6eda;
    inBuf[625] = 256'h01db70dce0de40e292e6c9eb5df1cff6d7fbddff97024b040305f804dd04eb04;
    inBuf[626] = 256'h34051d0695075209700bb00da80f47114a12491258118f0ff10ce909fc067104;
    inBuf[627] = 256'h9902ba01c1016c0296030d058606fa078c09350bf60cda0ead102d124613ed13;
    inBuf[628] = 256'h28144814a5145d157e16f1174a192e1a6d1ad11957183e1691135110af0c9808;
    inBuf[629] = 256'hfd0339ff99fa6ef648f36cf1d8f084f10df3f6f4f7f6c6f85cfa02fcdbfd1900;
    inBuf[630] = 256'hf30231069609fe0c1c10e2127915ec17721a3c1d1420b622c524b82548257423;
    inBuf[631] = 256'h6720981c8918a7143b113f0ea50b6009340726056f03f901cf00030019ffcafd;
    inBuf[632] = 256'hf6fb78f9a4f617f442f26cf1dff160f367f58df74af926fa20fa63f91ff8b4f6;
    inBuf[633] = 256'h63f524f4d2f249f162ef0ced76ea05e802e693e4e6e3dee314e45ae48de48ae4;
    inBuf[634] = 256'h9ce414e5f7e56ee777e98eeb83ed49ef9af0aff1f4f26df456f6def884fbf3fd;
    inBuf[635] = 256'he0ffa3001a0073feaefb42f8bff43af1faed0deb05e8e7e4b1e12ddec9dae2d7;
    inBuf[636] = 256'h63d59cd38ed2aad1e4d029d031cf71ce61ce12cfe7d0e7d383d773db5adfbee2;
    inBuf[637] = 256'hb1e554e8a8eaf5ec39ef2ff1bff29df38df3cbf27cf1dcef7dee82edd3ec8cec;
    inBuf[638] = 256'h5eecccebd8ea68e95fe73ee553e39ae172e0dedf6cdf30df23dfe9ded4de37df;
    inBuf[639] = 256'he0df0de1d5e2aee47de62be83fe9dde948ea5aea66ea9feab6eabdeaacea2dea;
    inBuf[640] = 256'h7ce9bde8cde713e7a3e631e6f5e5bae509e52ae41fe3c0e1b8e04de04ee028e1;
    inBuf[641] = 256'hb8e255e416e6d9e729e964eacaeb14ed7eee0df039f1e3f1fcf138f1c2ef01ee;
    inBuf[642] = 256'h23ec6aea1de92be862e7a4e6c1e567e47de216e018dd8fd9e2d52ed26cce08cb;
    inBuf[643] = 256'h24c882c570c329c25ac121c1b0c185c281c3dbc432c69cc7aec94dcc96cf1bd4;
    inBuf[644] = 256'h7cd953dfe6e5deecf2f3d5fbe4043b0f5f1b3529fc37f546f954c0606a69476e;
    inBuf[645] = 256'h266f756cdd66625f10579f4eae466a3f8738c1318a2a1c2228185e0c90fe50ef;
    inBuf[646] = 256'h4edf66cffcc032b5deaccca8fba8efacf6b3c7bc55c607d00dd961e18ce96ef1;
    inBuf[647] = 256'h4af9bf01690a0613e41b87249e2c8e34303c53434f4ad5505456b05a7b5d205e;
    inBuf[648] = 256'hb65c74595454ba4d6746b13eef36fa2f452acc25f922ed21ef218c2261236323;
    inBuf[649] = 256'h0822871fe31b8717831357101f0e2c0d300d5a0d5d0dee0c700b02090f067402;
    inBuf[650] = 256'h6afe72fa3df698f1d8ecd0e76fe253ddc2d8e7d452d23bd1a7d1c5d376d786dc;
    inBuf[651] = 256'hd7e206eabbf1a5f93b011e08150eed12de164a1a8a1d1c2132259729102e0a32;
    inBuf[652] = 256'hc834da35f334fd31512d562791208e199412f30bd5051200cefa29f6e7f124ee;
    inBuf[653] = 256'h0beb56e8f7e508e44ae2a2e034df06de24ddbfdcf1dca8ddd9de8ce094e2ebe4;
    inBuf[654] = 256'hd5e739ebf6ee3df3abf7a6fb2affd00117036003e602b1018400daffadff6300;
    inBuf[655] = 256'h14024804e906c9096b0cb50ea4100e1200139613d313cc13b613d5136d14c815;
    inBuf[656] = 256'h1a183e1bd71e72225b25f026fd266f257222a31e8c1a8c1602130010640d2b0b;
    inBuf[657] = 256'h43099c075d068b05f1047304d903d0024a0177ff84fdd6fbf1fa1afb7bfc1bff;
    inBuf[658] = 256'ha002a406da0adb0e8312fd155019861cc71fdf2273255f2773289228f027eb26;
    inBuf[659] = 256'hdb25fd2472241f24a923c3224f212d1f741c74194c161113de0f910c2909bd05;
    inBuf[660] = 256'h7d02a6ffa0fdb2fcd2fc14fe1200370233049e052f062006a805ed0453040204;
    inBuf[661] = 256'hd803d203d703b4037f0360035c0396030a0467045d04ae032102c4ffe0fcdef9;
    inBuf[662] = 256'h33f72df5f9f39bf3d4f376f465f56af67bf7b8f801fa46fb81fc61fdb7fd85fd;
    inBuf[663] = 256'hb2fc71fb2cfa09f93ff801f80ff82cf82bf8a7f77cf6d3f4c5f299f0a6eefdec;
    inBuf[664] = 256'h98eb5deaffe867e7abe5e3e36ae2a0e18ce12de268e3d0e422e653e73ce8fae8;
    inBuf[665] = 256'hd6e9d1eaf5eb54eda9eed2efe9f0d9f1cdf220f4d0f5daf735fa75fc3afe3cff;
    inBuf[666] = 256'h29ff05fe0bfc8bf910f7fcf47bf3b1f25bf223f2f4f18ef1e6f055f0e3efa4ef;
    inBuf[667] = 256'hceef13f037f044f0f3ef56efdfeea9eee8eedbef3bf1ccf260f4a0f588f62df7;
    inBuf[668] = 256'h9cf72df8eaf8c3f9b9fa8dfbf9fb04fca9fb0afb7efa3ffa78fa2cfb2efc47fd;
    inBuf[669] = 256'h15fe68fe4cfe9efda3fcbefbcbfafef981f9dcf838f8cdf746f708f75bf7c9f7;
    inBuf[670] = 256'h7cf85df9c5f9dff9a0f9c2f8d0f7f1f611f6b4f5b4f5b8f5eaf5e1f555f587f4;
    inBuf[671] = 256'h5af3f5f1baf0a7efeeee8dee36eeeeed62ed60ec55eb14eab8e8e9e733e75ae6;
    inBuf[672] = 256'hdde524e5ebe3efe2f8e1e3e05ae02ae0f2df01e032e030e03ee0aae057e165e2;
    inBuf[673] = 256'h4ee4d2e68ae9f1ece3f0f2f40cfaa1006e0854127e1ef22b643ae848cc554460;
    inBuf[674] = 256'h8d67116b416b9c68f063465e0c58df51024cf745d53f4e3984319f28671e4112;
    inBuf[675] = 256'he704c4f611e853da8dce59c5e9bf60be55c086c5b7ccefd4a4ddc2e53ced77f4;
    inBuf[676] = 256'h1dfbbb01e30812105f17df1edf25692cac327638103ea74306490a4e6052b655;
    inBuf[677] = 256'hb2570e58fe5675547050a04b2446fe3f083a8e349a2ff62bcd29cb28ec28b129;
    inBuf[678] = 256'h542a5a2a682973278324fa20941d681aa917d11538146e12aa101d0e9a0aea06;
    inBuf[679] = 256'hb00214fef0f9b8f542f116edade809e4d3dff8dbdad805d763d63cd79fd940dd;
    inBuf[680] = 256'h4ce292e8b2efc4f74600a408b310d117a81d6d220726be281b2b372d502f7231;
    inBuf[681] = 256'h3d337634a33441334e30ae2b9725bf1e76172b107309390381fd82f80af426f0;
    inBuf[682] = 256'h16ede0ea8ee906e911e97ee9e9e936ea8ceacbea30eb12ec25ed59eebbefcaf0;
    inBuf[683] = 256'h6ff1e9f116f22bf2a6f285f3b1f43ff6f2f748f91bfa70fa17fa4ff9bdf878f8;
    inBuf[684] = 256'haff8d5f9a2fbbefd66004b0323064809970ccc0f0413e8150e187319031ade19;
    inBuf[685] = 256'h76191a192019ad19941aaa1b841ca91c001c611ac5178d14ea10030d29095705;
    inBuf[686] = 256'h7901a2fdcff925f6e8f23ff065ee66ed0ded4aede0ed8fee6def8af0f7f1f4f3;
    inBuf[687] = 256'h92f6c8f983fd77017e0583095b0d2011dd146818c11ba81ebc20f4211d220221;
    inBuf[688] = 256'hf61e181c7a18b114fd10650d3f0a91071505dc02d900ddfe05fd64fbd6f963f8;
    inBuf[689] = 256'h0ff7b3f54ef40ff305f25df165f113f240f3ddf47af6b0f77ff8ccf89af842f8;
    inBuf[690] = 256'hd6f754f7d7f628f62df5faf367f2a0f0edee39edceebe5ea3deaf0e902eafee9;
    inBuf[691] = 256'hfce908eacfe9a2e9bbe9dde95cea5ceb6decaded20ef59f07af1abf2a5f378f4;
    inBuf[692] = 256'h12f50ef567f41df30ef18beee2eb25e9a6e682e46ce26fe07bde3fdce9d9b5d7;
    inBuf[693] = 256'h89d5b2d36cd266d1afd04cd0d3cf65cf42cf35cf8ccf92d0edd1a7d3cbd5c8d7;
    inBuf[694] = 256'h9ed967dbcedc16de79dfa9e0d7e1f9e293e3dae3e2e370e313e308e30fe38de3;
    inBuf[695] = 256'h6ee422e5e1e590e6c5e6f0e622e715e733e76fe761e750e71ae762e686e586e4;
    inBuf[696] = 256'h34e3fde1efe0e0df21df9dde11deb1dd6cdd1cdd12dd58ddcadd99dea6df9ce0;
    inBuf[697] = 256'h8fe175e21fe3d4e3cde4ece567e74ce943eb49ed54ef0af177f2a3f33cf461f4;
    inBuf[698] = 256'h23f447f31ef2e0f06bef24ee32ed4becb6eb72eb1debf6eaebea97ea44eadde9;
    inBuf[699] = 256'h0fe946e88ae7a2e610e6e6e5e4e56fe687e7d9e899eaaaeca6ee8ff030f237f3;
    inBuf[700] = 256'hb1f39ef3faf2faf1bff059efdced56ecd7ea5be9f0e7b4e67fe53ae4f4e268e1;
    inBuf[701] = 256'h6cdf35ddbcda03d87cd569d3d3d108d131d110d293d3b2d50dd880da26ddc6df;
    inBuf[702] = 256'h4fe210e5d8e77eea71edaef036f4cff8dcfe710609107f1b0a280f3585413b4c;
    inBuf[703] = 256'h7d54b459a05b955afe568f51254b4e44aa3d9037d231642ceb26b42085190f11;
    inBuf[704] = 256'hff06bbfbaaef4be3c5d7f0cd7ac644c26ac1a0c399c84bcfcdd69cdedde569ec;
    inBuf[705] = 256'ha8f262f8dafda3035409ce0e6914bb19ae1eb823af288a2d9e32af377f3c2741;
    inBuf[706] = 256'h5f45bf482f4b774c3d4c764a64473f43603e76390f356431c92e6f2d052d452d;
    inBuf[707] = 256'h012eb12ed72e5a2e022d902a4e278f23471fd21a97164312da0da40937059b00;
    inBuf[708] = 256'h5bfc3ef857f42ff15deeafeb7be94ee700e508e334e1a1dfefde15df57e041e3;
    inBuf[709] = 256'h9ee772eddff43afd1106210f8717c71ec2241229c02b372da62d672df02c6c2c;
    inBuf[710] = 256'he42b552b9f2a8229c4276d258022fa1e2e1b55176e13c90f9c0cca098107de05;
    inBuf[711] = 256'ha904dd039e03ca0343042805610681076b081809160950081d074705d3024400;
    inBuf[712] = 256'h59fd09faf9f60bf445f157ef2bee8cedceed77eef0ee65ef9aef70ef72efc6ef;
    inBuf[713] = 256'h89f038f2e0f4a6f8ecfd9204750c7715e01e022863304737443c5c3f88400140;
    inBuf[714] = 256'h433ea53b7e3838351c325c2f142d362b7b297827d1244a21e51cf317fb127b0e;
    inBuf[715] = 256'hd60a5108ef067c06d406d00711097c0a130c740d800e600fb40f600fce0ed20d;
    inBuf[716] = 256'h6b0c1c0bbc092908cf06930577040c0454044e054d070c0a3a0dca103e143617;
    inBuf[717] = 256'h9919221be71b331c241c2c1c901c431d831e3e201a221824ef252827d427d027;
    inBuf[718] = 256'hf2269125bd236321d21efd1bcd1889151f128c0e1f0bcd078d04a601fbfe71fc;
    inBuf[719] = 256'h3dfa5af8c1f6a8f5fbf481f41bf48ef3aef2a6f1c1f03ef077f0a1f194f311f6;
    inBuf[720] = 256'hdcf886fbb5fd4eff34005c00efff1bff06fee5fcf2fb5afb23fb51fbddfb79fc;
    inBuf[721] = 256'hf2fc51fd65fd34fd0bfdd1fc7cfc47fcfbfb8afb43fbf9fa94fa43faadf992f8;
    inBuf[722] = 256'h20f72ef5cbf25af0e7ed8eeb6fe94fe71fe5d3e23fe0aadd55db4ed9ffd789d7;
    inBuf[723] = 256'hbcd7bad85fda53dca6de21e171e3b6e5cee791e951eb1aede3eefdf060f3e2f5;
    inBuf[724] = 256'h95f83bfb85fd64ff9700fc00bf00e1ff89fe12fd8dfb05faadf869f70cf6b0f4;
    inBuf[725] = 256'h49f3b9f135f0d2ee71ed2cec08ebcce995e884e779e6ade550e533e575e529e6;
    inBuf[726] = 256'h03e70de850e982eab5ebfbec1fee44ef6ff063f136f2c7f2d4f296f20bf225f1;
    inBuf[727] = 256'h65f0dcef6aef64ef9eefbdeffdef43f068f0dcf09df188f2dff360f5aaf6dbf7;
    inBuf[728] = 256'hc1f822f956f982f9a3f905fac7fab3fba6fc73fdbdfd3cfde7fbc8f9faf6e2f3;
    inBuf[729] = 256'hdbf003ee8eeb85e99ce7c6e513e44ee29de04fdf2ede1ddd3ddc34dbb9d90cd8;
    inBuf[730] = 256'h3fd64ed4aad2a5d12ad168d180d223d44ad616d93ddcc0dfe5e363e820ed5ef2;
    inBuf[731] = 256'hcef747fd2d0388097d10aa184522492da739aa464653615eb066526be86b7468;
    inBuf[732] = 256'hb661b8586f4e04443c3a4b315e293722431b2d147d0cd7034cfae5eff7e44cda;
    inBuf[733] = 256'h7ad050c8c9c248c019c158c542cc23d542df47e989f2edfae0019907ef0cd211;
    inBuf[734] = 256'h67163e1bec1f0024be27e62a422d562f55312d3335357d37a2398a3b253d123e;
    inBuf[735] = 256'h2c3eb13da33c083b5139d0378136bb35d4358e36ce37a5398a3bef3cc43da33d;
    inBuf[736] = 256'h0e3c42396a356730b22aaf24281e371700102208b4ff2af799ee7ee685dfbcd9;
    inBuf[737] = 256'h46d552d276d079cf5ecfcdcfccd095d208d553d8b1dce7e111e850ef3ef7c8ff;
    inBuf[738] = 256'hde08cc11281ab821cd270d2c9c2e612f7a2e6a2c972937269822f51e311b2017;
    inBuf[739] = 256'hd412470e6909a40450007bfc89f9aaf782f615f666f6f0f6b0f7e6f843fabefb;
    inBuf[740] = 256'h9bfd97ff660114037104230520056b04d8025f0033fd5bf9d7f4f4efdceaa0e5;
    inBuf[741] = 256'hade057dcb4d828d6e2d4abd484d55ad7c0d9a0dc03e0b9e3d5e77eec9cf128f7;
    inBuf[742] = 256'h08fdfe02e4087a0e8313f217981b4a1e242030216e212a219a20c31fcb1ebf1d;
    inBuf[743] = 256'h751cd31ad018471627138a0f800b2407bf028ffec0faa0f764f503f48cf3f5f3;
    inBuf[744] = 256'heef443f6d9f76bf9cffa16fc46fd5dfe7fffd60061021204f105e007a409320b;
    inBuf[745] = 256'h7d0c670d070e6e0e980ea30e960e490ec70d0c0df30b980a2709b20765067605;
    inBuf[746] = 256'hf904ec043f05ea05c00692075d080b097509ac099a090e091e08c106eb04f302;
    inBuf[747] = 256'hfc0012ff7ffd2ffcecfacaf99bf836f7d7f57cf421f303f20bf128f07cefe5ee;
    inBuf[748] = 256'h78ee6eeeacee4bef6bf0bdf130f3c9f43cf690f7dcf8eaf9d7faa7fb20fc6bfc;
    inBuf[749] = 256'h9bfc85fc65fc53fc14fccdfb7ffbebfa3dfa7df981f87df774f62df5d4f36ef2;
    inBuf[750] = 256'hcaf023ef92ede2eb3aeaaae8f1e631e596e3fee194e08edfb5de0ade9edd27dd;
    inBuf[751] = 256'ha3dc37dcbbdb4edb1fdbfadaeada05db07db09db2ddb41db70dbc4dbeddb0fdc;
    inBuf[752] = 256'h2ddcffdbe0db06dc3ddcf0dc3bdeb1df84e1a5e39ae59de7b0e973eb28edcaee;
    inBuf[753] = 256'hf5efeaf0b0f108f252f29ef2b4f2c8f2b0f209f2f7f05bef12ed87eae0e719e5;
    inBuf[754] = 256'h98e25de031de4edcb2da36d92dd8bbd7bfd770d8e0d9c8db2ede16e12ae459e7;
    inBuf[755] = 256'h98ea8bed1bf03ff2b3f38ff4f5f4caf44ff4b1f3c3f2bff1bcf07bef44ee30ed;
    inBuf[756] = 256'hf7ebe5ea05eaf7e817e888e7f6e6d6e652e701e82ee9e1ea8fec66ee66f01bf2;
    inBuf[757] = 256'hb5f33cf553f628f7bcf7c1f76ff7d5f6c7f58ef44af3e6f1a5f0a8efd5ee43ee;
    inBuf[758] = 256'heaed8ded0ced56ec54eb10eac1e893e798e6fce5bee596e579e562e50ce590e4;
    inBuf[759] = 256'h42e4fde3bae3b2e39ee326e374e28de14ee011df2ede8bdd4fddb6dd6dde5ddf;
    inBuf[760] = 256'hbae029e286e32ee5efe6ade808eb2aee34f2fef7ebfffb096816cb243334b443;
    inBuf[761] = 256'h0a52ee5d7666ec6a346bc467516117594850ab47024063393b33212d4826d81d;
    inBuf[762] = 256'hbf13f707c6fa3bed2de06cd424cbcac4a9c124c2c1c5fccb70d4dfdd7ce7f6f0;
    inBuf[763] = 256'h56f97300e306610c2b111316c31afc1e16238426df28a12acd2b802c842d1b2f;
    inBuf[764] = 256'h2931e0330537e9393a3ccf3d573ee23dfd3c153c783b9f3bbd3c883eb8401443;
    inBuf[765] = 256'h1e457046fd46a4463445de42c93fd43b3a374332ca2cff263221141b9814e90d;
    inBuf[766] = 256'h9a06b7fedcf620ef14e8aae2ecdef9dc08dd52de53e0e9e250e57ce7f2e988ec;
    inBuf[767] = 256'ha2efe8f3ebf888feea044b0b4f1119171e1c21205b237c256326602668258023;
    inBuf[768] = 256'h01211a1ede1a7c172f14fe10dc0d0b0bbf08f10601064d06b707570a3e0edf12;
    inBuf[769] = 256'hc917b01cdd20ce238225e125e924062391208a1d131a6e167112030e67098c04;
    inBuf[770] = 256'h4affe6f962f49eeef6e89ce3afdec0da27d801d78ed7a6d9eedc25e1dce5e5ea;
    inBuf[771] = 256'h60f037f6b0fc2c04610c2b156e1e3b27df2e203548391f3b303ba239bd364233;
    inBuf[772] = 256'h5f2f0b2b972602221e1d1e181e13120e160941048cff06fbe3f67df343f1b5f0;
    inBuf[773] = 256'h57f253f66dfc3b04f90c96155e1dd4237a286a2b1e2db12d692dba2c712b4f29;
    inBuf[774] = 256'h8826f6228d1ee0193d15cf100d0d080a9107b70559045803e202170323043606;
    inBuf[775] = 256'h3d09240da6113716a81ac51e2222ec244e27ef28e7294f2a9c29b827d924cf20;
    inBuf[776] = 256'he91bcf16c411280d56092906720301018afe09fc97f962f7c7f5f3f4eff4dbf5;
    inBuf[777] = 256'h81f79bf931fc17ff120241057f08710bfd0def0ffa102b11ac109a0f370eb90c;
    inBuf[778] = 256'h300b9609d007c70562038d0074fd46fa24f76df462f2f8f04ff067f0e1f0a7f1;
    inBuf[779] = 256'hc1f2dcf3fcf460f6def76bf939fb0cfda7fe1f004701ec012502dd01ec0051ff;
    inBuf[780] = 256'hfafce6f93df631f216ee3beac4e6dde37fe160df75ddaadbd3d93bd838d7d6d6;
    inBuf[781] = 256'h6ad727d9b8dbfcded3e2c7e6b5eaa8ee71f218f6a5f9e2fcbaff06028a035204;
    inBuf[782] = 256'h58048f033b026300f5fd2efb0cf87cf4dbf04eede2e906e7dbe443e382e282e2;
    inBuf[783] = 256'hece2e0e34ae5d0e69de8c9ea0ced7fef2ff2b4f4e6f6b3f8caf92afa0cfa8df9;
    inBuf[784] = 256'he9f862f8fef7b1f74cf773f613f52bf3bcf02beec6eb95e9e2e7aee6aae5f0e4;
    inBuf[785] = 256'h87e435e443e4dde4cae537e728e940eb95ed29f0aef240f5cef7faf9c6fb05fd;
    inBuf[786] = 256'h68fd23fd44fcc6fa2af99df70ef6daf4e5f3cef2b2f166f099ee9aec94ea87e8;
    inBuf[787] = 256'he8e6ebe56be57fe507e697e61ae784e7aae7b0e7d4e70ee867e8fae89ee914ea;
    inBuf[788] = 256'h64ea88ea43eaa6e9e8e8cce735e666e43ee28ddfc6dc2adaabd7bcd5a4d41bd4;
    inBuf[789] = 256'h2cd4e6d4d7d5f1d66cd802dab3dbd5dd20e06ce212e513e88feb4bf0d0f679ff;
    inBuf[790] = 256'hb70a6d18f42760384a4844560c618c676169d26679609957a94dcb430d3bfd33;
    inBuf[791] = 256'h652edc29a525c220961ab512fb08e4fd08f239e6aadb39d3a7cdb3cb53cd30d2;
    inBuf[792] = 256'hc1d9bce212ec0ff5a5fca0028b07400b1f0e0e11cd132c16a818de1a831c251e;
    inBuf[793] = 256'hc41f582171230b26ec28422cce2f153304366e38f6398d3a663aa53977385137;
    inBuf[794] = 256'haa368a3609374b38e1395b3b943c073d503c943ac337e933932f052b5e260422;
    inBuf[795] = 256'hf61de719c6154611ff0b06067aff75f896f161ebf9e5c1e1d7ded5dca0db22db;
    inBuf[796] = 256'hf7da33db14dc71dd75df52e2a8e55fe98dedbff1cff5ebf9b5fde9009f038e05;
    inBuf[797] = 256'h8406c4067406bf050d059504560441043304e5031103bc01050004fe24fcecfa;
    inBuf[798] = 256'h84fa2ffb24fd0a008f036f07fd0ace0dc70f9b104110050fe50cf90988069b02;
    inBuf[799] = 256'h4afed1f955f5f6f0c8ecc2e8dee401e126dd7bd934d6a6d33cd221d268d305d6;
    inBuf[800] = 256'h97d9bfdd37e2a6e6f6ea40ef90f31df80dfd4202ac070f0de711f215ef18861a;
    inBuf[801] = 256'hd11a021a2b18b115f21201101f0d820a0e08db05090471020301c2ff89fe49fd;
    inBuf[802] = 256'h17fc0dfb57fa2bfab8fa10fc14fe99005e03f5051408a2096f0a8d0a4f0ad109;
    inBuf[803] = 256'h3209bf086b0804089e071a073d062e050e04d402b301e1005a00360096007101;
    inBuf[804] = 256'hb3027704a6060409810bf80d1a10cd111513d3130f140014a51302133a122a11;
    inBuf[805] = 256'hb30fe00d920bd108de05ca02bcffecfc3bfaa4f73bf5cef276f074eeb6ec6beb;
    inBuf[806] = 256'hd1eaa4ead1ea5bebd7eb3cecc5ec51ed0dee3fefb4f05cf225f4a9f5d9f6b3f7;
    inBuf[807] = 256'h02f8f8f7b5f718f767f6b4f5bef4d0f3f2f2daf1d7f0faeff4ee21ee9fed1bed;
    inBuf[808] = 256'he3ec0eed21ed43ed85ed7aed5eed6eed61ed63ed9bedb0eda0ed7eed10ed69ec;
    inBuf[809] = 256'ha9ebb9eab3e995e83ee7b9e5f8e3ede1d2dfb1dd8cdbaad911d8b3d6c9d549d5;
    inBuf[810] = 256'h17d560d507d6d6d6edd728d953daaadb1cdd81de20e0f1e1b2e39ae59be762e9;
    inBuf[811] = 256'h0ceb91eca7ed79ee19ef5aef76ef81ef4def12efdfee7dee34ee16eed7ede0ed;
    inBuf[812] = 256'h12ee18ee45ee68ee49ee0deec6ed44edc4ec70ec21ecf8eb10ec2eec58ec94ec;
    inBuf[813] = 256'hb7ecd0ece8ecf3ec16ed58ed9dedf9ed55ee7cee7aee59ee06eeb0ed7eed57ed;
    inBuf[814] = 256'h53ed7aed84ed5eed16ed7deca6ebdeea31ead5e913ead1ea03ec99ed38efc0f0;
    inBuf[815] = 256'h22f22bf306f4cbf467f515f6bcf611f745f727f77cf6baf5d7f4a8f3b3f2d5f1;
    inBuf[816] = 256'haff0b0efb9ee7fed8fecf4eb69eb50eb9debeceb56ecc8ec04ed16ed17ed15ed;
    inBuf[817] = 256'h21ed5eedf2edb7ee9cefa3f04ef165f11af123f0a1ee4bed1cec19ebafea81ea;
    inBuf[818] = 256'h0aea50e911e823e6e5e3aae1aadf3ede89dd76dde6ddb1de8fdf56e024e1f5e1;
    inBuf[819] = 256'hcfe228e450e685e980eec5f57fffe30baa1a072beb3bd24b5c595c63c3689269;
    inBuf[820] = 256'h33664f5f6d56f24ccd43f73bce35d6309c2c5c280a23431cd313cb0902ff40f4;
    inBuf[821] = 256'h74eadae2f7dd38dc02deb9e2d7e9eff296fcf305bb0ec815d41a7b1e6c20ef20;
    inBuf[822] = 256'h1e21ea205b202320fe1fa11f791f7a1f921f3520802147238a252128972aa72c;
    inBuf[823] = 256'h602eb72fa4309f31f53287349f367639a03cfd3f9343d4465949184bba4bf64a;
    inBuf[824] = 256'h0049034608426c3d8f387733502e50293a24f91eae1909140c0e18080f0238fc;
    inBuf[825] = 256'h33f7e7f276ef43edceebe7eac5eadcea32eb48ecc9ede1ef09f39af658fa6bfe;
    inBuf[826] = 256'hfd01be0401076508f1082e09090997083808ea07b707b407ef077a082f090e0a;
    inBuf[827] = 256'h220b010cac0c620dc60d0a0ebe0eb40f15114913e615b818ae1b2e1efe1fe820;
    inBuf[828] = 256'hbe208f1f621d6f1ae616f012b10e760a3f061d025afee2faadf7e8f46cf23ff0;
    inBuf[829] = 256'h8eee52edcbec1bed29ee31f006f343f6fbf9cffd4f01bd04e5079b0a740d5910;
    inBuf[830] = 256'h1313131602195d1b5f1db51ef31e751e3e1d371be418891643146f123811a810;
    inBuf[831] = 256'hd0109211ca123f14a615e116cf175518be185719501a1e1c181f1d230228712d;
    inBuf[832] = 256'h9332a33626398a399e37d933ac2e9f289422ff1c0218e2138310940d160bea08;
    inBuf[833] = 256'hfe06780549047a0334035603fb0364057d076f0a610ef812ff17251dab214025;
    inBuf[834] = 256'hb327a0284028f526bd24eb21c31e201b1c17ca12140e4509b4049e0078fd83fb;
    inBuf[835] = 256'hbdfa36fbaffccdfe5e01fd03620698087b0af60b3a0d2c0ead0ee70ec80e260e;
    inBuf[836] = 256'h510d370c930a8e080f06ea0240ff27fbbbf64ef227ee8aeabde7d3e5cce487e4;
    inBuf[837] = 256'hb2e42ce5e7e5b9e6b4e700e98fea6beca2ee08f17ef3e8f50bf8d1f935fb0efc;
    inBuf[838] = 256'h57fc27fc81fb87fa5df90af8adf652f5eaf389f234f1dbefa3ee94ed8feca7eb;
    inBuf[839] = 256'hdaeaf6e91de96de8d5e78ee7b7e721e8d2e8b8e985ea38ebc9eb0cec36ec65ec;
    inBuf[840] = 256'h7deca6ecdfeceaece7ecd7ec96ec65ec56ec47ec6fecbbeceaec1fed45ed24ed;
    inBuf[841] = 256'h02ede7ecbbecccec13ed57edc8ed4bee97eee6ee3aef5bef87efcdeff6ef2ef0;
    inBuf[842] = 256'h77f095f0b0f0d5f0cdf0c2f0d0f0c7f0caf0f6f01bf151f1adf1eff11ef242f2;
    inBuf[843] = 256'h16f2abf115f119f0e3ee9eed1cec92ea38e9dee7b3e6e2e522e597e460e42ce4;
    inBuf[844] = 256'h21e45ce491e4e4e464e5c5e537e6bfe60be75de7c9e705e852e8b4e8d5e8f9e8;
    inBuf[845] = 256'h20e9ffe8dfe8bfe85de80ee8d7e772e741e74de758e7bde782e852e95cea8feb;
    inBuf[846] = 256'h8dec74ed43eeb1eedfeee4ee9aee21ee9aedeeec20ec40eb36eae6e85ae79de5;
    inBuf[847] = 256'h9fe37ce17cdf9ddddfdb95dabfd91cd9d1d8dcd8ddd8ead825d94bd971d9d2d9;
    inBuf[848] = 256'h3ddabfda99db97dcb2dd31dfefe0f4e2b7e55fe914ee50f43efcd6050d11761d;
    inBuf[849] = 256'h6f2a2e379e42e24b445221558454e950d74a5a43963b2f34c62da22861249620;
    inBuf[850] = 256'hbe1c1e185e12720b860340fb5df3a6ecf8e7cfe57ae60feaf9ef9ef75300d908;
    inBuf[851] = 256'h60108316751a261c2d1c8f1acd17ed141512770fac0d840ccd0bc10b1c0cb70c;
    inBuf[852] = 256'he10d750f45117b13f1157e18311bfb1dd520cd23f126592af22d9d315e35e238;
    inBuf[853] = 256'hc53bf23d223f0b3fd33d863b28381734892f982a93259520981bbe16f211150d;
    inBuf[854] = 256'h4b08790389fec3f938f5f1f04fed64ea20e8c4e636e622e69de678e74ae83be9;
    inBuf[855] = 256'h4dea24ebf6ebf8ecdcedadee93ef3af08bf0a5f05ef0b5efe6ee0eee49edbbec;
    inBuf[856] = 256'h70ec62ec85ecd7ec4eedd1ed76ee4def39f05cf1d7f290f4a4f635f91afc50ff;
    inBuf[857] = 256'hd00247068609590c630e7f0f970f920e9e0ce5099006020370fff6fbd2f8f5f5;
    inBuf[858] = 256'h45f3dff0aaee97ecdeea82e994e850e8b7e8cbe9a6eb23ee2ef1bcf47ff845fc;
    inBuf[859] = 256'he0fff802720543074f08d208f408b7085d08020887071507b1062e06af053b05;
    inBuf[860] = 256'hc20466042604f90309046204fc04ec052c079d082b0aae0b0e0d460e3d0f0510;
    inBuf[861] = 256'hbf1061110112ae123e139e13c1137713bb12a21133109c0e110dad0b8f0acb09;
    inBuf[862] = 256'h580935095909c1096f0a500b5f0c9a0ddc0e1210471170128f13bf14f9152c17;
    inBuf[863] = 256'h4d183519be19c9192a19dd17f8158913b710bb0db10abc07ff0474021e0006fe;
    inBuf[864] = 256'h1bfc5afacbf85ff71af611f53af495f32bf3f1f2e1f208f35bf3ccf34ff4c5f4;
    inBuf[865] = 256'h1ff55cf571f569f55af549f537f525f504f5d5f4a1f462f41af4dbf3adf398f3;
    inBuf[866] = 256'h97f3a2f3b7f3d3f3eff3fff3f5f3cff397f348f3e8f28cf241f20cf2f4f1f3f1;
    inBuf[867] = 256'hfef10bf20cf2fbf1dff1bcf19af182f178f178f175f161f139f101f1bdf06bf0;
    inBuf[868] = 256'h23f0eaefabef6def22efb5ee1cee60ed88eca4ebcbea08ea6be9fee8b3e88de8;
    inBuf[869] = 256'h8ee8afe8fee886e933ea04ebfbebf2ece2edd5eebbefa1f0a7f1c8f20df47df5;
    inBuf[870] = 256'he8f639f863f93efacffa38fb79fbacfbeefb2ffc73fcb9fce0fce6fcd2fc8bfc;
    inBuf[871] = 256'h28fcc0fb3ffbb5fa2dfa8bf9e6f852f8bef740f7e2f688f647f62cf619f628f6;
    inBuf[872] = 256'h73f6d4f658f711f8d0f895f965fa15fbabfb32fc7dfc8ffc74fc06fc5bfb96fa;
    inBuf[873] = 256'ha5f9a1f8a7f792f66ff549f4fbf2a7f173f04def6deef6edc1ede8ed6dee09ef;
    inBuf[874] = 256'hccefb2f073f126f2cdf220f34cf363f328f3ddf2acf260f238f25cf28cf2ecf2;
    inBuf[875] = 256'h87f3fff355f482f42cf463f34af2d3f04aef02ee04ed87eca6ec31ed05eef8ee;
    inBuf[876] = 256'hb6ef0ff0e8ef37ef0eee7eecc4ea0be954e7e1e5d3e4fae37ce362e34be346e3;
    inBuf[877] = 256'h51e317e3c3e279e201e2aae1afe1cce145e25de3cae4c8e6b3e970ed3cf26ff8;
    inBuf[878] = 256'he8ffab08b6128a1dbf28d033c83def45bd4b844e2d4e1e4bc145f43ec737eb30;
    inBuf[879] = 256'hf82a4726a522c31f2d1d571afd16f6123f0e43095e040f001efde2fba8fcd0ff;
    inBuf[880] = 256'hde04480baf12cd19b51f38246a260f26f8231320c91a84157610ec0b01098707;
    inBuf[881] = 256'h3c07a0081e0b2b0e09121f16031a0c1edb214225ad28f32b112f6032bc352039;
    inBuf[882] = 256'h9b3cce3f8d42ac44b5459c456844ee416e3e3f3a83358c30b12b1427e7224c1f;
    inBuf[883] = 256'h461cdb19ee174b16de147913e1111710210ef50bc809cd0702069904af031403;
    inBuf[884] = 256'hc702d202da02d8020003cf025202db01e8007fff12fe3ffc17fa2cf845f673f4;
    inBuf[885] = 256'h3df37af21df273f244f35ef4d2f562f7e1f853faacfbe9fc13fe3aff6d00a601;
    inBuf[886] = 256'hf902840443064408980a230dc00f341234147815af15cb14ea121310af0c3609;
    inBuf[887] = 256'hcd05e002c60053ff9efea9fef9fe74ff0b005a00710073003f0024006100ec00;
    inBuf[888] = 256'h0802b603b8050908650a730c2d0e510fbd0fb40f2d0f3c0e420d400c300b4e0a;
    inBuf[889] = 256'h8309b208f7074a07a4062b06eb05f805630621072a087209dd0a510cb10ddf0e;
    inBuf[890] = 256'hcd0f6c10bc10d110bd109e109110ac10f6106211dc11491275124d12cf11f610;
    inBuf[891] = 256'he10fbf0eab0dda0c7d0c910c190d190e680fe5107112dc130415e7158816e516;
    inBuf[892] = 256'h1f174f177a17a717c617c2178a170f1745162d15d01329124610380efd0ba109;
    inBuf[893] = 256'h4207ee04bd02c30004ff8efd61fc6ffbc3fa68fa43fa48fa77faacfad2fae7fa;
    inBuf[894] = 256'hcffa88fa23fa8ff9d2f811f847f77cf6cff52bf58af4fff368f3b4f201f238f1;
    inBuf[895] = 256'h5cf09feff7ee79ee53ee66eea7ee2fefcfef7ef055f128f2f2f2bef352f4abf4;
    inBuf[896] = 256'hd8f4b9f471f427f4ccf392f389f380f38ef3aaf39af383f369f329f3f4f2c3f2;
    inBuf[897] = 256'h65f204f28ef1d5f013f04bef5eee8bedccecf3eb28eb66ea82e9b4e80fe87fe7;
    inBuf[898] = 256'h38e73ae74ee785e7d9e710e84ee8aee80ce986e92deac0ea45ebc8eb10ec34ec;
    inBuf[899] = 256'h5bec5bec52ec60ec54ec49ec5cec5fec7aecc9ec18ed86ed19ee8fee06ef7eef;
    inBuf[900] = 256'he3ef65f0e0f01bf14df179f16cf173f19bf1b6f105f285f2f6f287f32df4aff4;
    inBuf[901] = 256'h3cf5c5f512f647f658f61af6c5f569f5f8f4adf495f48ff4aef4e2f4f8f4fcf4;
    inBuf[902] = 256'he6f490f410f466f372f256f134f007ef0fee7fed3bed4fedb1ed02ee27ee16ee;
    inBuf[903] = 256'h96edcdecf7eb12eb64ea27ea35eaaeea99ebadecf7ed6befb9f0f1f101f3a1f3;
    inBuf[904] = 256'hfbf313f4c2f357f3eaf253f2ddf189f11af1c3f078f0fdef81ef03ef5beebeed;
    inBuf[905] = 256'h30ed98ec1fecc4eb70eb3eeb1eebfdeae7eac8ea9bea6cea25eacfe977e900e9;
    inBuf[906] = 256'h81e812e89ee745e725e71ee73de78be7dae72ce88fe8e6e840e9bee94deaffea;
    inBuf[907] = 256'hf7eb21ed95ee88f0fbf213f60afacefe5c04b60a84117f18691faf25e82ad42e;
    inBuf[908] = 256'h013156311030522d90297c257321dc1d111bf81867172d16d9142c130311430e;
    inBuf[909] = 256'h200bdf07d30486024b015e01ff02ef05ca09460e9e123516da180f1aad191818;
    inBuf[910] = 256'h5915b411df0d170ab00650040c03f6024f04c606ff09dc0dd1117c15d518951b;
    inBuf[911] = 256'had1d5c1f9c2088216e22472329243e255a2663275028ce28af28f02766261f24;
    inBuf[912] = 256'h5c213b1efb1aed172d15e1122911f50f440f0b0f0e0f300f480f0e0f780e880d;
    inBuf[913] = 256'h290c970a06096c070106da04b903b202cc01c400c1fff0fe20fe7afd28fde4fc;
    inBuf[914] = 256'hb4fcabfc7cfc28fcccfb3cfb93fa06fa8df94df96ef9cbf958fa02fb88fbd7fb;
    inBuf[915] = 256'hedfbc3fb7afb34fbfdfaecfa05fb3cfb99fb26fcebfcfbfd5fff0901d0028704;
    inBuf[916] = 256'hf705e3063107e7060406ac0418036301bdff62fe62fdd4fccefc2cfdc9fd8afe;
    inBuf[917] = 256'h2fff95ffc2ffb4ff89ff75ff98ff0c00de00ff015c03d8044b06a107ba087309;
    inBuf[918] = 256'hc0099909f208e8079f063405da03bb02df014e010501e100ce00c100a7008500;
    inBuf[919] = 256'h6e0069007e00b7000d017001d5012e027202940294027e0258022c0219022702;
    inBuf[920] = 256'h5302aa0219038303e5032a043c042c04ff03b20366032403ec02d602ed022d03;
    inBuf[921] = 256'ha4034f041b05f705cd068f073508c5085309e909860a300bd30b560cb50cda0c;
    inBuf[922] = 256'hbc0c6b0cda0b070b030ab9082a077805a003b701ebff36fe9ffc44fb08faeef8;
    inBuf[923] = 256'h17f86bf7eaf6aff68df669f650f617f6abf531f59cf4eef350f3c2f23ff2e4f1;
    inBuf[924] = 256'ha6f176f15cf143f119f1e2f094f031f0d3ef86ef5cef6aefa9ef1df0bdf070f1;
    inBuf[925] = 256'h3cf21df3fbf3e8f4ddf5b2f675f71df883f8c6f8f3f8f6f803f92bf950f995f9;
    inBuf[926] = 256'hf1f924fa3efa31fabef90cf92df8fef6c0f592f45bf352f284f1c2f02bf0bbef;
    inBuf[927] = 256'h38efc5ee66eef0ed8fed4ded04edd7ecc7ecb2ecb6ecd6ecfbec47edb6ed26ee;
    inBuf[928] = 256'ha9ee28ef74efa5efbaefacefb0efd9ef20f0aaf06df145f23ff341f41ff5eff5;
    inBuf[929] = 256'ha3f61bf785f7e8f731f893f816f994f92afacafa3afb95fbd9fbe1fbe6fbf8fb;
    inBuf[930] = 256'heefbf6fb0bfceefbbefb7ffbfafa5dfabaf9ebf822f87af7d5f666f642f63ef6;
    inBuf[931] = 256'h75f6e2f64af7bcf738f896f8f4f85cf9b2f90afa5ffa8cfaa3faa3fa77fa43fa;
    inBuf[932] = 256'h0cfabcf96df920f9baf85af810f8c4f792f77cf757f72ff703f7aff654f610f6;
    inBuf[933] = 256'hd3f5caf50df671f6fcf6a5f726f883f8bdf8b0f883f84df8fcf7bbf791f757f7;
    inBuf[934] = 256'h29f7fff6aff65ef613f6b5f574f553f533f52cf528f5fdf4b9f442f480f390f2;
    inBuf[935] = 256'h70f12df000eff6ed2eedd4ecd7ec3aedffede6eee1efdff09df11cf26ef270f2;
    inBuf[936] = 256'h4cf236f221f238f29ff232f3f6f3eaf4dbf5c7f6b9f79ef891f9b3fa02fc99fd;
    inBuf[937] = 256'h8dffd8018a04a107ff0a940e2d1281156918ac1a161cb81c9a1cc51b7f1aee18;
    inBuf[938] = 256'h1f174d158413b8110e10850e0a0dc80bbb0ad40947090e091c09a7099b0ae00b;
    inBuf[939] = 256'ha20db60ff6118a142b17a319101c1b1e8c1f98200321b9202220301ff41def1c;
    inBuf[940] = 256'h191c781b621b991bf01b861c001d341d541d301dd81ca41c791c701cc61c391d;
    inBuf[941] = 256'hca1d9b1e5d1f1c20ff20b9215422f522462353234b23ef225422bb21f4201520;
    inBuf[942] = 256'h571f821e981dba1c9f1b391aa918b5166e141a12ab0f560d720bee09e5088508;
    inBuf[943] = 256'h8908e808b309970a890bae0cb50da20ea60f7d102911e5116e12b912fc12ec12;
    inBuf[944] = 256'h7912d411bf103a0f8a0d930b72097c07a005f503b802c5011b01df00e3002601;
    inBuf[945] = 256'hc3018e028603c1040a065807b908f109ed0abc0b2d0c320ceb0b450b410a1609;
    inBuf[946] = 256'hc5075606f904b50385029401e80072004f007500c1003d01e3019c028603aa04;
    inBuf[947] = 256'hfd058d073f09ec0a8b0cf00d020fda0f6710a710c210a2103610a50fd90ed60d;
    inBuf[948] = 256'hd60cd70bdd0a150a6409b9083408ba074507f806c0069106810677066c067706;
    inBuf[949] = 256'h8906a806e8062f077707c607f80708080608dd0794074107d3064d06c3052e05;
    inBuf[950] = 256'h98041f04c60394039803c60313047c04f2046b05e7056806f60699075d084909;
    inBuf[951] = 256'h550a6e0b8c0c8c0d4e0ece0efa0ebd0e280e3a0de70b500a820885068a04b302;
    inBuf[952] = 256'h0a01b9ffc4fe09fe82fd0ffd7efcd2fb09fb1dfa3af975f8d2f76df736f70ff7;
    inBuf[953] = 256'hf7f6c9f66ef6fcf56ef5c7f42ef49bf309f388f205f27cf103f18ff02df0f3ef;
    inBuf[954] = 256'hd1efd4ef0ef06ef009f1e8f1f3f22cf482f5c1f6e6f7e6f8a2f942fad7fa51fb;
    inBuf[955] = 256'hcbfb43fc87fc9dfc80fc10fc6bfba4faacf99ff88cf75bf628f502f4dcf2d2f1;
    inBuf[956] = 256'hf4f02cf086efffee79eef8ed7fedfaec7fec1fecd4ebbdebeeeb56ec05edf4ed;
    inBuf[957] = 256'hf3eef1efd8f078f1d0f1eaf1b7f156f1e3f05df0ecefaeef9defd5ef5df009f1;
    inBuf[958] = 256'hd1f19cf232f397f3d1f3d5f3d0f3e2f302f450f4d3f465f516f6e6f6aaf770f8;
    inBuf[959] = 256'h30f9b3f9f7f9f7f98ef9def80df81ff746f6a4f51ff5bdf47af41ff4a9f326f3;
    inBuf[960] = 256'h7af2bdf116f175f0e9ef8fef49ef1fef2fef5fefbcef63f02cf110f21af317f4;
    inBuf[961] = 256'hfcf4e2f5a6f651f705f8a2f826f9a6f9f4f90efa10fad9f97ef927f9b5f83bf8;
    inBuf[962] = 256'hd6f75af7d6f667f6e1f55cf5f5f486f427f4f4f3bcf393f385f356f313f3caf2;
    inBuf[963] = 256'h48f2abf111f154f09befffee57eec1ed4bedc4ec4aece5eb64ebe4ea70ead9e9;
    inBuf[964] = 256'h47e9d0e851e8f4e7c8e79de78ce79ae799e7b2e7f7e74be8d3e890e94dea11eb;
    inBuf[965] = 256'hcdeb4deca9ece9ecfdec0fed2bed3fed69ed9fedc2edebed0cee06eef7edd1ed;
    inBuf[966] = 256'h79ed19edadec2beccdeb96eb7eebbbeb3fecf3ecfbed36ef7ef0eaf150f386f4;
    inBuf[967] = 256'ha3f57ff605f759f76ef74ef738f728f729f767f7b8f707f860f891f898f89ef8;
    inBuf[968] = 256'h9cf8b0f810f9a8f97dfa96fbbefcecfd2aff5b009501ef025604d6056a07e808;
    inBuf[969] = 256'h570aa30bb20c9e0d620ef30e7b0ff70f5610c01026116e11b811f111fc11fd11;
    inBuf[970] = 256'he4119e1159111311c710ad10c61008119a1165124a13571467155c164c171f18;
    inBuf[971] = 256'hc6186719ed194b1aac1af61a201b521b6e1b591b2f1bc41a021a1519f017a016;
    inBuf[972] = 256'h6a1547143e137a12d8114c11f910c110a610d4102b11a7115b121013b5135a14;
    inBuf[973] = 256'hc614fd141b15f3148d140c143d132612e810570f860da90bb309d50752061e05;
    inBuf[974] = 256'h4e04f403d003cc03df03d803bf03b503ae03c40308045504a404ea04ff04ec04;
    inBuf[975] = 256'hbf046a040804ab034103d9027e021f02c70180013201dc007e00030075ffe7fe;
    inBuf[976] = 256'h63fe03fedffdf7fd47fec4fe50ffd6ff46009200bd00cb00be00a10073002d00;
    inBuf[977] = 256'hd9ff77ff0affa9fe5dfe26fe0dfe06fef9fde2fdb1fd64fd10fdc5fc97fca0fc;
    inBuf[978] = 256'he2fc56fdf7fda7fe51ffebff58009700ad0094006200360016001a005300a900;
    inBuf[979] = 256'h10017901bd01d601cc01a20178016f018f01e70177022303dc038b0410056505;
    inBuf[980] = 256'h840566052205c70460040d04d703b803be03e003090440047c04a304b604a604;
    inBuf[981] = 256'h5404c6030103080201010f0038ff93fe1dfeb3fd4cfdd8fc43fc9efb01fb6ffa;
    inBuf[982] = 256'h06fad2f9c3f9dff921fa6dfaccfa3afb9cfbfffb5ffca2fcd6fcfafcf5fcd8fc;
    inBuf[983] = 256'ha3fc43fccefb4dfbbafa37fad3f989f973f98ff9caf92dfaaafa27fbaffb33fc;
    inBuf[984] = 256'ha2fc0cfd69fdacfdeafd18fe2bfe35fe31fe12fef5fdd8fdb5fda6fda6fda6fd;
    inBuf[985] = 256'hb4fdc3fdbefdb2fd94fd54fd05fda5fc2efcbafb50fbedfaaafa8afa82fa9ffa;
    inBuf[986] = 256'hd6fa10fb50fb84fb96fb91fb70fb30fbecfaa9fa66fa30fafef9bdf975f920f9;
    inBuf[987] = 256'hc0f870f83df828f83ef874f8b3f8faf83ef97bf9c1f917fa76fadffa43fb8dfb;
    inBuf[988] = 256'hb9fbc7fbb5fb95fb70fb41fb0cfbcbfa72fa0afa9cf92ff9d3f892f864f845f8;
    inBuf[989] = 256'h32f81df806f8f8f7ecf7e7f7f1f7fbf704f814f825f83df870f8b6f814f98ef9;
    inBuf[990] = 256'h12fa97fa1dfb8efbe6fb27fc43fc3afc1afcdbfb87fb32fbd0fa66fafcf97bf9;
    inBuf[991] = 256'he2f836f868f786f6a5f5c5f400f470f310f3edf20ef356f3bff33cf4a9f403f5;
    inBuf[992] = 256'h48f569f57ef599f5b4f5e5f531f680f6d5f622f749f74df72ef7e1f682f61ff6;
    inBuf[993] = 256'hb8f563f520f5daf49af454f4f9f39bf33af3d4f282f241f20ff204f21ff261f2;
    inBuf[994] = 256'he1f290f35cf443f51ff6d6f670f7dcf727f875f8c4f822f9a6f936facefa79fb;
    inBuf[995] = 256'h19fcb4fc58fde6fd65fedefe2eff63ff91ffa6ffc4ff0a006500f200b9018c02;
    inBuf[996] = 256'h76036c043d05fe05b8064c07e8079c084a09160aff0ad90bc60cc50daf0eb20f;
    inBuf[997] = 256'hc810c511cc12c71382142615a315d215ed15ea15ab1573154015ff1400154015;
    inBuf[998] = 256'ha1155b1647172a182b19211ae11ab01b791c231df51dcf1e8a1f66203921e021;
    inBuf[999] = 256'h9b223d23a02300242b240224d2237a23f12291223622d221ae21972174218c21;
    inBuf[1000] = 256'ha621ae21e4210722fe210422d7216b210b218d20f81fa51f681f401f6b1f9a1f;
    inBuf[1001] = 256'hb21fd91fbc1f4c1fca1e021e0a1d321c4b1b5e1aa419d418eb171c172b162915;
    inBuf[1002] = 256'h5e149d13fc12b01272123d122912e7117511fe104e10810fce0e060e3c0d960c;
    inBuf[1003] = 256'hd90b150b750ac7092709bc084c08e10791071e079a062c06af0545051305eb04;
    inBuf[1004] = 256'hda04ee04f004f20408050c05120527051905ef04b3044004b8033c03c0026902;
    inBuf[1005] = 256'h4c024402590285029d02a902ac028a0256021502b3014401cf004900cbff65ff;
    inBuf[1006] = 256'h0fffe4feecfe17ff72ffefff7300f7006b01b501dd01e201c301970163012a01;
    inBuf[1007] = 256'hfb00d300af00990089007d007a0076006b005c0041001700e5ffa1ff4efff4fe;
    inBuf[1008] = 256'h90fe2ffee8fdbffdc7fd0bfe7afe0cffafff3e00b000010128013c0154017301;
    inBuf[1009] = 256'haf010c027902f4027403de03350476048d0482045804fa037703d20202021f01;
    inBuf[1010] = 256'h3a004bff6dfea9fdeffc50fccefb55fbf5fab3fa74fa43fa19fad2f977f907f9;
    inBuf[1011] = 256'h6bf8bff713f75df6bef545f5e1f4acf4b1f4d4f428f5a7f520f695f6f7f614f7;
    inBuf[1012] = 256'h00f7c5f650f6cef55bf5e5f491f469f448f43ff44df441f430f421f4f1f3caf3;
    inBuf[1013] = 256'hc4f3c8f3fbf365f4d1f448f5bbf5ecf5ecf5c4f54ff5bcf425f471f3d0f25bf2;
    inBuf[1014] = 256'hf0f1b8f1bbf1c0f1d5f1eff1caf17ef11cf18af00af0c9efb3eff9efa1f065f1;
    inBuf[1015] = 256'h4df23ff3edf364f4a4f479f40ff481f3b4f2eaf148f1b7f06cf077f09cf0ecf0;
    inBuf[1016] = 256'h54f187f192f177f108f179f0ebef44efbbee67ee1beefeed18ee36ee7ceef4ee;
    inBuf[1017] = 256'h68eff5ef9df025f1acf139f29ef200f36df3aff3e2f30af4eef3b5f377f314f3;
    inBuf[1018] = 256'hc8f2b2f2abf2d4f22ef375f3b8f3f5f3f0f3cef39ff340f3e0f29df257f23bf2;
    inBuf[1019] = 256'h60f298f2fff296f31af497f407f52cf521f5f4f485f408f4a3f344f320f352f3;
    inBuf[1020] = 256'haaf339f4eef478f5d3f5f0f596f5e9f40af4f0f2e2f110f169f01df034f076f0;
    inBuf[1021] = 256'hedf085f1fef163f2b5f2caf2caf2c8f2aaf296f299f28af281f27df24df209f2;
    inBuf[1022] = 256'hb1f123f183f0deef1def6aeed2ed36edb7ec53ece8eb94eb56eb14ebefeae7ea;
    inBuf[1023] = 256'he1eaf9ea2ceb63ebc1eb47ece1eca8ed8bee63ef36f0e6f055f19bf1b6f1a9f1;
    inBuf[1024] = 256'ha2f1aaf1c3f10ef27cf2fbf295f327f499f4f1f41af513f502f5f0f4f9f44bf5;
    inBuf[1025] = 256'he3f5c6f6f5f745f99dfaf5fb26fd34fe32ff1300ec00d101ac02890370044705;
    inBuf[1026] = 256'h22060e07f307e808e909d10aa80b5d0ccc0c0f0d280d0e0df00cdd0cc60cd40c;
    inBuf[1027] = 256'h020d320d850ded0d510edb0e850f3c1034115f12a4132515bb1631189719ba1a;
    inBuf[1028] = 256'h701be51b081cdc1bb11b861b591b631b7a1b781b7a1b481bc91a341a72199018;
    inBuf[1029] = 256'he41765171f175817e417aa18c619ec1af31bf61cb41d1d1e661e5e1e0b1eaa1d;
    inBuf[1030] = 256'h121d541cb11b061b601af51988190f19a61807182c1747163015031407131612;
    inBuf[1031] = 256'h4511bd103b10bc0f590fd10e2e0e9b0dec0c3d0cbf0b440be10ab60a850a550a;
    inBuf[1032] = 256'h3a0af50992092b099308e50746079006e1055505c0043604c8034503c3025302;
    inBuf[1033] = 256'hcc014c01e7007f00330018000c00250064009900c200cd008700faff2eff1dfe;
    inBuf[1034] = 256'hfffc02fc37fbccfacffa1efbadfb52fcd0fc16fd11fdb2fc1bfc69fbb6fa32fa;
    inBuf[1035] = 256'hf3f9fdf957faeefaa0fb55fce7fc33fd2ffdc9fc06fcfbfabef972f83ff73cf6;
    inBuf[1036] = 256'h7ff511f5e3f4ecf419f552f599f5e9f53ef6a5f614f778f7c8f7e9f7c7f771f7;
    inBuf[1037] = 256'hf1f662f6fdf5ddf512f6aef68ff784f866f9ecf9dcf924f9a7f76df5b3f2aeef;
    inBuf[1038] = 256'hb9ec4eeac1e863e875e9e5eb7aefdff376f8a7fcf6ffe70147023401e3fecafb;
    inBuf[1039] = 256'h8ef8acf59bf3b8f201f354f46bf6c4f8e5fa76fc17fdabfc51fb2ff9a3f62af4;
    inBuf[1040] = 256'h22f2eef0e1f005f246f46df7fdfa72fe5001150375036a021100c6fc18f98af5;
    inBuf[1041] = 256'h9cf2baf00cf08ff01ff265f4fbf68bf9b5fb37fdf9fdf1fd32fdf3fb6cfad3f8;
    inBuf[1042] = 256'h6cf75ef6baf58cf5c4f537f6cbf65bf7bef7f4f701f8ecf7e0f700f855f8fcf8;
    inBuf[1043] = 256'hf3f917fb58fc95fd9efe67ffe4fffbffbcff34ff5afe4efd2dfcfcfae6f90af9;
    inBuf[1044] = 256'h61f801f8e5f7e3f7f4f70af801f8ecf7dcf7c5f7cbf7f8f730f87df8d3f807f9;
    inBuf[1045] = 256'h21f91ff9e2f881f805f857f796f6d0f5f5f42ef48cf3fdf29ef272f251f24cf2;
    inBuf[1046] = 256'h5bf25bf26af28df2b1f2f8f268f3e3f382f43bf5ecf5a7f664f701f894f814f9;
    inBuf[1047] = 256'h62f998f9b3f9a1f986f96bf949f945f963f991f9e6f955fac0fa38fbaefb0afc;
    inBuf[1048] = 256'h65fcb6fcedfc22fd4cfd5afd64fd64fd52fd4ffd5afd70fdacfdfffd56febafe;
    inBuf[1049] = 256'h10ff42ff5fff59ff35ff11fff0feddfef0fe21ff67ffc7ff27007800bc00e000;
    inBuf[1050] = 256'he400da00be00a00096009e00c400150181010a02ae025303f5038d0403055905;
    inBuf[1051] = 256'h91059c058b0564051d05c8046404e3035603bf0217027e01ff009b0071007e00;
    inBuf[1052] = 256'hb10011018701f0015702a802d502fa0214031c0332034a035a037f03ae03e003;
    inBuf[1053] = 256'h3704a7042405c6056f0603079207fc07300852085a08490856087a08af081e09;
    inBuf[1054] = 256'hac09430a010bc30b740c3a0df70d9d0e550f011093103811d1115112e5126a13;
    inBuf[1055] = 256'hcf133c148c14b014da14ee14e514fa140d1512153a1557155515671565154815;
    inBuf[1056] = 256'h50155f157415cd154316c9168f175d181719e719911afe1a641b951b8c1b911b;
    inBuf[1057] = 256'h7d1b551b611b761b911bf31b631cd41c771d061e691ecf1ef51ed11ea91e521e;
    inBuf[1058] = 256'hdd1da11d7a1d761ddc1d6c1e161f0320d7207a21122252223a220d229821ef20;
    inBuf[1059] = 256'h5f20b31ff71e6f1edb1d431de61c821c211cf71bbb1b6d1b3c1bdc1a571ae619;
    inBuf[1060] = 256'h4b199e181e188e170117ab164816eb15c2158c155c155e1548152a152515ec14;
    inBuf[1061] = 256'h91143c14ab1301136d12b9110c1191101010a80f760f340ff40ec50e600ede0d;
    inBuf[1062] = 256'h570d9b0cd70b300b7f0af0099d095209320948095c098809c709db09d309a609;
    inBuf[1063] = 256'h200964088107600639051d04f302e601f600070040ffa3fe1afec9fda1fd7efd;
    inBuf[1064] = 256'h6efd53fd0bfdaefc31fc8cfbe8fa44fa99f90df990f819f8c3f777f72ff700f7;
    inBuf[1065] = 256'hd3f6a7f697f691f698f6c4f6f6f629f765f784f78bf78df776f75cf755f744f7;
    inBuf[1066] = 256'h32f71ef7e0f682f610f67af5e4f46cf4fef3b4f391f367f342f31df3d5f287f2;
    inBuf[1067] = 256'h3df2dff18bf143f1e2f083f023f0a8ef39efe1ee8eee6fee86eebaee2eefd5ef;
    inBuf[1068] = 256'h8bf067f155f22af3fff3bff449f5bcf50ff624f623f604f6b1f55bf505f5a5f4;
    inBuf[1069] = 256'h73f46df47ff4c6f428f579f5cef50ef620f62ef636f62df641f66ff6a1f6fcf6;
    inBuf[1070] = 256'h72f7e4f76cf8f1f849f985f98ef946f9d4f83cf87bf7caf635f6b2f569f54ef5;
    inBuf[1071] = 256'h3ef54bf55df54bf528f5eaf477f4f9f37df3fbf2a4f284f284f2bef229f396f3;
    inBuf[1072] = 256'h16f49ef406f56cf5d4f524f67ff6eff64ff7bcf732f883f8c0f8e6f8cbf88bf8;
    inBuf[1073] = 256'h37f8b2f728f7b0f629f6b6f561f5f9f497f445f4d8f378f33df308f303f33ef3;
    inBuf[1074] = 256'h80f3d8f339f453f431f4d3f305f3faf1d9f08def57ee5ded79ecdaeb8beb50eb;
    inBuf[1075] = 256'h47eb6eeb7deb8beb92eb4eebe4ea64eaaae9fce884e827e825e88fe824e9fce9;
    inBuf[1076] = 256'h04ebe8ebbfec81edf3ed45ee89ee92ee9beeb5eeb2eec9ee02ef25ef62efb4ef;
    inBuf[1077] = 256'hdeef0ef042f04bf05ff085f08ff0aff0dcf0def0e2f0e2f0b3f092f085f067f0;
    inBuf[1078] = 256'h6df08df093f0a8f0bdf0a5f093f081f04bf023f000f0bcef88ef5cef1aeff6ee;
    inBuf[1079] = 256'he5eec6eec5eed1eecaeedeee03ef24ef71efdaef46f0d9f07af10df2b6f25ff3;
    inBuf[1080] = 256'hf3f396f433f5b8f546f6c7f62ef79cf7fef74cf8a5f8f7f83af98cf9d8f917fa;
    inBuf[1081] = 256'h60fa9afac0fae7fafbfa00fb13fb29fb4bfb93fbeffb61fcf3fc8bfd27feccfe;
    inBuf[1082] = 256'h63ffefff7b00f5006601d8013a029502ef0235037203ab03d503030440048604;
    inBuf[1083] = 256'heb0473050e06c7068e074a080209a909320ab30a2e0ba00b240cb60c4b0df90d;
    inBuf[1084] = 256'hb40e760f57104f1155127613941491156916f616231704179416e21521155a14;
    inBuf[1085] = 256'ha1131d13c51292129512b012cf120013241335134e1360137413af1301146a14;
    inBuf[1086] = 256'hfb148d150b167816a91694165616de154115ae141b1496133a13e8129a126212;
    inBuf[1087] = 256'h1e12cf118e114111ef10b310751042103c1050108a1003118f112112b7121b13;
    inBuf[1088] = 256'h42134113ff1292122212a0111e11b7104f10ed0fa70f580f040fb30e380e940d;
    inBuf[1089] = 256'hd70cec0bef0a100a4709ad0856081308d907a3074207c4064706c10556052305;
    inBuf[1090] = 256'h0a050f052d0530051805eb048c0415049f031e03ad0263022902120224023b02;
    inBuf[1091] = 256'h580277026d024202fb018501fb007300e4ff69ff0effbffe8bfe77fe6afe75fe;
    inBuf[1092] = 256'h98febafee5fe12ff27ff2fff29ff03ffd0fe93fe3bfedcfd74fdf3fc6bfcd8fb;
    inBuf[1093] = 256'h2bfb74faaef9d0f8f3f721f75ff6d3f57ef55af56df59cf5cbf5f9f515f620f6;
    inBuf[1094] = 256'h34f654f683f6cef61bf756f77cf776f744f7fef6a4f648f604f6d2f5b7f5bff5;
    inBuf[1095] = 256'hd9f505f647f685f6bdf6edf6fcf6f0f6d5f6a0f667f638f608f6e3f5cef5b6f5;
    inBuf[1096] = 256'ha6f5a2f59af59af5a2f59af58df579f550f52af513f504f511f538f55ef587f5;
    inBuf[1097] = 256'ha5f5a7f5a2f5a0f5a3f5c6f506f64af692f6c0f6b8f688f635f6cdf580f563f5;
    inBuf[1098] = 256'h80f5ebf595f65ff745f829f9f2f9a5fa35fb96fbd9fbf8fbf2fbe4fbd3fbcafb;
    inBuf[1099] = 256'he4fb1efc6efcd6fc37fd78fd94fd77fd1dfd9afcf2fb31fb74fabef918f995f8;
    inBuf[1100] = 256'h32f8f3f7e3f7f7f729f879f8d1f828f97cf9bef9eef913fa27fa30fa34fa30fa;
    inBuf[1101] = 256'h2ffa3dfa61faaafa25fbccfb9cfc82fd60fe1effa5ffe8ffeaffb6ff5efffafe;
    inBuf[1102] = 256'h9cfe50fe21fe0cfe0ffe29fe4ffe7cfeaefed9fefefe1fff34ff46ff59ff6aff;
    inBuf[1103] = 256'h83ffa8ffd6ff14006400ba0016016c01a701be01a7015701d90038007dffc0fe;
    inBuf[1104] = 256'h12fe74fdf9fca2fc67fc4dfc4bfc50fc59fc59fc3efc10fccffb7dfb30fbf0fa;
    inBuf[1105] = 256'hbffaaafaacfabafad9fa03fb31fb6bfbadfbeefb34fc77fcb0fceafc24fd63fd;
    inBuf[1106] = 256'haffd05fe5bfeacfee8fe03ff02ffe6febcfe98fe84fe88fea7fed8fe12ff47ff;
    inBuf[1107] = 256'h6cff77ff64ff2fffd9fe66fedefd4ffdc2fc46fce5fb9bfb67fb40fb13fbddfa;
    inBuf[1108] = 256'h9cfa4efa00fac0f98df973f976f98af9b8f902fa5cfacffa57fbd9fb51fcb0fc;
    inBuf[1109] = 256'hdbfcdffcc9fc97fc71fc67fc6bfc8bfcbdfcdbfcf4fc09fd10fd33fd86fdfefd;
    inBuf[1110] = 256'hb6fe9fff8b007c015a02fc028003e70325046804b504f6044d05b20508067506;
    inBuf[1111] = 256'hf60674071b08e208a4097e0a530bf80b8b0cfa0c2a0d520d6d0d6b0d820da80d;
    inBuf[1112] = 256'hc20dfe0d480e800ed50e320f7c0fe40f5610b4103011b01114128f1209136c13;
    inBuf[1113] = 256'hf3138d142715fa15e716cd17d118c619821a2e1ba21bc51bcf1ba71b431be51a;
    inBuf[1114] = 256'h791afb19ae197c1956197319a619d419201a581a621a6b1a4e1a021ac0196c19;
    inBuf[1115] = 256'h0419c2188918541858186c188118ba18de18d718c3187118db1732175b166315;
    inBuf[1116] = 256'h8814b413f4127b122812f7110612201234125612571234121412e011a8119811;
    inBuf[1117] = 256'h95119f11d011ff1126125c127e128e12a112941266122b12c9114d11d8105910;
    inBuf[1118] = 256'hde0f750ffb0e690ec00de80cf00bf80a040a300992081408af075707ea066306;
    inBuf[1119] = 256'hca051a056804c8033603bc025c020302b5016c011f01d10082002a00ceff6dff;
    inBuf[1120] = 256'h03ff98fe2cfebefd56fdf2fc94fc45fc04fcd5fbbcfbacfb9ffb8efb6afb35fb;
    inBuf[1121] = 256'hfcfac4faa6fab4fae5fa37fb99fbe0fbfcfbddfb75fbdafa28fa6af9c7f84cf8;
    inBuf[1122] = 256'hedf7aef780f743f7f9f699f615f680f5e6f43ff4a9f32cf3bcf270f24bf23af2;
    inBuf[1123] = 256'h50f289f2cff22df39af3f7f34df493f4b2f4c1f4c6f4b5f4acf4aff4a5f49cf4;
    inBuf[1124] = 256'h88f449f4f5f393f319f3b3f272f24af253f282f2aef2dcf2fdf2eef2caf29af2;
    inBuf[1125] = 256'h52f21af202f2f9f11df272f2d7f25ef3fdf38af40ef57ff5b4f5c1f5adf564f5;
    inBuf[1126] = 256'h0cf5bbf462f423f407f4ebf3dff3e0f3c2f39bf370f328f3e4f2b6f285f26bf2;
    inBuf[1127] = 256'h71f26ff278f290f292f29bf2bcf2dcf21cf38ef30ff4b0f472f51ef6baf642f7;
    inBuf[1128] = 256'h84f794f785f739f7d9f688f62bf6e8f5d4f5c5f5cff5f9f50cf616f61df6ebf5;
    inBuf[1129] = 256'h96f52ef590f4e1f344f39bf210f2b8f166f12bf10ff1dcf0a9f08bf05df045f0;
    inBuf[1130] = 256'h59f069f089f0baf0c0f0aef095f04af0f9efc0ef79ef45ef34ef13effaeef9ee;
    inBuf[1131] = 256'he2eed6eee6eee2eee3eeeeeeceee9eee74ee30ee03ee12ee40eeb4ee76ef4af0;
    inBuf[1132] = 256'h33f122f2cef244f389f376f33ef300f3acf270f25df248f243f249f226f2f2f1;
    inBuf[1133] = 256'hb7f157f1f9f0acf04df0f5efa4ef30efb8ee47eec9ed6ded47ed41ed7aededed;
    inBuf[1134] = 256'h6eee0aefb3ef3ff0c0f031f173f19ff1b6f1a2f185f169f145f140f165f1a6f1;
    inBuf[1135] = 256'h1bf2b9f25ff312f4b9f434f58ff5c3f5c9f5c6f5c3f5c9f5f6f547f6b0f637f7;
    inBuf[1136] = 256'hc7f74df8d0f844f9a5f905fa5efaaefa04fb56fba5fb04fc6efcebfc88fd33fe;
    inBuf[1137] = 256'he5fe95ff26009000d800f6000301180137017701da014602b502140344034c03;
    inBuf[1138] = 256'h3103f302b90299029602cd023b03c3036a041705a9052e069906df061f075907;
    inBuf[1139] = 256'h8407bf07030842089b0804097209050ab10a620b330c060dc00d760e0c0f6e0f;
    inBuf[1140] = 256'hc10ff70f0c102f1055107610ba1008115011b71123128612091391130d149d14;
    inBuf[1141] = 256'h1b156f15b815d415b81596155b150815d314a6147a147d149114ab14f8145215;
    inBuf[1142] = 256'hac1528169a16ec1640176d17681762173a17f016b51667160016b1155515ed14;
    inBuf[1143] = 256'ha914681425140b14ed13be13a413751330130813e012c112df1211135213be13;
    inBuf[1144] = 256'h19144f147c146b142014d0136413f512be129e129812c312e012db12c7127212;
    inBuf[1145] = 256'he5115311a110e80f560fc20e330ec00d3a0da50c210c8a0bf10a780afd098d09;
    inBuf[1146] = 256'h49090c09e808fc0826097409fa09870a1c0bbe0b370c890cc20cbd0c920c5f0c;
    inBuf[1147] = 256'h100cc50b970b670b440b310b000bb90a5f0ad60937099b08f3076307fd06aa06;
    inBuf[1148] = 256'h7d06770673067b06860670064506020693051805a1043004ed03e20300045104;
    inBuf[1149] = 256'hbb0410054c054f0502057d04c103d602e601f40003002fff6cfeb4fd1cfd98fc;
    inBuf[1150] = 256'h25fcd9fba2fb7afb6efb61fb48fb31fb03fbc2fa88fa4bfa16fa02faf9f9f9f9;
    inBuf[1151] = 256'h08fa02fae1f9b4f964f906f9b9f874f84bf851f863f883f8aff8bef8b8f8aaf8;
    inBuf[1152] = 256'h7ef84ef830f810f8fef702f8faf7f0f7e9f7c7f79ef77df748f715f7ecf6abf6;
    inBuf[1153] = 256'h60f611f69ef520f5a8f422f4b1f368f32ef31af331f34cf377f3aff3cdf3e0f3;
    inBuf[1154] = 256'heff3dbf3c3f3b6f3a0f3a5f3d1f30bf464f4d9f43df594f5d8f5e0f5c3f58ef5;
    inBuf[1155] = 256'h33f5d8f493f455f43af44bf469f4a5f401f55af5c0f534f691f6e6f635f75bf7;
    inBuf[1156] = 256'h6ef778f765f753f757f75ef783f7cff71ef879f8dcf81bf943f95df950f93af9;
    inBuf[1157] = 256'h36f92bf931f94ef956f94af928f9cbf845f8b2f704f765f6f5f5a2f580f597f5;
    inBuf[1158] = 256'hbcf5f1f538f666f688f6adf6b7f6bdf6d3f6ddf6f0f620f749f780f7d0f713f8;
    inBuf[1159] = 256'h56f8a3f8cdf8e5f8f5f8dbf8b2f894f86af856f86ff893f8d3f82ef971f9a0f9;
    inBuf[1160] = 256'hbcf99bf959f909f997f828f8d1f775f72ef701f7c4f68cf65bf609f6b1f55bf5;
    inBuf[1161] = 256'hecf487f43df4f6f3d8f3e5f3f9f325f459f467f462f445f4faf3aff373f33ff3;
    inBuf[1162] = 256'h3ff374f3c0f335f4b7f41cf570f59af583f54ff5fff494f445f416f407f43df4;
    inBuf[1163] = 256'ha1f41bf5b5f547f6baf61ff75df772f784f783f776f780f78bf799f7c6f7f4f7;
    inBuf[1164] = 256'h23f86bf8a6f8d7f811f92df935f942f934f924f92ff938f958f9a5f9f8f962fa;
    inBuf[1165] = 256'hebfa63fbdcfb5cfcb5fc06fd5bfd8cfdc1fd05fe30fe6afebdfefdfe5affdbff;
    inBuf[1166] = 256'h59000301db01b102aa03b904a00582064e07d1073f089708b908ef083b097f09;
    inBuf[1167] = 256'hfc09a30a440b130cf20cae0d810e550f0410d210ac1169124b133114ed14bf15;
    inBuf[1168] = 256'h82160d17a7172e188018e6183b195c198f19ad1998199a199019631966197319;
    inBuf[1169] = 256'h7819c119201a791a0b1b9c1b0a1c941c021d401d9b1de61d181e801eed1e4c1f;
    inBuf[1170] = 256'hde1f5f20b72020215d2162217621662135212a211321ec20f720f920ed201221;
    inBuf[1171] = 256'h2a213221632179216f21782154210321c1205920d71f791f0a1f911e3f1ed81d;
    inBuf[1172] = 256'h5d1dfb1c761cd61b491b981acd1915193b184f177d169615ad14f0132e137a12;
    inBuf[1173] = 256'hf91177110211b6105d10ff0fb40f470fc60e4f0ebb0d280dbb0c560c130c0c0c;
    inBuf[1174] = 256'h150c360c760c9d0caf0cb20c780c110c900bd90a090a3e0964089c07f8065b06;
    inBuf[1175] = 256'hd6056605e6045f04d20325037402ca011c0185000f00a5ff59ff28fffafedbfe;
    inBuf[1176] = 256'hc5fea0fe7afe48fef6fd93fd1afd7ffcddfb32fb7bfad4f935f99af814f895f7;
    inBuf[1177] = 256'h16f7a7f63bf6d0f57bf530f5f3f4d5f4c5f4c2f4d7f4eef406f52df551f579f5;
    inBuf[1178] = 256'hb7f5f9f542f6a0f6f1f634f76df779f75cf722f7b6f62bf69cf5fdf469f4f9f3;
    inBuf[1179] = 256'h99f356f338f314f3ebf2bbf25af2d9f14af19ef0f9ef7cef14efdceeddeee9ee;
    inBuf[1180] = 256'h06ef30ef33ef1feffeeeb0ee56ee06eea6ed58ed2cedfdece4ece9ece0ece1ec;
    inBuf[1181] = 256'hf4ecebece7eceeecd9eccaecccecb7ecb2ecc9ecd6ecfdec47ed85edd4ed36ee;
    inBuf[1182] = 256'h76eeb7eefeee25ef59efa8efe8ef41f0aff0f9f036f161f144f10bf1c8f05ff0;
    inBuf[1183] = 256'h0cf0e4efc3efceef02f01df039f04cf01ff0dfef9aef2fefdceeb1ee8cee9bee;
    inBuf[1184] = 256'he1ee27ef8eef0df069f0c6f022f14ef178f1a9f1b8f1d8f10ef22df261f2aaf2;
    inBuf[1185] = 256'hd9f218f367f39cf3dff332f467f4a3f4e6f401f51df53cf534f532f53af524f5;
    inBuf[1186] = 256'h1cf527f51ef52ff560f589f5d4f53cf691f6eff64cf773f787f785f74bf708f7;
    inBuf[1187] = 256'hc9f676f641f631f625f63df673f694f6b7f6cff6aff678f62ff6bbf54df5f5f4;
    inBuf[1188] = 256'h9ff473f473f475f48ff4b3f4b0f49cf472f414f4aaf341f3c8f26ef23ef21bf2;
    inBuf[1189] = 256'h21f248f261f27ef293f27ff262f246f21bf209f219f231f267f2b1f2e6f215f3;
    inBuf[1190] = 256'h36f32af30ef3e9f2a8f26ff244f211f2f2f1e2f1c7f1b3f1a0f175f147f116f1;
    inBuf[1191] = 256'hcff08df052f00ff0dfefbfef9def91ef93ef8fef98efa3ef9cef99ef92ef80ef;
    inBuf[1192] = 256'h81ef98efc2ef19f095f021f1c3f15ef2d7f236f36ef37df384f389f39af3d7f3;
    inBuf[1193] = 256'h39f4b9f461f512f6bbf65ff7e4f749f8a1f8e1f819f962f9b0f90efa87fa04fb;
    inBuf[1194] = 256'h86fb16fc9afc21fdb9fd50fefafebeff840055013202fb02c10389043c05f405;
    inBuf[1195] = 256'hb90671073408fe08af095f0a0b0b980b2a0cc00c400dcb0d5a0ec80e340f920f;
    inBuf[1196] = 256'hc40ff80f2b104e1099100a11881140121b13ed13d814bc1573162c17d7175f18;
    inBuf[1197] = 256'h0519ba19681a461b341c0c1dfb1dd91e851f3720ce203721b32121226c22d222;
    inBuf[1198] = 256'h2a235c23a823e523022445248424b1240b256325a32508265c268c26d6260527;
    inBuf[1199] = 256'h0c272c272f270b270127d92688265026f62574250c258724e1236123ca221c22;
    inBuf[1200] = 256'h9621f9204320b31f0a1f4c1ebb1d171d671ce41b4a1b9e1a181a7919cf185a18;
    inBuf[1201] = 256'he017721748171c17f016ed16c41678163616bd151f159914f1134513ca124312;
    inBuf[1202] = 256'hc41174110b1195103510a40ff70e570e8c0db50c000c360b750ae1093e09a408;
    inBuf[1203] = 256'h3008a7072107ba063706b3054405b3041a048f03e1022f029201dd003400aeff;
    inBuf[1204] = 256'h23ffb3fe70fe2dfe03fefbfde2fdcefdc6fda0fd79fd5efd2dfd09fdfafce1fc;
    inBuf[1205] = 256'hdbfceafceffc03fd26fd38fd4efd63fd56fd3cfd13fdc1fc65fc02fc8cfb23fb;
    inBuf[1206] = 256'hcafa74fa3dfa1ffa0bfa12fa2bfa41fa63fa83fa92faa2faa9fa9ffa9cfa97fa;
    inBuf[1207] = 256'h8cfa8ffa95fa98faa8fab6fabcfac7fac6fab6faa1fa79fa3ffa04fabef974f9;
    inBuf[1208] = 256'h3bf909f9e5f8dff8e8f804f939f974f9b2f9f5f926fa45fa59fa52fa3dfa2afa;
    inBuf[1209] = 256'h10fa01fa09fa17fa34fa64fa8dfab5fae0faf5fa01fb07fbf3fad4fab1fa7bfa;
    inBuf[1210] = 256'h48fa23fa01faf5f905fa17fa30fa49fa3dfa14fad0f95ff9dff866f8ecf792f7;
    inBuf[1211] = 256'h64f746f747f75ef765f768f765f743f71df7fff6d5f6bdf6bdf6b9f6c5f6e1f6;
    inBuf[1212] = 256'hfaf626f759f779f79ef7cff7f0f71bf84ef86bf884f89bf892f884f878f85ef8;
    inBuf[1213] = 256'h4ef855f85af86df892f8a9f8bff8d8f8daf8d3f8cdf8aef886f865f832f802f8;
    inBuf[1214] = 256'he6f7c8f7b8f7c6f7d0f7def7f9f7fbf7eaf7daf7aff777f74ef720f7fdf6faf6;
    inBuf[1215] = 256'hf7f6f9f613f719f713f71bf70ff7fcf609f718f736f77ef7c3f706f85af890f8;
    inBuf[1216] = 256'habf8cdf8d1f8cbf8e8f806f935f997f9f8f95ffae5fa4efb9dfbeffb10fc10fc;
    inBuf[1217] = 256'h12fcecfbb9fba0fb71fb49fb4cfb3cfb2bfb35fb1cfbf5fad9fa92fa3efafaf9;
    inBuf[1218] = 256'h96f936f9f9f8abf86ef858f82df809f8f5f7bbf782f75ef721f7fbf6fbf6edf6;
    inBuf[1219] = 256'hf5f616f716f712f707f7c7f680f638f6d7f597f57bf562f582f5cdf50bf66ef6;
    inBuf[1220] = 256'hc9f6eff61af71cf7e5f6b2f671f616f6dff5c6f5b2f5caf5f9f52cf67ef6cef6;
    inBuf[1221] = 256'h11f75cf78bf798f79ff782f74ef72ff714f711f74ef7b3f748f814f9e9f9c3fa;
    inBuf[1222] = 256'h97fb37fcb7fc1dfd4efd76fdadfde5fd46fed7fe79ff42002001ed01c5029403;
    inBuf[1223] = 256'h3a04e1047905ed056d06e4064607c5074808c1086609170ac60aa40b850c570d;
    inBuf[1224] = 256'h3e0e090fac0f5710da103711a71100124b12c3123713ad135814fb149b156516;
    inBuf[1225] = 256'h1517b2176418ea184e19be19fd19251a6b1a931ac11a251b7c1be01b761cf11c;
    inBuf[1226] = 256'h611de11d241e491e731e651e4d1e561e461e471e7d1e9d1eca1e161f361f4c1f;
    inBuf[1227] = 256'h6c1f531f2d1f141fce1e891e601e151ed51daf1d631d171dd91c6a1cf71b911b;
    inBuf[1228] = 256'h071b881a201a9a192019bc183218a91728177416ba15071526144f138f12b311;
    inBuf[1229] = 256'hf3105510a00f020f7b0ecd0d260d860cb60bed0a330a56099408f10734079506;
    inBuf[1230] = 256'h0e066405ce0442048d03e8024e028d01e200460087ffe4fe58feb4fd31fdc0fc;
    inBuf[1231] = 256'h35fcc4fb5bfbc9fa45fac0f913f97df8f2f74ff7cff663f6ecf596f549f5e3f4;
    inBuf[1232] = 256'h91f438f4c0f360f309f3abf279f261f24ff260f26df263f25ff23ff200f2c7f1;
    inBuf[1233] = 256'h82f137f10ef1eef0d3f0d2f0cdf0c8f0d0f0c7f0b4f0adf096f07bf06ef053f0;
    inBuf[1234] = 256'h39f02ff01ef018f02af036f04ff081f0a4f0c7f0eff0f7f0f6f0fbf0ecf0ecf0;
    inBuf[1235] = 256'h08f121f155f1a6f1e7f12cf27af2a3f2bef2daf2d9f2def2f8f205f32cf35ff3;
    inBuf[1236] = 256'h7ff3acf3d0f3c8f3b2f394f34bf307f3dbf29ff27ef288f288f299f2bbf2b7f2;
    inBuf[1237] = 256'haaf2a2f270f23cf21af2e1f1b9f1aff194f185f18df177f162f159f130f108f1;
    inBuf[1238] = 256'hf1f0b9f082f05af011f0c6ef88ef30efdfeea6ee5cee21ee03eed4edb1eda2ed;
    inBuf[1239] = 256'h74ed42ed19edd1ec8eec60ec24ecfeebfdebf5eb01ec28ec3bec53ec71ec74ec;
    inBuf[1240] = 256'h73ec79ec6cec62ec66ec57ec58ec6cec6fec8becc8ecf8ec3fed99edd4ed0fee;
    inBuf[1241] = 256'h47ee52ee56ee5dee4aee4dee6cee83eebdee18ef67efc9ef30f070f0aff0e7f0;
    inBuf[1242] = 256'hfaf018f147f167f1a3f1f6f13df296f2f3f234f380f3d5f316f46cf4ccf415f5;
    inBuf[1243] = 256'h61f5a6f5c0f5ccf5c8f5a8f597f598f59ef5caf516f65ff6b5f60af73ff769f7;
    inBuf[1244] = 256'h82f77bf777f77df77df793f7bff7eef72cf874f8aef8e9f824f94af96ff99bf9;
    inBuf[1245] = 256'hb9f9dff90ffa36fa61fa96fac3faf8fa34fb63fb93fbc7fbebfb0cfc28fc2cfc;
    inBuf[1246] = 256'h28fc20fc07fceafbcefbabfb91fb83fb73fb73fb83fb94fbaefbc8fbd2fbd8fb;
    inBuf[1247] = 256'hd6fbc3fbadfb97fb82fb80fb8dfba5fbcdfbf5fb0ffc1ffc18fcf7fbc8fb89fb;
    inBuf[1248] = 256'h46fb0cfbd8fab1fa9efa8ffa84fa80fa77fa72fa7afa83fa9afac4faf3fa31fb;
    inBuf[1249] = 256'h80fbcffb2cfc96fcfefc77fdfcfd79fefdfe82fff1ff5f00ce002c0194010802;
    inBuf[1250] = 256'h7b020803a3033304cd046205d00537069506d6062a079007f70789083709da09;
    inBuf[1251] = 256'h920a430bc90b540cd20c2a0d9c0d1b0e880e1d0fc10f4c10f3109f113012e612;
    inBuf[1252] = 256'ha813561435152016e816ca179b183219db19751ae61a841b311cd21cb21d9c1e;
    inBuf[1253] = 256'h621f43200621862117228d22d5224e23cc233224d3246f25dc256426ca26f926;
    inBuf[1254] = 256'h4d279427c2273328a72802298f29fc29272a5e2a632a2e2a232a0f2aef291e2a;
    inBuf[1255] = 256'h532a782acc2af72ae62ae22aa52a302adf297329f528b6286b280b28db278d27;
    inBuf[1256] = 256'h1527b72637269d253025a324ff238323e02220228521c620fb1f5f1fa91ef11d;
    inBuf[1257] = 256'h6b1dca1c201c981be41a1c1a6f199618b317f5161b1643158f14b813d9120b12;
    inBuf[1258] = 256'h0e110610120ff90dea0c020c050b160a4509550863077c067005670473036a02;
    inBuf[1259] = 256'h7601a100c1fff6fe3ffe71fdadfcf5fb2afb73fad4f932f9aaf836f8b9f747f7;
    inBuf[1260] = 256'hcff63af6a6f50cf567f4dbf367f304f3cbf2a9f290f287f271f245f20ff2bef1;
    inBuf[1261] = 256'h5cf103f1aff071f05ef061f082f0c5f006f145f17ef196f19af193f16ff14cf1;
    inBuf[1262] = 256'h32f10ef1fcf001f100f110f130f145f167f191f1a8f1caf1f2f105f221f240f2;
    inBuf[1263] = 256'h47f259f272f27af294f2bff2e4f225f37df3ccf329f488f4cdf414f556f57ef5;
    inBuf[1264] = 256'hb7f5fff53bf68ef6f4f64ef7b8f72af888f8eff857f9a7f9f9f944fa6bfa89fa;
    inBuf[1265] = 256'h9afa86fa6efa58fa32fa20fa28fa2ffa4cfa7afa95faa9faaffa89fa50fa0cfa;
    inBuf[1266] = 256'hacf955f913f9d1f8acf8a7f89af892f88bf866f837f805f8b9f76bf72af7dcf6;
    inBuf[1267] = 256'h98f664f61df6d7f59ef556f51df5fff4e1f4d9f4f0f4fff40df518f5fbf4c6f4;
    inBuf[1268] = 256'h87f428f4d0f398f36df36cf39df3d2f311f451f464f457f431f4d9f374f318f3;
    inBuf[1269] = 256'hb2f264f237f206f2e7f1d8f1b4f196f183f15bf13ef132f116f102f1f2f0c1f0;
    inBuf[1270] = 256'h8bf054f003f0c7efaaef90ef9fefd4ef03f03cf072f07af073f063f035f018f0;
    inBuf[1271] = 256'h18f018f03df07ef0aef0e6f01df12df140f15bf160f17cf1b1f1d9f111f24ef2;
    inBuf[1272] = 256'h67f27cf28ff283f288f2a7f2c3f204f369f3c1f323f483f4b5f4daf4f7f4f3f4;
    inBuf[1273] = 256'hf9f416f529f552f58cf5aef5d1f5f2f5f2f5f5f504f605f618f640f658f671f6;
    inBuf[1274] = 256'h8bf68bf68af694f697f6b5f6f9f647f7b1f72ff896f8eff833f946f93ef92af9;
    inBuf[1275] = 256'h00f9e0f8d9f8def8fdf836f96ff9acf9e7f908fa1ffa2ffa2bfa25fa25fa23fa;
    inBuf[1276] = 256'h2bfa42fa5ffa8cfac4fafdfa3ffb82fbbbfbf1fb1efc39fc48fc45fc31fc13fc;
    inBuf[1277] = 256'he6fbb0fb7dfb49fb24fb18fb1afb34fb68fba0fbe1fb25fc52fc72fc88fc8bfc;
    inBuf[1278] = 256'h98fcbbfcecfc4efde4fd92fe66ff4d001e01e50194020f037b03dd0329049004;
    inBuf[1279] = 256'h13059a054b061807dd07b9089a095b0a230be50b820c270dc90d4c0ee40e850f;
    inBuf[1280] = 256'h1410c61086113012f512ba135a140715a7151c16a0161f17811703188818f118;
    inBuf[1281] = 256'h7819f719501abc1a1a1b551bb11b101c611ce01c621dc81d451ea31eca1ef51e;
    inBuf[1282] = 256'hff1ee91e001f231f521fcb1f5920e32092211f227822cf22f322ea22fc22fe22;
    inBuf[1283] = 256'hf82225234b2363239423992372235123fc2283221d229521fa207a20dc1f2f1f;
    inBuf[1284] = 256'h9d1eef1d391da61cfa1b491bb21af51923195c1866176216771578148913cc12;
    inBuf[1285] = 256'h0c126211db1038108c0fe20e040e160d2f0c2b0b360a68099808e9075c07c306;
    inBuf[1286] = 256'h3706b3050a055d04aa03d202f7011c0126003aff59fe6efd9dfcdffb20fb7bfa;
    inBuf[1287] = 256'hdef931f98bf8d8f708f738f65ff578f4abf3ebf238f2abf12df1b9f05ff001f0;
    inBuf[1288] = 256'ha0ef4feff2ee93ee47eef2ed9bed53edfbeca1ec53ecf6eb9deb5aeb11ebd9ea;
    inBuf[1289] = 256'hc0eaa5ea9feab6eac4eaddea02eb0aeb0deb0cebe9eac6eaadea8aea86eaabea;
    inBuf[1290] = 256'hd8ea2deba1eb08ec77ece3ec22ed59ed87ed98edbdedfded40eeb1ee49efdeef;
    inBuf[1291] = 256'h8ff04bf1e7f185f21cf38df302f476f4c8f420f574f5a4f5d8f50ef62bf65ef6;
    inBuf[1292] = 256'ha7f6edf654f7d1f73bf8abf80ff942f964f977f965f960f971f981f9b4f904fa;
    inBuf[1293] = 256'h49fa96fadefafdfa11fb1efb0cfb03fb08fb01fb07fb1dfb1dfb22fb2cfb1ffb;
    inBuf[1294] = 256'h14fb12fbfbfae7fad9faaffa83fa5cfa1cfae0f9b5f97ef951f938f90bf9d8f8;
    inBuf[1295] = 256'ha4f849f8ddf770f7eaf66df610f6b8f57cf563f541f51df5fbf4b2f456f4f9f3;
    inBuf[1296] = 256'h82f30cf3b3f259f210f2e0f19ff15bf120f1cef07ef046f00cf0e9efe7efe0ef;
    inBuf[1297] = 256'he0efe5efcaefa3ef7eef45ef1eef1fef30ef6aefd0ef36f0a6f014f15cf18ff1;
    inBuf[1298] = 256'hb0f1adf1a6f1a6f19df1a9f1cff1f6f135f286f2ccf218f360f38bf3aff3c7f3;
    inBuf[1299] = 256'hc4f3caf3daf3e9f319f463f4b0f414f579f5c6f50af638f644f64ff65bf668f6;
    inBuf[1300] = 256'h9bf6eef653f7ddf770f8f4f871f9d4f911fa44fa69fa85fab8fafbfa46fbaafb;
    inBuf[1301] = 256'h10fc68fcbffc02fd2cfd52fd6dfd7ffd9bfdb7fdcdfdecfd03fe10fe23fe33fe;
    inBuf[1302] = 256'h44fe67fe95fec8fe09ff46ff77ff9fffb4ffb5ffb1ffa5ff97ff96ff99ffa1ff;
    inBuf[1303] = 256'hb3ffc4ffd3ffe5fff6ff080021003a0053006a00760077006e0058003f002c00;
    inBuf[1304] = 256'h200025003a0056007800930099008c006b003300faffc7ff9eff90ff9bffb1ff;
    inBuf[1305] = 256'hd9ff04002300440062007a00a400de001f017701da0130028b02de021f036b03;
    inBuf[1306] = 256'hc3031d049b042d05b8055206dd063f079607d807fb0732087c08cc084b09e309;
    inBuf[1307] = 256'h720a160baf0b1e0c920cfa0c430da70d150e6f0ee90e630fbb0f28109110e010;
    inBuf[1308] = 256'h5a11e81170122e13f7139d145315eb153f169616d916f9164e17c0173918fe18;
    inBuf[1309] = 256'hdd19a81a961b6a1cfc1c931d051e3f1e971eea1e251f991f142079201121a221;
    inBuf[1310] = 256'h1222ac22332391230b2464248324af24b0247a2463243a240024072415241c24;
    inBuf[1311] = 256'h5b2483247e2485245024dc237123dd223022b4213321b52076202c20d81faa1f;
    inBuf[1312] = 256'h5d1ff81eac1e3a1eaf1d3d1da21cf21b5a1ba11ae3195019b1182118c4175717;
    inBuf[1313] = 256'he6168216e71525155514461323121411f40ff30e280e600db10c1a0c590b830a;
    inBuf[1314] = 256'h990972083a070606c0049b039f02ac01e0002e006dffb8fe03fe32fd6afca6fb;
    inBuf[1315] = 256'hd1fa12fa59f997f8ecf746f799f607f67df5f1f481f413f49cf335f3c2f23df2;
    inBuf[1316] = 256'hc3f139f1a5f028f0a5ef27efc7ee65ee09eec7ed7eed3aed0cedd1ec96ec67ec;
    inBuf[1317] = 256'h1deccaeb7ceb12ebabea5dea0eeadfe9dfe9e8e910ea52ea81eaafeadbeadfea;
    inBuf[1318] = 256'hdceae0eaceead5eaffea2eeb86eb03ec7bec06ed98ed06ee70eed1ee0bef47ef;
    inBuf[1319] = 256'h87efafefe9ef34f072f0c9f035f196f10bf28bf2f2f25ef3c4f303f43ff476f4;
    inBuf[1320] = 256'h8ff4b3f4e4f408f543f58ef5ccf519f66bf6a5f6e5f625f74af777f7aaf7c9f7;
    inBuf[1321] = 256'hf5f72cf856f88ef8d5f812f95ef9b9f906fa5dfab9fafafa38fb70fb8afb9efb;
    inBuf[1322] = 256'hb3fbb2fbb6fbc3fbc2fbc7fbd5fbd1fbd1fbd7fbcbfbc2fbc0fbacfb99fb88fb;
    inBuf[1323] = 256'h60fb2ffbfafaacfa5bfa14fac9f993f97ef974f97ef997f99af989f961f90af9;
    inBuf[1324] = 256'h99f826f8adf74ef71ff70df724f75ef793f7c1f7e2f7d9f7b6f788f745f70af7;
    inBuf[1325] = 256'he5f6c8f6c4f6d7f6e8f6fef617f71df720f725f71af710f70af7f5f6ddf6c5f6;
    inBuf[1326] = 256'h9bf673f651f62cf615f60ef607f60af614f611f60df609f6f9f5eff5edf5eaf5;
    inBuf[1327] = 256'hf4f508f616f62df649f65bf677f69cf6c1f6f4f631f765f798f7c1f7d2f7d9f7;
    inBuf[1328] = 256'hdaf7d3f7dff701f832f87bf8cdf80df93cf94bf92ff9fcf8bff882f865f870f8;
    inBuf[1329] = 256'h9df8f1f857f9b2f9fbf923fa1cfafcf9cef9a1f991f9a9f9e7f94ffacffa4efb;
    inBuf[1330] = 256'hc6fb22fc55fc6efc6efc5efc56fc61fc82fcc2fc19fd7dfdecfd55feacfef8fe;
    inBuf[1331] = 256'h31ff56ff77ff94ffb1ffdcff120051009c00e7002c0169019201a601af01aa01;
    inBuf[1332] = 256'ha001a001a901c001e5010d023502570267026e02730275028c02c1020d037603;
    inBuf[1333] = 256'hf3036b04dd0438056f059605b605d3050e066e06e5067d072408b3082f098709;
    inBuf[1334] = 256'haa09b909bd09ba09d9091c0a700ae50a610bbe0b0b0c340c2a0c170c010ce60b;
    inBuf[1335] = 256'hf30b220c5b0cb60c140d530d8e0dae0da40da10d9f0d970dba0df90d400eb00e;
    inBuf[1336] = 256'h2c0f960f12108010cd1027117811b51117128612f61295134114e01492152b16;
    inBuf[1337] = 256'h9116ed161f172117301739173e177a17ca1718188618db18f9180219cd185b18;
    inBuf[1338] = 256'hf0177e171717fa16051728177a17b517bb17a5174717ac1616167915f614c314;
    inBuf[1339] = 256'hb914d01414153f153a151915af1412147513ce124112f911d211cd11f111fa11;
    inBuf[1340] = 256'hde11a61126117810c10ff30e350ea80d2d0dd20c9b0c540c000c9c0b010b470a;
    inBuf[1341] = 256'h7c098e08a607d70611066f05f20478040a049a0305035f02a801d4000b0056ff;
    inBuf[1342] = 256'haefe33fed8fd83fd41fdf6fc89fc0dfc76fbc5fa21fa8af903f9aef875f847f8;
    inBuf[1343] = 256'h2cf8fcf7a1f72ef78ef6cdf517f567f4d4f37ff349f329f322f300f3b8f256f2;
    inBuf[1344] = 256'hbff108f15cf0b2ef2aefe3eebfeec3eef1ee10ef1eef1befdeee7bee0fee8ded;
    inBuf[1345] = 256'h1dede0ecc2ecdbec30ed8aedeeed4bee6cee61ee38eedced7ded3eed14ed29ed;
    inBuf[1346] = 256'h85edf8ed8dee2def9aefe1efffefd7ef97ef5eef20ef0def31ef67efbdef22f0;
    inBuf[1347] = 256'h5ef080f084f04af003f0c3ef7eef62ef77ef9defe3ef38f06ef09bf0b6f0a8f0;
    inBuf[1348] = 256'h9ff0abf0bcf0fdf06ff1eff18cf234f3baf333f495f4c9f4f7f429f550f591f5;
    inBuf[1349] = 256'hedf547f6b5f62cf788f7e0f72ef856f875f88cf885f87df877f85ef852f855f8;
    inBuf[1350] = 256'h51f85ff87cf88cf8a0f8b2f8a7f896f883f85ef844f83bf832f83ef85df873f8;
    inBuf[1351] = 256'h90f8b1f8bef8cef8e5f8f4f812f942f96ff9a8f9e7f911fa32fa47fa3dfa2bfa;
    inBuf[1352] = 256'h19fafbf9eaf9e9f9e5f9e9f9f2f9e5f9d0f9b6f983f94ff91ef9dbf898f855f8;
    inBuf[1353] = 256'hf8f795f732f7c3f662f61bf6e2f5c7f5c6f5bef5b4f59cf559f5fdf494f41af4;
    inBuf[1354] = 256'hb3f374f359f375f3c4f329f49ff414f567f59ef5baf5aff59af58cf583f595f5;
    inBuf[1355] = 256'hc5f506f663f6cdf62bf786f7d4f702f81ff82df824f81bf816f811f81ef838f8;
    inBuf[1356] = 256'h52f879f8a2f8bef8dcf8f4f801f916f931f94bf973f9a0f9c6f9edf90afa14fa;
    inBuf[1357] = 256'h1cfa1cfa18fa28fa4afa7efacffa31fb99fb05fc5efc9dfccbfcddfcddfce2fc;
    inBuf[1358] = 256'hedfc0efd51fdaafd16fe91fefefe5bffa6ffd2ffecff0500170039007300b300;
    inBuf[1359] = 256'h02015c01a601e8012102410262028a02b102f0024803a2030a047604c7040f05;
    inBuf[1360] = 256'h490568059005c70506066f06fd06980750080c09ab09410aba0a030b430b790b;
    inBuf[1361] = 256'ha00be50b420ca60c320dcb0d500edc0e4e0f890fb40fbc0f970f7e0f660f490f;
    inBuf[1362] = 256'h5f0f910fc90f2c109310dc102a11571151114b113011fe10f61004111b116f11;
    inBuf[1363] = 256'hda114012c6123d138c13e51324143e147414a714ce1423158015d1154616b016;
    inBuf[1364] = 256'hfb165b17a317ca170818391852188b18b618c418e918f118cf18bc188e184018;
    inBuf[1365] = 256'h1218da1796177f176117321727170617c4169c165d160716d915aa157c158915;
    inBuf[1366] = 256'h9e15b415fc153b166616ac16d416dc16f516ef16cf16cb16bc16a616bd16d316;
    inBuf[1367] = 256'he7161f173f173e1740171217b5165a16da154a15dc146d140914d513a0136913;
    inBuf[1368] = 256'h471303139c122d128b11c9100c10390f690ec60d2f0db40c6c0c2a0cf20bcc0b;
    inBuf[1369] = 256'h890b2e0bcf0a460aa90916097808ea0788073707080708071007260748075007;
    inBuf[1370] = 256'h46072d07e9068c062306a1051c05a3042904c403790333030003d50297024e02;
    inBuf[1371] = 256'hea015a01ae00e7ff05ff29fe59fd9bfc09fc9bfb47fb15fbecfab9fa84fa38fa;
    inBuf[1372] = 256'hd1f961f9e4f860f8eef785f727f7e4f6acf680f66cf65ef658f666f670f676f6;
    inBuf[1373] = 256'h80f670f64af61cf6d5f588f546f508f5e3f4e2f4ebf407f536f552f563f56af5;
    inBuf[1374] = 256'h52f52bf503f5c9f496f472f446f423f410f4f0f3dbf3d6f3cbf3cff3e9f3fdf3;
    inBuf[1375] = 256'h1af43df445f443f439f410f4e8f3d0f3bbf3caf306f454f4bff43bf5a3f5fef5;
    inBuf[1376] = 256'h4cf672f685f691f686f681f68bf68ef6a2f6c3f6daf6fcf628f745f767f78cf7;
    inBuf[1377] = 256'h9af7a0f79bf775f745f711f7c9f690f674f665f67cf6b8f6fbf651f7abf7e5f7;
    inBuf[1378] = 256'h0ff829f820f814f811f80cf822f855f88bf8d5f82bf96ff9b0f9f1f91cfa46fa;
    inBuf[1379] = 256'h72fa8efaa9fac3fac3fabefab5fa96fa79fa6cfa5cfa59fa68fa6dfa71fa6dfa;
    inBuf[1380] = 256'h46fa0afabef954f9eaf88df82df8e5f7b7f788f761f73ff709f7d2f69ff65ff6;
    inBuf[1381] = 256'h31f619f601f6fcf509f609f60ef619f615f618f625f629f638f64ff655f65cf6;
    inBuf[1382] = 256'h65f65af651f652f64cf655f66ff680f699f6b1f6aaf694f66ef628f6e1f5a4f5;
    inBuf[1383] = 256'h6af551f55cf573f5a1f5d6f5f2f5fef5f2f5bdf57af531f5ddf4a1f482f473f4;
    inBuf[1384] = 256'h8df4c5f40af568f5cdf524f67df6c9f6f7f61ef73af744f75df784f7b5f70bf8;
    inBuf[1385] = 256'h7af8f4f884f916fa92fa03fb59fb8afba9fbb5fbaefbaffbb7fbc4fbe7fb15fc;
    inBuf[1386] = 256'h44fc7efcb3fcdefc0dfd38fd5bfd85fdadfdccfde8fdf7fdfbfd00fe01fe09fe;
    inBuf[1387] = 256'h29fe5cfea7fe0eff80fff7ff6f00d400260165018c01a801c701e70118026102;
    inBuf[1388] = 256'hb50219038603ec034d04a504ed0432057105a705e0051906460672069806b306;
    inBuf[1389] = 256'hcf06eb06060731076707a207f10747089708ea082d0957097409730954092d09;
    inBuf[1390] = 256'hfb08c808ad08a508b508ee0839098709df091f0a390a3a0a100abf096a091209;
    inBuf[1391] = 256'hc408a508ab08d3082a098a09e0092d0a530a490a270ae5098f0948090709d008;
    inBuf[1392] = 256'hb808aa089e08a308a108950895088f088208860885087f0885087f086a085908;
    inBuf[1393] = 256'h3e081e08130810081b084a088508c1080d094c0973099309990989097a095f09;
    inBuf[1394] = 256'h400934092a09230936094a095b0977098b09900995098709680948091809dd08;
    inBuf[1395] = 256'hab08730836080908db07ac0787075f0735071007e406b6068f0660062e060006;
    inBuf[1396] = 256'hca058c054f050a05c5048a0452042a0417040d0411042004280427041b04f703;
    inBuf[1397] = 256'hc60388033c03f302af027002430222020602f701ea01d201b30183013b01e500;
    inBuf[1398] = 256'h7900f7ff73ffe5fe51feccfd50fddffc87fc3bfcf9fbc6fb8afb42fbf5fa8efa;
    inBuf[1399] = 256'h13fa99f914f992f82af8cef78af76bf758f756f76bf776f778f779f759f724f7;
    inBuf[1400] = 256'he8f68ff62df6daf583f53bf515f5f7f4eef401f50bf513f51ff50bf5e5f4b9f4;
    inBuf[1401] = 256'h71f423f4e4f39df367f34df332f329f335f336f340f355f356f358f361f351f3;
    inBuf[1402] = 256'h3ef32df302f3daf2bdf293f27cf27df279f28cf2b4f2ccf2ecf215f328f33ff3;
    inBuf[1403] = 256'h5af35ff36af37cf377f379f384f37ef387f3a1f3b3f3dcf31df455f49bf4e9f4;
    inBuf[1404] = 256'h1cf549f569f564f559f54cf52cf520f52af535f55af597f5ccf50df655f689f6;
    inBuf[1405] = 256'hbff6f1f604f712f71af701f7e7f6d0f6adf69df6a6f6b4f6e3f62cf771f7c4f7;
    inBuf[1406] = 256'h16f849f86ff882f870f856f83df81af810f823f83df873f8c1f808f956f9a5f9;
    inBuf[1407] = 256'hdbf90bfa36fa45fa4bfa4bfa32fa17fa01fae1f9d4f9e3f9fef936fa89fadefa;
    inBuf[1408] = 256'h38fb8cfbc1fbe0fbeafbcefba6fb7efb50fb36fb39fb4bfb79fbbbfbf8fb38fc;
    inBuf[1409] = 256'h6efc85fc89fc80fc5cfc30fc02fccafb9cfb7afb58fb46fb47fb4afb57fb69fb;
    inBuf[1410] = 256'h6dfb6bfb62fb43fb20fbfffad9fabffab2faa6faa2faa3fa9afa8ffa83fa72fa;
    inBuf[1411] = 256'h6afa72fa87fab2faf0fa35fb7dfbbbfbe2fbf6fbf6fbe7fbdafbd9fbf1fb28fc;
    inBuf[1412] = 256'h7bfce5fc60fdd9fd45fea1fee3fe0eff26ff2cff2aff29ff27ff2fff45ff63ff;
    inBuf[1413] = 256'h90ffcdff0e0052009600ca00f10007010201ec00cc00a1007d00680062007900;
    inBuf[1414] = 256'hac00ee004701ac0108026002ad02e3020e032c03370347035c036f039a03da03;
    inBuf[1415] = 256'h23048b0405057d05fc057006c306070732073a07450751075a078307c2070608;
    inBuf[1416] = 256'h6708d1082d099109ee09340a820aca0afe0a420b830bac0be00b0d0c210c400c;
    inBuf[1417] = 256'h5f0c700c9e0cd90c100d670dc50d120e6e0ebb0ee40e0f0f260f1a0f1c0f1a0f;
    inBuf[1418] = 256'h0b0f210f460f710fcd0f37109c1022119b11ed113f126e1267125d123b120112;
    inBuf[1419] = 256'heb11e311e2111f127312c7124213b4130014501479146f1467144214fc13d513;
    inBuf[1420] = 256'hb11388139513b513dc133a149e14f2145e15a915bc15c21594152c15cc145f14;
    inBuf[1421] = 256'hec13b813a413a913ef133e148114d514ff14f114dc149c143414e01385132813;
    inBuf[1422] = 256'hfd12de12c712e112fa120b133b135913571362134c130f13d71281121612cc11;
    inBuf[1423] = 256'h821143113b1140114b1173118611781168113011d7108b103610e40fbb0f9c0f;
    inBuf[1424] = 256'h830f870f790f540f310fed0e900e400ee50d8d0d540d1d0dec0cce0ca00c640c;
    inBuf[1425] = 256'h2d0cdb0b750b160ba50a2f0ac8095909f208a90866083408230815080c080a08;
    inBuf[1426] = 256'hee07bb0776070d078f0616069a053305f304cd04cc04ec040f0532054b054105;
    inBuf[1427] = 256'h1705d0046604ec036e03ec027d022602df01b401a30199019c019c0187016201;
    inBuf[1428] = 256'h1d01ab001f0078ffbafe06fe5ffdcefc6afc25fcf8fbe5fbd2fbacfb7afb28fb;
    inBuf[1429] = 256'hb2fa2ffa9bf900f97af802f89df75df72ff711f70af702f7f9f6fbf6f0f6ddf6;
    inBuf[1430] = 256'hcdf6aef686f660f62af6eff5bef584f550f531f512f501f506f508f510f524f5;
    inBuf[1431] = 256'h20f50ff5f6f4b7f466f412f4a7f343f3fdf2c2f2acf2c3f2e1f212f354f377f3;
    inBuf[1432] = 256'h86f384f354f315f3d8f288f24bf231f21ef228f252f276f2a7f2e5f209f32ef3;
    inBuf[1433] = 256'h59f369f37af392f38ef38ef396f38bf38ff3aaf3c3f3fcf353f4a3f403f56bf5;
    inBuf[1434] = 256'hadf5ddf5fbf5e8f5cbf5a9f573f553f551f54ff570f5b0f5e5f529f674f69ff6;
    inBuf[1435] = 256'hc3f6daf6cbf6b5f69cf66bf64af643f63bf657f695f6d2f61ff774f7a7f7c8f7;
    inBuf[1436] = 256'hd4f7b1f782f74ef709f7dbf6cdf6c5f6d9f605f725f745f760f75ef756f74cf7;
    inBuf[1437] = 256'h2ff71cf714f7fff6f4f6f1f6dff6d3f6d3f6cdf6d6f6f1f607f728f74af753f7;
    inBuf[1438] = 256'h4ff73df70bf7d4f6a6f678f666f679f69cf6d5f61df752f777f787f76df73ef7;
    inBuf[1439] = 256'h0af7caf69bf68ff695f6b7f6f6f634f770f7a3f7b4f7acf792f75bf71bf7e4f6;
    inBuf[1440] = 256'hb0f692f694f6a6f6cdf606f737f75ff77bf778f760f73af702f7cdf6a8f68ef6;
    inBuf[1441] = 256'h91f6b4f6e9f633f789f7d6f71ef858f876f884f888f87df877f87ef88ff8baf8;
    inBuf[1442] = 256'h00f953f9b9f926fa86fadcfa20fb42fb50fb4ffb41fb38fb3efb51fb7dfbbffb;
    inBuf[1443] = 256'h09fc5bfcaafce6fc13fd2cfd2ffd27fd1afd0bfd07fd12fd2bfd58fd92fdd2fd;
    inBuf[1444] = 256'h1afe61fea2feddfe0bff2eff4eff68ff83ffa9ffdaff1d007500d5003a01a101;
    inBuf[1445] = 256'hf8013f0275029402a802bd02d302f7022f037103bf030f044e047c0497049504;
    inBuf[1446] = 256'h860473045f045b0467047e04a104c704e104f504fb04f004e504da04cd04cc04;
    inBuf[1447] = 256'hd104d604e204eb04ee04f604fc0404051a05360555057f05a405bc05d005d605;
    inBuf[1448] = 256'hd005ce05cd05d305f005170644067d06ad06cd06e306e306cb06ae0686065a06;
    inBuf[1449] = 256'h39061e06080603060006fe0508060b060506fd05e505b70580053805e804a204;
    inBuf[1450] = 256'h65043f043d0451047804af04dc04f204ef04c20472041404aa0348030403de02;
    inBuf[1451] = 256'hdd02ff022b0358037e03830367033403e5028a023202e0019f0177015d015501;
    inBuf[1452] = 256'h5e01640169016c015d0143011c01e400a60064001c00ddffabff82ff6dff66ff;
    inBuf[1453] = 256'h63ff67ff65ff52ff36ff0affd1fe9afe65fe35fe18fe07fef9fdf5fdedfddbfd;
    inBuf[1454] = 256'hc3fd9efd6dfd3efd0cfddbfcb6fc95fc76fc64fc4efc33fc1bfcf7fbcafb9dfb;
    inBuf[1455] = 256'h60fb1bfbd9fa91fa4dfa1dfaf6f9e1f9e7f9f2f9fff90efa05fae7f9bcf974f9;
    inBuf[1456] = 256'h22f9daf892f85df84cf84bf85ff88cf8b0f8ccf8e4f8daf8b7f88cf843f8f3f7;
    inBuf[1457] = 256'haff766f72bf70ff7fcf6fff620f73df761f78bf797f78cf76ff727f7ccf66ef6;
    inBuf[1458] = 256'h03f6abf579f559f55ef587f5aef5dbf505f608f6f6f5d2f58bf541f5fff4b8f4;
    inBuf[1459] = 256'h89f477f46bf479f4a0f4c2f4f3f42af54bf568f57df56df552f531f5f9f4ccf4;
    inBuf[1460] = 256'hb1f497f49bf4bdf4ddf407f533f53cf533f51bf5e2f4a9f47ef455f448f458f4;
    inBuf[1461] = 256'h66f47df496f492f482f46bf441f422f41bf41df43cf474f4a7f4dcf409f513f5;
    inBuf[1462] = 256'h0ef501f5e1f4cff4d4f4e1f40bf54bf584f5c3f500f624f647f66af67ff69ef6;
    inBuf[1463] = 256'hc7f6e5f607f729f738f74af760f770f792f7caf706f853f8a8f8e8f81bf93cf9;
    inBuf[1464] = 256'h38f925f90ff9f2f8e9f8f8f813f947f98ef9ccf90afa45fa6efa90faaefabffa;
    inBuf[1465] = 256'hd2fae8faf5fa08fb21fb38fb5efb96fbd8fb2efc91fcf2fc4cfd90fdaffdb3fd;
    inBuf[1466] = 256'h9bfd6ffd4bfd3cfd47fd7cfdd2fd38fea4fefdfe34ff4cff41ff1efffcfee6fe;
    inBuf[1467] = 256'he4fe06ff42ff91ffecff3e008400be00e300fd0017012e014b0172019901c601;
    inBuf[1468] = 256'hf701220252028702b902f3022f035e038903a803ae03ad03a903a303b603e003;
    inBuf[1469] = 256'h18046c04cb0417055a05820583057a056a0552055a058105b90515067e06da06;
    inBuf[1470] = 256'h3a078907b407dc07fc070b082a0855087d08bd0803093f098c09da091a0a6f0a;
    inBuf[1471] = 256'hc80a150b6e0bbe0bf20b240c430c460c570c6b0c7c0cb10cf60c380d8f0dde0d;
    inBuf[1472] = 256'h120e480e670e660e6d0e690e520e510e4d0e3f0e4b0e570e5e0e860eb20ed70e;
    inBuf[1473] = 256'h140f4a0f670f8a0f920f790f6d0f590f3d0f4b0f690f920fe40f36107510bc10;
    inBuf[1474] = 256'he810ed10f410e810ca10c810c510bb10d110e210e010f110f510e910f6100011;
    inBuf[1475] = 256'hfe1016111f110e110711e710ad1088105f103610351039103b105a1067105710;
    inBuf[1476] = 256'h50103010f70fd50fae0f860f830f7e0f6f0f780f6e0f4d0f400f290f090f0e0f;
    inBuf[1477] = 256'h170f1d0f3d0f4b0f410f420f290ffa0ee70ed30ec00ed40ee60eeb0eff0ef80e;
    inBuf[1478] = 256'hd00eb00e7d0e3f0e250e0f0efb0d060e050eeb0dd60da70d5b0d200de10ca40c;
    inBuf[1479] = 256'h910c870c7d0c8f0c930c7f0c730c530c1f0c040ce80bcb0bd10bd50bcf0bdc0b;
    inBuf[1480] = 256'hda0bca0bcf0bd10bd40bfb0b210c3d0c640c6e0c540c360cff0bbd0b9c0b8a0b;
    inBuf[1481] = 256'h8d0bbb0bed0b140c3b0c3a0c0e0cd80b880b2f0bf30ac60aac0ab60ac10ac20a;
    inBuf[1482] = 256'hc40aa90a750a440a0b0ad609be09ab099e09a009900969093d09fe08b6087f08;
    inBuf[1483] = 256'h51083608390840084808530846082208f907c0077e0746070b07d606aa067406;
    inBuf[1484] = 256'h3c060706c505840552052005f404d204a5046e042904c9035d03ed0276021002;
    inBuf[1485] = 256'hc401870164015501440137012101f700c400890042000400c8ff82ff43fffffe;
    inBuf[1486] = 256'haefe62fe16fecffda1fd84fd70fd6dfd60fd3bfd01fd9efc14fc7dfbd7fa38fa;
    inBuf[1487] = 256'hbdf95ef923f912f909f900f9f4f8c5f878f818f896f707f783f6fdf584f52af5;
    inBuf[1488] = 256'hd9f49cf47cf45af442f440f434f426f421f405f4ddf3b9f380f346f322f3fcf2;
    inBuf[1489] = 256'heaf2fef218f341f380f3aef3d5f3fbf302f4fdf3fbf3def3bcf3a6f37af34ff3;
    inBuf[1490] = 256'h32f309f3edf2ecf2e5f2eef20cf314f31af31df3f7f2c5f293f246f207f2e5f1;
    inBuf[1491] = 256'hc0f1b8f1d1f1e1f101f22af233f23ff250f243f240f24df247f252f269f268f2;
    inBuf[1492] = 256'h6ff27ef274f279f291f29cf2bef2f1f211f336f35af35df35ff360f347f339f3;
    inBuf[1493] = 256'h38f328f325f32cf323f321f323f313f30ef317f317f327f344f352f364f371f3;
    inBuf[1494] = 256'h64f353f341f321f313f321f33bf37bf3daf33cf4aef422f57bf5cdf512f639f6;
    inBuf[1495] = 256'h60f68cf6aef6e4f62cf773f7d1f73ff8a4f813f981f9d4f91dfa52fa5bfa50fa;
    inBuf[1496] = 256'h34fafef9d1f9b2f996f998f9b2f9d0f9f9f91bfa21fa17faf6f9b2f968f922f9;
    inBuf[1497] = 256'hddf8b1f8a3f8a6f8c2f8e8f805f91df929f91ef909f9f1f8d5f8c4f8c1f8c8f8;
    inBuf[1498] = 256'hdef801f926f955f98af9b8f9e3f909fa22fa31fa32fa26fa1dfa1bfa1efa37fa;
    inBuf[1499] = 256'h6afaa9faf5fa43fb7ffba6fbaefb8efb56fb11fbc6fa93fa82fa91faccfa2afb;
    inBuf[1500] = 256'h93fb00fc62fca5fcd0fce2fcddfcd7fcd9fce6fc10fd53fda4fd09fe7cfef0fe;
    inBuf[1501] = 256'h67ffdaff3e009600d900010113010e01f300cf00ac00900088009500b400e600;
    inBuf[1502] = 256'h1e014f0172017b0166013601f0009c004a000200cdffb1ffadffbbffd8fffcff;
    inBuf[1503] = 256'h23004a006e008a009f00ab00b000ae00a700a400aa00bd00e2001b016101b201;
    inBuf[1504] = 256'h07025902a402e40217034003610377038c039e03a703a803a30394037e036703;
    inBuf[1505] = 256'h510349034e035c0374038e039c03970378033b03e80287022202cd0195017b01;
    inBuf[1506] = 256'h8301a501d601100244026a0284028e02860276025f02420225020902f301ea01;
    inBuf[1507] = 256'hed01fd011e024b027b02aa02ca02d102c0028f023f02dd0172010801b0006f00;
    inBuf[1508] = 256'h490043004f0064007c008b00890076004c001200d2ff8dff48ff0cffe0fec7fe;
    inBuf[1509] = 256'hc8fee1fe0dff4bff91ffd3ff0c003100410042003500220018001d0032005b00;
    inBuf[1510] = 256'h9400d7001a0156018801ad01c301ce01d001ca01be01ad019601770149011001;
    inBuf[1511] = 256'hd000890042000200c7ff90ff5fff2bfff1feb1fe67fe16fec7fd77fd2dfdedfc;
    inBuf[1512] = 256'hb1fc7dfc52fc2afc07fcf3fbedfbf6fb15fc3ffc70fca4fccafcdffce2fccffc;
    inBuf[1513] = 256'haefc8dfc70fc63fc74fc9cfcdafc2cfd82fdd3fd15fe3cfe4bfe46fe2cfe05fe;
    inBuf[1514] = 256'hdffdb8fd9afd8efd8ffda2fdc8fdf8fd2ffe66fe8bfe9cfe96fe6cfe2afedefd;
    inBuf[1515] = 256'h89fd43fd1bfd0cfd20fd54fd90fdd1fd0afe25fe2cfe1ffef7fdccfda8fd88fd;
    inBuf[1516] = 256'h7bfd7ffd87fd97fdaafdadfdaafda0fd85fd65fd41fd12fde4fcb5fc7afc3efc;
    inBuf[1517] = 256'h05fcc8fb90fb62fb35fb11fbeffac4fa96fa67fa2ffafdf9d7f9bdf9b8f9c6f9;
    inBuf[1518] = 256'hdef9fef91ffa35fa40fa40fa34fa2bfa2cfa34fa4efa7dfabafa06fb59fba8fb;
    inBuf[1519] = 256'hfbfb49fc89fcc3fcf4fc15fd2efd3dfd3cfd3cfd3efd41fd58fd86fdc2fd13fe;
    inBuf[1520] = 256'h6cfeb4fee9fefefee1fe9efe3dfec5fd58fd04fdccfcc5fcebfc2dfd83fdd9fd;
    inBuf[1521] = 256'h19fe3ffe43fe1efedffd91fd39fdeefcbdfca9fcbafcecfc38fd96fdf9fd55fe;
    inBuf[1522] = 256'ha3fed9fef3fef2fed9feb3fe88fe61fe4bfe4afe5cfe81feb3feeafe23ff58ff;
    inBuf[1523] = 256'h83ffa6ffc1ffd0ffd4ffd1ffbfffa1ff7bff4eff26ff0eff09ff22ff5cffadff;
    inBuf[1524] = 256'h0d007400ca00040123011e01fc00cd009e0081008600ab00f3005f01d8015602;
    inBuf[1525] = 256'hd2023b039103d303fb03150425042b04300438043f04500469048304a804d504;
    inBuf[1526] = 256'h0305380568058805a305ab059705770548050805cd0494045f04450440044b04;
    inBuf[1527] = 256'h7904bc0406056205ba05fd05360654064e063e0622060006f705080634069106;
    inBuf[1528] = 256'h1107a2074c08f4088109f609410a570a4e0a290aed09bf09a2099a09c0090a0a;
    inBuf[1529] = 256'h6a0ae50a620bc70b160c380c1e0cda0b6e0be00a570adb0978094d094e096b09;
    inBuf[1530] = 256'had09f309200a3c0a2f0af509aa094909df0893085d083d084d087308a008e008;
    inBuf[1531] = 256'h150936095809660963096f0978097e099709ab09b309c309c009a90998097a09;
    inBuf[1532] = 256'h5409420932092509350949095a0977098309770965093909f208af0866082208;
    inBuf[1533] = 256'hfc07e907ec0715084a088008c408f908140923091809f408cd089d086c085308;
    inBuf[1534] = 256'h450846086c089f08d80826097009ab09de09f209e509c40982092709cf087108;
    inBuf[1535] = 256'h1c08eb07ce07c407da07f207ff070608e807a6074c07d0064206c1054605e104;
    inBuf[1536] = 256'ha804870480049704b004c604e004e404d704c804a904870471045c0454046304;
    inBuf[1537] = 256'h73048604a804c204d304e804f50403051805280538054e05570553054a052c05;
    inBuf[1538] = 256'hfc04c9048b0449041204e503c903c303c603ce03d903d303b8038c034703f102;
    inBuf[1539] = 256'h97023b02e701a70177015b015701600175019601b301ca01db01dc01d201bf01;
    inBuf[1540] = 256'h9f017c015c013c0125011e012201380160018f01c401f701170223021702e801;
    inBuf[1541] = 256'ha0014801e30082003000edffc6ffb9ffbfffd5fff1ff01000100eaffb1ff61ff;
    inBuf[1542] = 256'hfdfe90fe2bfed7fd9bfd7ffd84fd9efdc9fdfbfd28fe4bfe59fe51fe37fe0ffe;
    inBuf[1543] = 256'hddfdacfd82fd65fd59fd5afd65fd79fd8dfd9ffdaafda8fd99fd80fd58fd27fd;
    inBuf[1544] = 256'hf6fcc0fc8dfc62fc3bfc18fcfcfbdcfbbcfb9afb6dfb3efb12fbe4fabbfa9dfa;
    inBuf[1545] = 256'h83fa6efa61fa4ffa3bfa26fa0afaeaf9d0f9b8f9acf9b5f9cbf9f3f92ffa71fa;
    inBuf[1546] = 256'hb4faf8fa30fb59fb76fb7ffb7afb72fb66fb62fb6cfb85fbb1fbf0fb36fc7efc;
    inBuf[1547] = 256'hc6fcfdfc20fd2dfd20fd01fdd4fc9cfc6cfc49fc34fc37fc54fc80fcb9fcfbfc;
    inBuf[1548] = 256'h31fd5afd6ffd67fd48fd16fdcffc86fc46fc0cfcebfbedfb06fc3afc83fcc9fc;
    inBuf[1549] = 256'h05fd31fd35fd19fde6fc95fc39fce5fb97fb64fb57fb63fb8cfbcefb0ffc44fc;
    inBuf[1550] = 256'h6cfc71fc55fc22fcd4fb7bfb2cfbe5fab3faa3faadfad0fa0bfb4dfb8ffbcefb;
    inBuf[1551] = 256'hf8fb0dfc10fcfcfbdefbc5fbb1fbaefbc2fbe6fb19fc5bfc9afcd4fc09fd2cfd;
    inBuf[1552] = 256'h41fd50fd4efd47fd45fd40fd3ffd46fd46fd48fd4bfd41fd37fd34fd2afd27fd;
    inBuf[1553] = 256'h30fd33fd39fd40fd36fd22fd08fdd8fca1fc6afc26fcecfbc6fba3fb91fb98fb;
    inBuf[1554] = 256'ha2fbb4fbc9fbc8fbb9fb9cfb64fb1efbd7fa8bfa4cfa26fa0ffa12fa32fa58fa;
    inBuf[1555] = 256'h83faaffac8fad0fac8faaafa83fa5cfa33fa15fa0afa08fa17fa39fa60fa8efa;
    inBuf[1556] = 256'hc2faeffa1afb40fb57fb65fb68fb5bfb4cfb3ffb2ffb2ffb43fb65fb9dfbe8fb;
    inBuf[1557] = 256'h33fc82fccafcf7fc12fd18fd00fde1fcbffc99fc84fc86fc93fcb8fcedfc22fd;
    inBuf[1558] = 256'h5cfd94fdb6fdcffdd9fdcefdbcfda4fd82fd69fd59fd4efd55fd69fd84fdadfd;
    inBuf[1559] = 256'hdffd10fe45fe76fe9bfebafec8fec4feb5fe9cfe79fe58fe3dfe30fe3bfe5cfe;
    inBuf[1560] = 256'h92fedffe36ff88ffcaffedffedffcaff86ff30ffdcfe97fe70fe74fea2fef4fe;
    inBuf[1561] = 256'h63ffdbff4a00a200d600e200ca0094004d000700ccffa8ffa8ffc9ff06005d00;
    inBuf[1562] = 256'hc3002a018c01de01120228021c02f201b40167011b01e400c800ca00f1003601;
    inBuf[1563] = 256'h8b01e4013002650277025c021902b9014101c3004e00eeffabff8cff90ffafff;
    inBuf[1564] = 256'hdeff110040005d005b003e000400b3ff54fff6fea6fe70fe58fe62fe8dfed0fe;
    inBuf[1565] = 256'h22ff78ffc5ff06003600510058004e0037001a00fbffdfffd0ffd2ffe7ff1600;
    inBuf[1566] = 256'h5d00b40014017201c101f7010502eb01b0015b01fe00aa006d0053005e008600;
    inBuf[1567] = 256'hc40007013e015c0156012c01e6008b002900d1ff8fff67ff59ff60ff76ff92ff;
    inBuf[1568] = 256'ha8ffb1ffb1ffa6ff92ff7dff6bff5fff59ff59ff5aff57ff4dff38ff19fff2fe;
    inBuf[1569] = 256'hc6fe9dfe81fe73fe77fe8efeb2fedafefcfe0dff05ffe5feadfe65fe1cfedefd;
    inBuf[1570] = 256'hb4fdaafdbdfdedfd33fe80fec9fe06ff2cff3aff36ff23ff0bfff7feebfeecfe;
    inBuf[1571] = 256'hfafe10ff33ff5fff91ffcdff110057009e00e100150136013a012001f400b700;
    inBuf[1572] = 256'h73003c001b0014002d005f009e00e00014012b012401f4009f003500c0ff48ff;
    inBuf[1573] = 256'hdffe90fe5efe4dfe58fe78fea8fedafe00ff18ff1dff0affe0fea6fe62fe1efe;
    inBuf[1574] = 256'he4fdbafda6fdacfdcbfd00fe46fe90fed8fe17ff46ff60ff62ff4cff22ffecfe;
    inBuf[1575] = 256'haffe77fe4efe3dfe49fe74feb7fe0fff6fffc8ff0f00380040002800f3ffadff;
    inBuf[1576] = 256'h69ff30ff0bff07ff20ff54ff9ffff4ff48009600d100f50006010201e900c400;
    inBuf[1577] = 256'h9600630035001000f7fff9ff16004b009500ed0043018b01b501b80194014901;
    inBuf[1578] = 256'hdf006a00f8ff96ff51ff34ff3cff61ff97ffd2ff050020001900f2ffb2ff5dff;
    inBuf[1579] = 256'hfefea2fe55fe1ffe02fe00fe1afe48fe85fecbfe11ff50ff86ffaaffc1ffcbff;
    inBuf[1580] = 256'hc6ffb8ffa8ff97ff8aff87ff8effa6ffd2ff0f005f00c10029018f01e9012b02;
    inBuf[1581] = 256'h4e024e022802e8019d0152011a01060119015801be013902b70224036c038203;
    inBuf[1582] = 256'h6403110399020c027c010001a60077007a00a800f5005601b9010b0241024f02;
    inBuf[1583] = 256'h3102ec01890111019a003300ebffd2ffe6ff23008300f8006c01d10117023302;
    inBuf[1584] = 256'h2602f00199013701d10073003300180021005300ab001b01990113027c02cb02;
    inBuf[1585] = 256'hf202e902bf0278021a02bf017901510158019001ef016a02ed026103bf03f303;
    inBuf[1586] = 256'hf303cc0387032b03cf028102480232023f026802ac0201035c03ba030b044304;
    inBuf[1587] = 256'h690473045b042d04ee03a3035f032803030301031c034d039603e0031a044504;
    inBuf[1588] = 256'h50043304fe03b30359030403b8027c025f025d027002a102df021e0362039a03;
    inBuf[1589] = 256'hb803c403b6038e035c032103e702c302b002af02ca02f3021f034f0377039003;
    inBuf[1590] = 256'ha103a5039e039a0394038d038e038e038a038a03880386039103a303bf03ea03;
    inBuf[1591] = 256'h190444046d0485048604780457042704f703c8039f0387037b0375037c038603;
    inBuf[1592] = 256'h8d039b03a703ae03bb03c203be03b903a803870362033a031103f702e902eb02;
    inBuf[1593] = 256'h0b03370366039c03c803df03e503d103a4036c032703dc02a0026d0249024102;
    inBuf[1594] = 256'h4c0267029602c602f4021d03300327030a03d20289024002fa01c601b201b601;
    inBuf[1595] = 256'hd4010d024c028a02c202e502ef02e802cb029c0265022702eb01bd0199018801;
    inBuf[1596] = 256'h9401b501e80130027d02c002f5020d030203d7028e023402de0192015d014e01;
    inBuf[1597] = 256'h5c017f01b201e40104020f02fe01d5019d0159011301d5009a0066003f001f00;
    inBuf[1598] = 256'h0700feff02001500370063009500c900f00008010e01fd00da00af0080005a00;
    inBuf[1599] = 256'h47004b006a00a100e50031017a01b701de01ec01dc01b40177012d01df009c00;
    inBuf[1600] = 256'h6f005d0068008e00c300fd002d01460143012201e40091003600ddff8fff51ff;
    inBuf[1601] = 256'h24ff07fff8feedfee5fee0fed9fed4fed2fed2fed3fecdfebafe98fe68fe2afe;
    inBuf[1602] = 256'heafdb3fd8ffd89fda1fdd6fd20fe72febefef2fe06fff8fecefe8dfe44fe01fe;
    inBuf[1603] = 256'hd1fdbcfdc5fde6fd1cfe5afe99fed1fefafe11ff17ff0ffffcfee5feccfeb7fe;
    inBuf[1604] = 256'hacfeacfebafed3fef3fe1aff44ff6bff8dffa8ffb8ffc0ffc2ffbcffb5ffa9ff;
    inBuf[1605] = 256'h98ff88ff77ff67ff5fff5fff6aff83ffa6ffccfff2ff0a000e00ffffd7ff9bff;
    inBuf[1606] = 256'h57ff15ffe1fec2feb9fec7fee6fe08ff21ff2eff29ff0fffe5feb6fe8cfe6ffe;
    inBuf[1607] = 256'h61fe61fe6efe83fe9afeadfebdfec7fecdfed2fed4fed6fed9fedcfeddfedffe;
    inBuf[1608] = 256'he0fee2fee4fee5fee9fef0fef4fef7fefafefbfefbfefefe01ff0dff22ff3aff;
    inBuf[1609] = 256'h54ff6dff7dff85ff83ff76ff66ff59ff4dff48ff4cff55ff63ff70ff76ff79ff;
    inBuf[1610] = 256'h79ff70ff67ff63ff5dff59ff58ff55ff53ff4fff47ff41ff42ff46ff51ff64ff;
    inBuf[1611] = 256'h78ff8aff99ff9cff92ff7fff62ff3eff18fff0fecafeacfe90fe7bfe6ffe63fe;
    inBuf[1612] = 256'h5bfe59fe54fe50fe4bfe3efe29fe0bfee1fdb5fd8dfd68fd55fd59fd6dfd92fd;
    inBuf[1613] = 256'hc0fde6fd02fe0efe03fee5fdb9fd84fd57fd3afd27fd28fd3dfd5bfd7efd9ffd;
    inBuf[1614] = 256'hb6fdc6fdd0fdd0fdcefdd1fdd5fddffdeefdfdfd0ffe24fe36fe46fe57fe64fe;
    inBuf[1615] = 256'h72fe81fe8afe91fe98fe9afe99fe95fe89fe78fe62fe42fe1ffefefdddfdc3fd;
    inBuf[1616] = 256'hb9fdb9fdc5fddcfdf4fd08fe13fe0afef2fdcefda0fd74fd55fd42fd43fd5afd;
    inBuf[1617] = 256'h7cfda4fdcdfde9fdf6fdf3fddafdb9fd96fd6ffd51fd42fd3bfd41fd54fd68fd;
    inBuf[1618] = 256'h82fda1fdbbfdd4fdeffd00fe0ffe1afe1bfe19fe1afe18fe1bfe28fe35fe47fe;
    inBuf[1619] = 256'h5ffe6ffe79fe7dfe71fe5dfe44fe1efef5fdcffda5fd82fd6bfd55fd47fd44fd;
    inBuf[1620] = 256'h44fd4afd55fd5afd5dfd5cfd50fd3efd29fd0efdfbfcf3fcf3fcfefc14fd28fd;
    inBuf[1621] = 256'h3cfd46fd3dfd25fd03fdd6fcaafc86fc69fc60fc6bfc7dfc97fcb6fccbfcd9fc;
    inBuf[1622] = 256'he1fcdbfcd1fcc9fcc0fcc2fcd0fce0fcf8fc17fd2ffd41fd50fd4ffd44fd33fd;
    inBuf[1623] = 256'h18fdfcfce4fcc8fcb2fca6fc97fc8cfc89fc82fc7bfc7afc75fc70fc74fc77fc;
    inBuf[1624] = 256'h81fc94fca4fcb5fcc6fcc9fcc5fcbefcabfc98fc8cfc83fc85fc94fca2fcb2fc;
    inBuf[1625] = 256'hc1fcc0fcb4fc99fc6afc39fc0cfce3fbccfbcffbe5fb0ffc46fc79fcacfcd2fc;
    inBuf[1626] = 256'hdefcdafccafcaafc88fc6efc5afc58fc69fc84fcacfcdafc01fd21fd35fd34fd;
    inBuf[1627] = 256'h27fd12fdeffccdfcb3fca1fc9cfcabfcc6fceefc1dfd46fd6dfd8efd9efda3fd;
    inBuf[1628] = 256'ha4fd9dfd94fd8ffd8afd8dfd97fda3fdb5fdccfdddfdeefd01fe0efe1bfe28fe;
    inBuf[1629] = 256'h31fe3bfe46fe4cfe53fe5cfe64fe72fe84fe97feb1fed3fef3fe13ff34ff54ff;
    inBuf[1630] = 256'h71ff85ff90ff98ff9aff91ff86ff7dff74ff6fff6eff71ff7bff89ff95ffa2ff;
    inBuf[1631] = 256'hadffb1ffaeffa2ff8cff73ff59ff3eff28ff1eff1eff2bff40ff5bff7aff97ff;
    inBuf[1632] = 256'hadffbeffc6ffc2ffb8ffabff9fff97ff98ffa2ffb6ffd3fff9ff24004d007000;
    inBuf[1633] = 256'h8e00a300ae00b000ac00a700a500a800b300c600df00020129014a0168018101;
    inBuf[1634] = 256'h8e0191018c017e01710165015c015b015f01640170017d0185018c0190018e01;
    inBuf[1635] = 256'h8b0185017e017c017c017e018a019701a301b201c001c701d001d301d101d301;
    inBuf[1636] = 256'hd401d301db01e801f90111022602370247024e02490241023502290228022e02;
    inBuf[1637] = 256'h3b02550274029502b902d202e002e802e202d102c002ad029e029b02a102ac02;
    inBuf[1638] = 256'hc202d702e802fb0208030b030903fe02ec02e102d502c802c802d202de02f502;
    inBuf[1639] = 256'h0f0325033c034a034e0355035303460340033a033203340339033b0343034703;
    inBuf[1640] = 256'h45034803470342034a03570365037f039903ac03c403d403d603d603d003c303;
    inBuf[1641] = 256'hbf03be03c003d403ec03030421043a0445044a04400427040c04ec03c803b103;
    inBuf[1642] = 256'ha503a303b803d703fc032c0454046e04810482046e04550433040d04f403e203;
    inBuf[1643] = 256'hd803e403f8030f042c043d043d04390429040a04e903c603a3038f0382037803;
    inBuf[1644] = 256'h80039103a403c503e503ff031d0433043b043f043a042a041d040e04fd03f803;
    inBuf[1645] = 256'hfb0302041504270432043f04440439042e041f040a04fa03ed03e003e003e703;
    inBuf[1646] = 256'hed03fa0305040904120418041504160416041104110412040a040404f903e603;
    inBuf[1647] = 256'hd603c103a2038c0379036503600365036c0380039503a003a903a70395038103;
    inBuf[1648] = 256'h68034d0341033e0342035c037e039e03bf03d403d603cd03b3038b0366034503;
    inBuf[1649] = 256'h28031e031d03220332033e033e033b0330031d030c03fa02e902e602e902ef02;
    inBuf[1650] = 256'h000312031e032b0330032b03240319030b03070307030b031a032c033e035103;
    inBuf[1651] = 256'h5a03560349032f030c03e802c402a30295029802ab02ce02f7021e0341035303;
    inBuf[1652] = 256'h500340031f03f302ca02a6028c0286029102a702c902ec02070319031a030503;
    inBuf[1653] = 256'he302b10276023f021002eb01dc01e101f501190243026b028c029e029d029002;
    inBuf[1654] = 256'h76025102300219020b020d021a022f024b02620270027602700260024d023402;
    inBuf[1655] = 256'h19020202ec01d801cd01c301b801b401b301b501b901c001cc01de01eb01f201;
    inBuf[1656] = 256'hf501ef01df01ca01af0194017c0169015c01570156015c016501690169016601;
    inBuf[1657] = 256'h58013f011f01fa00d700b700a100970098009f00ae00c000cd00d400d300c800;
    inBuf[1658] = 256'hb3009700760057003b00230010000000f4ffecffe3ffd8ffceffc7ffbeffb5ff;
    inBuf[1659] = 256'haeffa5ff98ff87ff74ff63ff52ff43ff3dff3eff46ff54ff65ff75ff82ff87ff;
    inBuf[1660] = 256'h87ff81ff75ff66ff58ff4cff43ff3fff3eff3dff3fff40ff3eff3cff37ff32ff;
    inBuf[1661] = 256'h30ff2cff28ff25ff21ff18ff0dff00fff3fee7fedafed0fecdfecbfec9fecbfe;
    inBuf[1662] = 256'hcefecefecbfec3feb7fea9fe95fe7cfe66fe52fe41fe3afe38fe3bfe44fe4efe;
    inBuf[1663] = 256'h55fe58fe51fe41fe2ffe18fe01feeffde1fddcfde3fdebfdf1fdfafdfcfdf6fd;
    inBuf[1664] = 256'hecfddbfdc8fdbafdaffdaafdaffdb6fdbffdccfdcffdccfdc6fdb9fda7fd98fd;
    inBuf[1665] = 256'h8afd84fd88fd90fda0fdb4fdc1fdccfdd6fdd2fdc2fdaffd98fd82fd70fd5ffd;
    inBuf[1666] = 256'h5afd62fd6dfd7dfd91fd9cfd9efd98fd84fd68fd48fd24fd06fdf3fce6fce4fc;
    inBuf[1667] = 256'heefcf8fc05fd10fd10fd06fdf7fcdcfcbefca2fc87fc74fc6cfc67fc67fc6dfc;
    inBuf[1668] = 256'h6ffc71fc74fc70fc6bfc68fc5dfc54fc51fc4dfc4bfc4cfc4cfc4dfc50fc4bfc;
    inBuf[1669] = 256'h46fc44fc3cfc34fc2ffc27fc20fc1efc19fc16fc17fc13fc0efc0cfc03fcf9fb;
    inBuf[1670] = 256'hf4fbe9fbe3fbe5fbe6fbebfbf5fbfbfb02fc0bfc09fc04fc00fcf4fbe8fbdefb;
    inBuf[1671] = 256'hd0fbc6fbc2fbb8fbaffbadfba7fba3fba5fba3fba2fba5fb9ffb99fb93fb85fb;
    inBuf[1672] = 256'h79fb75fb6cfb68fb6bfb6ffb7dfb90fb9afba5fbb1fbb2fbaffba9fb99fb8afb;
    inBuf[1673] = 256'h80fb75fb6ffb70fb6efb74fb80fb88fb93fba1fba6fbaafbb1fbb0fbaffbb0fb;
    inBuf[1674] = 256'hadfbadfbb2fbb5fbc0fbd1fbdefbeffb04fc11fc19fc1dfc1bfc19fc14fc09fc;
    inBuf[1675] = 256'h01fcfefbf9fbf8fbfefb02fc0bfc1bfc28fc37fc49fc57fc65fc73fc7afc82fc;
    inBuf[1676] = 256'h8bfc8afc88fc8cfc8ffc96fca3fcb0fcc2fcdafcecfcfafc04fd03fdfffcf7fc;
    inBuf[1677] = 256'he3fccdfcbdfcabfc9ffc9dfc9efca9fcbdfcd2fce9fc00fd0efd17fd1bfd12fd;
    inBuf[1678] = 256'h04fdf7fce7fcdcfcddfce6fcfafc1bfd3efd64fd88fd9efdaafdadfda1fd8dfd;
    inBuf[1679] = 256'h79fd66fd59fd57fd5ffd74fd95fdb9fddffd07fe28fe41fe53fe58fe57fe53fe;
    inBuf[1680] = 256'h4cfe49fe4ffe5cfe72fe8efeadfecffeeffe03ff0cff0eff08fffcfeeefee2fe;
    inBuf[1681] = 256'hdafed8fedefeeafef9fe08ff15ff23ff2fff38ff3fff4bff5cff70ff84ff99ff;
    inBuf[1682] = 256'hacffbcffc4ffc7ffc6ffc1ffbeffbdffbcffc1ffcbffd4ffddffe6ffe9ffe7ff;
    inBuf[1683] = 256'he0ffd3ffc3ffb5ffa9ffa3ffa6ffafffc1ffdbfff8ff16003300490059006100;
    inBuf[1684] = 256'h60005d005a00570059006200710083009900ab00b900c200c400bf00b800b100;
    inBuf[1685] = 256'haf00b500c500dc00fa001a01380154016701710175017401740178017b017f01;
    inBuf[1686] = 256'h8c019e01b001c101cc01d201d001c301af019a0180016701580150014f015c01;
    inBuf[1687] = 256'h74019201b301cf01e601f601f601ea01dd01cd01c001be01c501d501f0010e02;
    inBuf[1688] = 256'h28023e02470246023f022c021302fd01ea01db01d701d801db01e401ec01f301;
    inBuf[1689] = 256'hfb01fe01fd01ff01fe01fd01020207020b0215021c021f0221021d0216021102;
    inBuf[1690] = 256'h0902000201020602100225023d0253026a0276027702710260024b023b023102;
    inBuf[1691] = 256'h330249026a029402c502f20217032f03330329031603f702d502bf02b302b302;
    inBuf[1692] = 256'hc302dc02fb021c033803490350034b033c0325030803ee02dd02d002cb02d602;
    inBuf[1693] = 256'hec02040320033b035203610363035c0355034b033b0330032a03250325032503;
    inBuf[1694] = 256'h21031f0319030f030803ff02f802f602f402ef02f102ee02e102d402c102a902;
    inBuf[1695] = 256'h97028a0284028d029d02b502d702f5020a031b031f0315030503ea02c902ad02;
    inBuf[1696] = 256'h9502870289029602b002d8020203270349035c035c034e0333031003f002d502;
    inBuf[1697] = 256'hc602cd02e10201032b03550377038f0391037f03620338030703d902b2029602;
    inBuf[1698] = 256'h880284028a029a02ab02b902c602ce02cf02c902b802a00288026e0254024102;
    inBuf[1699] = 256'h3702340238024302520263026f02740275026d025d0246022b020d02f201dd01;
    inBuf[1700] = 256'hce01c801c901d301e401fa010f0226023502390237022a021202f801de01c701;
    inBuf[1701] = 256'hbb01b601b801c401d501e401f001f301ee01e401d301bf01b001a3019b019e01;
    inBuf[1702] = 256'ha401ad01ba01c201c701cf01d201d101d301d101cd01cd01c901c201bc01b101;
    inBuf[1703] = 256'ha7019e0193018a018801850185018801890189018d0191019401970197019901;
    inBuf[1704] = 256'h990192018b0185017a017001680162015d01590154014f0148013c012e012101;
    inBuf[1705] = 256'h11010101f600ed00e500df00db00d800d500d200cd00ca00cb00ce00d200d300;
    inBuf[1706] = 256'hd300d600d500cf00c800c000b400a7009b009100890081007b007a007a007e00;
    inBuf[1707] = 256'h860090009d00ac00b700bc00ba00af009c008700710060005b00610072008e00;
    inBuf[1708] = 256'haa00c300d500d900cb00af00870056002400f7ffd7ffcbffd0ffe4ff02002500;
    inBuf[1709] = 256'h4900630068005e0047002200f5ffc7ff9eff82ff78ff7dff94ffb5ffd9fffaff;
    inBuf[1710] = 256'h110016000900ecffc4ff97ff6aff43ff2bff1eff1dff28ff36ff44ff53ff5eff;
    inBuf[1711] = 256'h62ff62ff60ff59ff52ff4aff40ff35ff2aff20ff17ff0fff0dff14ff21ff32ff;
    inBuf[1712] = 256'h4aff62ff73ff7cff7bff6dff52ff2eff09ffe7fec8feb3feaefeb4fec3fedcfe;
    inBuf[1713] = 256'hfbfe1bff36ff46ff4aff3eff22fffdfed7feb3fe95fe87fe88fe99feb4fed3fe;
    inBuf[1714] = 256'hf1fe08ff11ff0cfff6fed0fea4fe77fe4efe32fe28fe2afe38fe50fe6cfe88fe;
    inBuf[1715] = 256'ha2feb6fec5fed0fed7fedafed9fed3fecdfec7febdfeb6feb5feb6febafec5fe;
    inBuf[1716] = 256'hd1fedafee1fee3fedffed4febffea4fe8afe6dfe50fe39fe29fe22fe27fe37fe;
    inBuf[1717] = 256'h50fe70fe8ffeacfec2fecbfec9febcfea2fe7ffe60fe44fe31fe2efe39fe51fe;
    inBuf[1718] = 256'h72fe91fea9feb7feb6fea8fe91fe73fe5afe4dfe47fe4efe65fe83fea8feccfe;
    inBuf[1719] = 256'he8fe01ff14ff18ff18ff12ff04fff9fef2fee8fee5fee7fee4fee4fee5fee1fe;
    inBuf[1720] = 256'hddfed7fecbfec3febdfeb7feb9febffec5fed4fee3feeffefcfe02ff00fffffe;
    inBuf[1721] = 256'hfcfef6fef7fe00ff0cff1eff31ff3dff44ff46ff3dff2fff1eff0cfffefef3fe;
    inBuf[1722] = 256'heafee7fee6fee6fee9feecfeeffef4fefafefefe05ff0bff0eff13ff16ff12ff;
    inBuf[1723] = 256'h0cff08ff01fffbfef8fef7fefdfe09ff14ff20ff2cff30ff32ff31ff2bff27ff;
    inBuf[1724] = 256'h24ff1aff10ff08ff00ff00ff02ff07ff1bff38ff53ff6fff87ff94ff9aff96ff;
    inBuf[1725] = 256'h85ff72ff5cff45ff38ff31ff30ff3dff51ff68ff84ff9dffadffb6ffb6ffa9ff;
    inBuf[1726] = 256'h95ff78ff57ff39ff1fff0cff0bff1bff39ff65ff99ffcafff2ff0a000d00faff;
    inBuf[1727] = 256'hd5ffa8ff7aff53ff3dff3cff4cff6bff94ffbcffdcfff1fff6ffeeffd9ffb8ff;
    inBuf[1728] = 256'h92ff6fff53ff40ff36ff38ff42ff54ff6cff85ff9bffafffc0ffc8ffcaffc8ff;
    inBuf[1729] = 256'hbcffa6ff8fff7aff66ff58ff52ff54ff5dff6dff82ff9cffb7ffd2ffe7fff5ff;
    inBuf[1730] = 256'hf9ffeeffd7ffb8ff96ff77ff64ff60ff72ff9cffd2ff0d00470073008d008d00;
    inBuf[1731] = 256'h740048001400ddffb2ff9aff97ffacffd5ff07003a00680085008e0084006800;
    inBuf[1732] = 256'h46002100ffffe4ffd6ffd3ffdcffefff070020003600470050004c003f002b00;
    inBuf[1733] = 256'h1300fcffe9ffdcffd8ffdfffebfffaff0600100018001b001d00220026002b00;
    inBuf[1734] = 256'h320038003b003a003200260018000700f8fff1fff1fff9ff08001b002e003b00;
    inBuf[1735] = 256'h40003f00360028001a000e0009000b00100015001d00230028002f0034003700;
    inBuf[1736] = 256'h3900390035002c001f0012000500fafff3fff1fff3fffbff0700110019001f00;
    inBuf[1737] = 256'h240024002300230027002f0037003e00440046003f00310020000900f3ffe8ff;
    inBuf[1738] = 256'he4ffe7fff4ff02000f00180016000b00fbffe5ffcfffbdffaeffa5ffa4ffaaff;
    inBuf[1739] = 256'hb7ffc9ffdefff7ff0c00190020001f001000f7ffdbffbbff9fff89ff7bff78ff;
    inBuf[1740] = 256'h81ff92ffa6ffb9ffcaffd1ffc9ffb7ffa1ff88ff70ff60ff56ff53ff56ff5aff;
    inBuf[1741] = 256'h5eff63ff69ff70ff78ff82ff8eff96ff96ff8fff7eff61ff3fff1dfffefee7fe;
    inBuf[1742] = 256'hdffee3fef4fe0fff2dff47ff61ff73ff78ff71ff61ff4bff34ff1dff0bff01ff;
    inBuf[1743] = 256'h01ff0dff23ff3fff60ff85ffa6ffbfffcdffc9ffb2ff8dff5cff29fffffee3fe;
    inBuf[1744] = 256'hdafeeafe09ff32ff5dff7eff97ffa4ff9cff86ff6bff4aff2aff13ff01fffcfe;
    inBuf[1745] = 256'h06ff19ff35ff58ff7aff98ffadffb4ffafff9aff78ff55ff33ff12fffefef8fe;
    inBuf[1746] = 256'hfbfe0cff29ff45ff5dff6cff71ff6eff63ff55ff4eff4dff51ff5bff6aff77ff;
    inBuf[1747] = 256'h7fff7eff79ff76ff74ff74ff7cff88ff94ffa2ffadffb0ffabffa0ff8fff7aff;
    inBuf[1748] = 256'h68ff5bff59ff60ff70ff89ffaaffcdffedff08001c0028002d0029001e001200;
    inBuf[1749] = 256'h0600fdfffafffeff0d00260042005b0071007b0077006900510034001e000f00;
    inBuf[1750] = 256'h0c001a0031004d0069007e008c00940094009300960099009f00aa00b500bc00;
    inBuf[1751] = 256'hbf00bb00b000a100910083007b007c0086009500a500b100b700b700b300a800;
    inBuf[1752] = 256'h9a008f008a008d009500a100b200c200ce00da00e300e800ea00e600de00d600;
    inBuf[1753] = 256'hca00bc00b400b100b200b900c300cf00db00e000df00dd00d600d000d300da00;
    inBuf[1754] = 256'he600fb0010011f012b0130012b0123011501060100010501120125013b014f01;
    inBuf[1755] = 256'h5b015c0152013f0124010901f600ee00ef00fb000c011e01320143014a014c01;
    inBuf[1756] = 256'h4b0144013c01310124011a0112010c010e0115011d012a013a0144014a014a01;
    inBuf[1757] = 256'h43013701280117010d0106010101070113011e012801300132012f0127011c01;
    inBuf[1758] = 256'h160116011a0124012f0135013b013b0135012f012a01260128012b0131013a01;
    inBuf[1759] = 256'h4301490150015301510150014d01470143013b012f0125011f011b011e012201;
    inBuf[1760] = 256'h2c013d014e015c01670166015c014d0136011b010801fb00f600fd000b011f01;
    inBuf[1761] = 256'h3601430149014a01400132012601160107010001fa00f700fc0002010a011801;
    inBuf[1762] = 256'h2901390147014e0151014f014501330120010e01fc00f400f500f90005011301;
    inBuf[1763] = 256'h1d0125012801200116010e010101f700f100e800df00db00d300cc00c800c400;
    inBuf[1764] = 256'hc400c700cd00d600db00d900d600cc00b800a50093007d006f006a006a007000;
    inBuf[1765] = 256'h7a00850092009b00a000a1009d009400870077006500530045003c0036003600;
    inBuf[1766] = 256'h40004f005d00690070006f006600520037001e000a00fdfffbff040016002c00;
    inBuf[1767] = 256'h3f004d00540051004600360028001c0012000f00120016001a001d001e001c00;
    inBuf[1768] = 256'h140009000300fffffafffaff0000060011001d002200230021001b0013000700;
    inBuf[1769] = 256'hfbfff3ffefffeffff3fff9ff000009000c000700fbffe6ffcaffaeff96ff86ff;
    inBuf[1770] = 256'h82ff89ff9dffb7ffd1ffe6fff2fff0ffe4ffd0ffbaffa7ff97ff91ff97ffa4ff;
    inBuf[1771] = 256'hb4ffc6ffd1ffd3ffcdffbdffa9ff97ff84ff75ff6fff71ff77ff82ff8eff98ff;
    inBuf[1772] = 256'h9effa0ff9fff9bff97ff94ff93ff93ff96ffa0ffaaffb3ffbfffc8ffc9ffc7ff;
    inBuf[1773] = 256'hbeffabff9bff90ff88ff85ff8bff96ffa5ffb5ffc2ffc9ffcaffc4ffb9ffacff;
    inBuf[1774] = 256'ha2ff9eff9dffa3ffb3ffc4ffd2ffe2ffebffe8ffe4ffdaffcbffbdffb0ffa5ff;
    inBuf[1775] = 256'h9eff9aff98ff9aff9cff9dffa1ffa3ffa0ff9dff99ff94ff8eff88ff85ff84ff;
    inBuf[1776] = 256'h84ff89ff92ff9affa1ffa7ffa9ffa7ffa1ff99ff93ff8fff8cff8bff90ff99ff;
    inBuf[1777] = 256'ha1ffa5ffa6ffa2ff9cff95ff8aff7eff77ff78ff7dff84ff8fff9cffa9ffb4ff;
    inBuf[1778] = 256'hb9ffbcffbaffb4ffadffa3ff99ff94ff94ff98ffa1ffb0ffbeffcbffd7ffdaff;
    inBuf[1779] = 256'hd7ffceffbdffa9ff9aff8dff83ff85ff8fff9dffafffc4ffd5ffe1ffe2ffddff;
    inBuf[1780] = 256'hd6ffccffc2ffbbffb9ffbdffc5ffceffd6ffdeffe1ffdeffdbffd6ffcfffc9ff;
    inBuf[1781] = 256'hc5ffc1ffc1ffc3ffc3ffc4ffc6ffc5ffc2ffc0ffbbffb8ffbaffc0ffc9ffd6ff;
    inBuf[1782] = 256'he5fff5ff04000d000d000400f6ffe3ffceffbaffabffa5ffa9ffb4ffc6ffdaff;
    inBuf[1783] = 256'hebfff5fff8fff0ffe0ffccffb5ffa1ff95ff92ff9cffb1ffc9ffe5ff03001900;
    inBuf[1784] = 256'h25002a0021000f00faffe3ffcdffc0ffbaffbaffc2ffd0ffe2fff3ffffff0500;
    inBuf[1785] = 256'h0500fffff5ffe8ffdaffd0ffcaffc8ffceffd8ffe3fff1fffdff020003000100;
    inBuf[1786] = 256'hfbfff1ffe6ffdcffd2ffc5ffbdffb9ffb5ffb2ffb1ffafffacffacffaeffafff;
    inBuf[1787] = 256'hafffaeffadffabffa6ffa0ff9bff97ff93ff90ff8cff8bff8aff85ff80ff7eff;
    inBuf[1788] = 256'h76ff6bff63ff5aff50ff48ff41ff3cff3bff39ff35ff37ff37ff34ff30ff2dff;
    inBuf[1789] = 256'h2cff2bff2bff2dff30ff32ff36ff3aff3bff39ff36ff30ff28ff20ff17ff10ff;
    inBuf[1790] = 256'h0dff0cff0fff15ff19ff1eff22ff1eff1aff17ff0eff04fffefef9fef5fef5fe;
    inBuf[1791] = 256'hf8fefbfefbfefcfefdfefbfef5feeefee8fee1fed9fed4fed2fed0fecafec5fe;
    inBuf[1792] = 256'hc3fec0febbfeb9febbfebbfebbfebefec2fec3fec3fec2fec1febcfeb3feabfe;
    inBuf[1793] = 256'ha8fea3fea0fea2fea6feaefeb8febdfebffec1febcfeb4feadfea4fe9dfe97fe;
    inBuf[1794] = 256'h92fe91fe96fe9bfea2feabfeb4febcfec1febffebefebcfeb6feb0feacfea7fe;
    inBuf[1795] = 256'ha7feaafeabfeb1febafec3fecefed7fedefee4fee8fee5fedffedafed4fecdfe;
    inBuf[1796] = 256'hc7fec5fecbfed7fee4fef2fe03ff13ff1eff21ff1dff17ff10ff05fffafef5fe;
    inBuf[1797] = 256'hf5fefbfe07ff12ff1eff2cff34ff35ff32ff28ff1cff11ff07ff01ff03ff0bff;
    inBuf[1798] = 256'h18ff29ff37ff44ff4eff4fff4cff48ff40ff3cff3aff39ff42ff52ff5eff6cff;
    inBuf[1799] = 256'h78ff7dff7eff78ff6dff61ff55ff4eff4fff55ff5fff70ff83ff93ffa0ffa9ff;
    inBuf[1800] = 256'habffa9ffa2ff9aff96ff95ff9affa3ffafffc1ffd6ffe6ffeffff5fff7fff2ff;
    inBuf[1801] = 256'hebffe2ffdaffd8ffd9ffdaffe0ffecfff6ff01000b00110016001c0021002600;
    inBuf[1802] = 256'h2d00370042004900500056005500510051004e00470049004d00510059006400;
    inBuf[1803] = 256'h6f00780079007500710069005c0053004c004b005500640078009300ad00c000;
    inBuf[1804] = 256'hd100d900d700cd00be00ad009f00950090009400a200b600ca00dd00ef00fb00;
    inBuf[1805] = 256'hfe00fa00f300e700d700cb00c600c800d000e000f4000c012401390147014f01;
    inBuf[1806] = 256'h51014b01420139012e0123011f01210125012f013f015001610171017c018401;
    inBuf[1807] = 256'h850181017d0176016e016d017001740182019401a401b801c801d101d901da01;
    inBuf[1808] = 256'hd101c901c101b801b201af01b001ba01c501d001e001ea01ee01f101ee01e801;
    inBuf[1809] = 256'he501e001db01de01e301e901f60102020b02140218021902180214020f020c02;
    inBuf[1810] = 256'h0a020b02110216021d0227022b022e02320231022c022b022702220224022802;
    inBuf[1811] = 256'h2a023002360238023e0242024102440246024202430244024402470248024702;
    inBuf[1812] = 256'h4b024d024a024f025202510259025d025b02600263025f025f025c0253025302;
    inBuf[1813] = 256'h53024e02520255025702600267026b02740275026f026f026c0261025c025802;
    inBuf[1814] = 256'h53025302530254025c026002620268026a02680266025f0255024d0242023802;
    inBuf[1815] = 256'h33022c0227022a02300236023f02440247024b0247023e02330221020d02ff01;
    inBuf[1816] = 256'hf301e901ea01ef01f9010c021a0223022a02260217020602f101da01c601b601;
    inBuf[1817] = 256'hb001b701c001cf01e401f401fe010302fb01ea01d701be01a301910186018101;
    inBuf[1818] = 256'h89019701a701b801c101c101c201b901a50191017c0168015c01550152015801;
    inBuf[1819] = 256'h5e0164016b016c0166015c014d013b012e012201160112011101120117011801;
    inBuf[1820] = 256'h1801190114010c010401fc00f400ed00e600e200df00d900d300cb00be00b400;
    inBuf[1821] = 256'haa009a008c0083007a0073006f006b0066006000580051004b00420037002f00;
    inBuf[1822] = 256'h290024001f001a0016000f000300f8ffecffdcffcbffbeffb2ffa8ffa4ffa3ff;
    inBuf[1823] = 256'h9eff97ff91ff8bff82ff76ff6bff5fff55ff4eff4fff54ff59ff60ff65ff69ff;
    inBuf[1824] = 256'h69ff63ff57ff48ff37ff27ff1aff0dff04ff01ff01ff04ff05ff04ff00fffafe;
    inBuf[1825] = 256'hf0fee4fed6fecafec0feb8feb4feb3feb3feb7febcfebdfebcfebefebbfeb3fe;
    inBuf[1826] = 256'haafe9efe91fe86fe79fe69fe5dfe52fe46fe3afe32fe2cfe28fe24fe23fe23fe;
    inBuf[1827] = 256'h20fe1cfe15fe0dfe05fefdfdf2fde7fde1fddffddffde3fde8fdecfdf0fdf0fd;
    inBuf[1828] = 256'hecfde6fddafdc9fdbbfdacfd9ffd97fd91fd91fd97fd9dfda3fdacfdb1fdb2fd;
    inBuf[1829] = 256'hb3fdadfda7fda1fd9afd95fd95fd91fd91fd97fd9afd9dfda2fda1fda2fda6fd;
    inBuf[1830] = 256'ha2fd9afd95fd8cfd83fd7dfd72fd6bfd69fd65fd65fd69fd69fd6dfd76fd78fd;
    inBuf[1831] = 256'h79fd79fd73fd6cfd67fd5ffd58fd56fd56fd5bfd64fd6bfd74fd7cfd7dfd7bfd;
    inBuf[1832] = 256'h79fd70fd63fd5afd51fd4dfd4efd4cfd50fd5bfd60fd60fd63fd60fd57fd4ffd;
    inBuf[1833] = 256'h47fd3ffd3cfd3afd3ffd47fd4cfd53fd5afd58fd54fd50fd47fd3dfd34fd2cfd;
    inBuf[1834] = 256'h2bfd2efd2ffd34fd3afd3bfd3cfd3bfd32fd2afd26fd1ffd19fd18fd1bfd22fd;
    inBuf[1835] = 256'h2bfd34fd3ffd48fd4cfd4ffd4ffd4cfd4cfd4cfd49fd4afd4efd4ffd51fd52fd;
    inBuf[1836] = 256'h50fd52fd55fd52fd51fd54fd50fd4ffd53fd51fd4ffd50fd4efd4efd4ffd4efd;
    inBuf[1837] = 256'h53fd5cfd63fd6cfd76fd7afd80fd82fd7afd75fd71fd65fd5dfd5afd57fd5cfd;
    inBuf[1838] = 256'h62fd67fd71fd78fd77fd78fd75fd68fd5ffd59fd52fd51fd56fd5cfd68fd79fd;
    inBuf[1839] = 256'h84fd8dfd93fd92fd8cfd84fd7bfd72fd6dfd6dfd73fd7efd89fd94fd9ffda7fd;
    inBuf[1840] = 256'ha8fda6fda1fd98fd93fd8efd8bfd92fd9cfdaafdbdfdcbfdd2fdd9fdd8fdd0fd;
    inBuf[1841] = 256'hc9fdc0fdb9fdb9fdbafdc0fdd0fdddfdeafdf9fdfffd01fe02fefafdf0fdeafd;
    inBuf[1842] = 256'he3fde2fde9fdf1fd01fe14fe1ffe29fe2ffe2cfe27fe20fe16fe10fe0ffe11fe;
    inBuf[1843] = 256'h1bfe27fe34fe46fe54fe5bfe60fe64fe62fe5efe5cfe5dfe64fe6dfe79fe88fe;
    inBuf[1844] = 256'h95fe9efea5fea8fea3fe9afe92fe8afe87fe8afe8efe97fea5feb0feb8fec2fe;
    inBuf[1845] = 256'hc7fec4febffebafeb5feb3feb3feb8fec7fed7fee7fef7fe03ff07ff06fffdfe;
    inBuf[1846] = 256'heefee2fed6feccfecafeccfed4fee3fef4fe02ff0fff16ff18ff18ff14ff0fff;
    inBuf[1847] = 256'h0bff0aff11ff1dff2cff41ff57ff69ff79ff84ff86ff84ff81ff7aff71ff6cff;
    inBuf[1848] = 256'h6eff72ff78ff83ff90ff9cffa5ffadffb2ffb2ffafffadffabffaeffb7ffc1ff;
    inBuf[1849] = 256'hcdffdbffebfff7fffeff02000200fffff9fff2ffebffe7ffe8ffeaffeffff6ff;
    inBuf[1850] = 256'hfbfffdfffdfff8fff0ffe8ffe0ffdaffdaffe1ffedfffdff0c001e002f003900;
    inBuf[1851] = 256'h400042003c0033002c00250025002b0034004200530063007000780076006f00;
    inBuf[1852] = 256'h640055004a00430043004c005d0073008e00a900bc00c800cc00c900c000b600;
    inBuf[1853] = 256'hac00a500a700b100c100d600eb00ff000f01160114010a01fb00ec00e100d800;
    inBuf[1854] = 256'hd800e300f30005011d01340144014d014d0147013f0136013101330139014801;
    inBuf[1855] = 256'h5f0177019001a401b001b801b601ac01a4019b01920192019a01a601bc01d301;
    inBuf[1856] = 256'he401f501000201020002fa01ee01ec01ef01f401020216022a0243025b026902;
    inBuf[1857] = 256'h76027b02770274026e02650266026b026f027e0290029c02aa02b502b802bc02;
    inBuf[1858] = 256'hbb02b602b702ba02b902c202d102df02f4020803160329033c03460353035d03;
    inBuf[1859] = 256'h62036d037803810391039d03a203ae03bc03c203ca03d403da03e503ee03f403;
    inBuf[1860] = 256'hff0308040a0416042204280437044704530465047704830493049e04a404ac04;
    inBuf[1861] = 256'hb004af04b304b404b504bd04c004c304d004d704d504da04dd04db04de04e004;
    inBuf[1862] = 256'he004eb04f8040305190530053f0556056a0574057f0588058905900598059b05;
    inBuf[1863] = 256'ha805b805c205d505e605ed05f905010601060406050602060b0615061c063006;
    inBuf[1864] = 256'h440655067006830689069806a1069e06a406a606a006a906b406b906c706d306;
    inBuf[1865] = 256'hd606e106e606e006e206dd06d106d206d306d106df06eb06f306080717071a07;
    inBuf[1866] = 256'h240728072007230724071f07280733073a074d075e0766077407790772077107;
    inBuf[1867] = 256'h69075a075a075b07580769077d0789079e07ad07b007b707b207a10799078d07;
    inBuf[1868] = 256'h7b077a077e0781079407a407a907ba07c007b007a40792077507630753074307;
    inBuf[1869] = 256'h4807510754076707770778077c0776076107500739071c070f070607ff060b07;
    inBuf[1870] = 256'h17071e073107380730072e0722070a07ff06f106e006e406ea06ec06fd060807;
    inBuf[1871] = 256'h0a0712070e07fc06f306e006c506bb06b106a606ab06ad06ab06b106a9069506;
    inBuf[1872] = 256'h87067006520641062f061e061f0620061f0629062a06200617060306e305c705;
    inBuf[1873] = 256'ha6058405730567055f0567056d056e056d056005460528050205d704b5049904;
    inBuf[1874] = 256'h860485048c049704ad04be04c104be04ac04890464043a041104f703e703e003;
    inBuf[1875] = 256'heb03fe030c04170416040404e803bf038a0358032a030403f302f002f7020903;
    inBuf[1876] = 256'h1b03250328031b03fa02cd029a0267023b0217020302ff0103020c0217021b02;
    inBuf[1877] = 256'h1302fe01d801a80174013f011001ec00d500ce00d100d900e200e500de00cc00;
    inBuf[1878] = 256'hae0086005c0034001000f4ffe2ffdcffdeffddffddffd9ffccffb5ff96ff6eff;
    inBuf[1879] = 256'h45ff1efff8fedbfec7feb6feabfea1fe90fe7dfe66fe44fe1dfef7fdd1fdadfd;
    inBuf[1880] = 256'h90fd76fd62fd54fd43fd31fd20fd04fde2fcbefc95fc6bfc4afc2bfc11fc00fc;
    inBuf[1881] = 256'hf0fbe3fbd6fbbffba4fb88fb5efb33fb0bfbe1fabffaa9fa94fa87fa86fa7cfa;
    inBuf[1882] = 256'h73fa6cfa53fa33fa15faebf9c2f9a5f986f971f96af95ff95bf95df950f940f9;
    inBuf[1883] = 256'h2ef907f9dbf8b5f883f855f834f811f8f8f7eef7ddf7d0f7c8f7aff795f77df7;
    inBuf[1884] = 256'h52f729f70df7e7f6c7f6b7f69ef68cf687f678f668f65cf63df61ff609f6e1f5;
    inBuf[1885] = 256'hbaf5a0f578f557f545f524f509f5fdf4dff4c4f4bbf4a2f48ff48bf476f467f4;
    inBuf[1886] = 256'h66f451f43df437f41ef407f4fff3e5f3d1f3d0f3bef3b2f3b3f39ff38cf383f3;
    inBuf[1887] = 256'h5ff33bf321f3f2f2cdf2baf29af28cf293f28af28df29ef292f287f285f264f2;
    inBuf[1888] = 256'h46f234f20bf2f0f1edf1dbf1d8f1ecf1eaf1ecf1f6f1dff1c5f1b2f17ff151f1;
    inBuf[1889] = 256'h35f10bf1f4f0f9f0f0f0f9f017f11cf124f135f125f112f106f1ddf0c1f0bdf0;
    inBuf[1890] = 256'ha8f0a5f0bcf0c2f0d5f0f4f0f2f0eff0eef0caf0a8f094f066f047f041f02df0;
    inBuf[1891] = 256'h2ff049f050f061f07af074f06ff06ff04df034f02bf00ef005f015f013f021f0;
    inBuf[1892] = 256'h3ff042f04bf05df04bf038f02ff00ef0f7eff6efe4efe4effbef01f013f033f0;
    inBuf[1893] = 256'h33f036f042f033f02af030f023f025f03bf041f057f07cf085f095f0aef0a6f0;
    inBuf[1894] = 256'ha2f0abf09af096f0a6f0a5f0b4f0d8f0e6f0fbf01bf11ef123f131f122f11cf1;
    inBuf[1895] = 256'h26f11ef128f148f154f16df195f1a4f1b8f1d0f1caf1caf1d1f1c3f1c5f1dbf1;
    inBuf[1896] = 256'he1f1f7f11ff236f256f27df288f293f2a4f29ef29ff2acf2a9f2b3f2d0f2e3f2;
    inBuf[1897] = 256'h03f32ff347f365f389f394f3a0f3b3f3b2f3baf3d1f3dbf3f6f322f43ef464f4;
    inBuf[1898] = 256'h95f4b0f4cff4f4f4fef40df525f529f535f550f55ef579f5a3f5bef5e3f510f6;
    inBuf[1899] = 256'h28f643f664f672f685f69df6a9f6c1f6e3f6f9f61cf74af76cf797f7c6f7e4f7;
    inBuf[1900] = 256'h07f82bf83df855f872f882f89cf8bdf8d6f8fcf826f942f968f994f9b4f9d7f9;
    inBuf[1901] = 256'hfcf916fa38fa5dfa78fa9afac1fae2fa0cfb38fb5cfb85fbaffbd2fbfbfb24fc;
    inBuf[1902] = 256'h45fc6bfc91fcaefccffcf0fc0afd29fd48fd67fd8efdb5fdd8fd04fe32fe5afe;
    inBuf[1903] = 256'h85feaefed2fef6fe13ff2dff4dff6aff88ffb0ffdaff06003a0067009200c200;
    inBuf[1904] = 256'he700060125013d01550171018b01ac01d801030236026e02a202d7020a033003;
    inBuf[1905] = 256'h540374038a03a503c103da0300042d0456048d04c904fb04310563058705ad05;
    inBuf[1906] = 256'hcc05db05f4050f06240649067806a506e206210755078f07c007dd07fd071508;
    inBuf[1907] = 256'h1a082b0840084e0871089f08cb080a0948097709af09d909e909020a120a100a;
    inBuf[1908] = 256'h220a3d0a560a890ac10af10a350b750b9d0bcb0be60be80bf50bfa0bf30b0c0c;
    inBuf[1909] = 256'h2a0c440c7f0cbc0cec0c2d0d5d0d720d920da30d9c0dab0db70dbd0de60d130e;
    inBuf[1910] = 256'h3a0e800ec00eea0e1e0f410f480f580f590f4b0f5a0f690f720f9e0fce0ff30f;
    inBuf[1911] = 256'h2f105f107a10a310b610ae10bb10c010b610cd10e510f7102d1160118311be11;
    inBuf[1912] = 256'he811f31110121b120a1212121212031218122e123c126c129612ac12db12fa12;
    inBuf[1913] = 256'hfb120c130b13f412fb12fa12ee120c1328133c1373139e13b113d813ea13df13;
    inBuf[1914] = 256'he613d813b713b513ae13a113bf13db13eb131b143c1440145714551438142f14;
    inBuf[1915] = 256'h1714f413f913fc13f9131f14411452147b148f1485148c147a144b143b142414;
    inBuf[1916] = 256'h02140a141414141437144e144e1464146214421437141b14ee13e513d713c013;
    inBuf[1917] = 256'hd213de13dd13fa130414f413f913e813c013b4139a137513781371135f137013;
    inBuf[1918] = 256'h7313611369135e133c1334131b13f212e812d412b412b612ab12931299128f12;
    inBuf[1919] = 256'h6e12671252122c1222120d12ec11e911d911bb11ba11a81184117b1165113d11;
    inBuf[1920] = 256'h32111c11f810f010dd10ba10b3109f1079106c1052102a101d100310e00fdd0f;
    inBuf[1921] = 256'hcc0fad0faa0f970f720f650f470f1d0f0d0fef0eca0ec30eb00e930e920e830e;
    inBuf[1922] = 256'h620e540e330e010ee40dba0d850d6d0d500d320d310d290d170d180d060de10c;
    inBuf[1923] = 256'hc70c9a0c600c380c080cd80bc80bb70ba60bb00baf0ba10b9b0b7c0b480b1a0b;
    inBuf[1924] = 256'hd50a870a540a230af609ec09e809e609f809f809e409d309a80964092609dd08;
    inBuf[1925] = 256'h920862083c0823082b0835083b084b0843082208f807b4075d071007c0067b06;
    inBuf[1926] = 256'h56063b0630063e064b06500653063c060d06d40587053105e804a40472045d04;
    inBuf[1927] = 256'h5504580467046f04680456042b04ee03a90356030303c1028902620255025302;
    inBuf[1928] = 256'h570261026202520236020502c3017b012f01e800b00085006900610063006900;
    inBuf[1929] = 256'h6d00660050002d00f6ffb0ff63ff16ffd4fe9efe76fe65fe64fe68fe70fe74fe;
    inBuf[1930] = 256'h68fe4cfe1cfedafd90fd40fdf0fcb0fc80fc63fc5dfc62fc6dfc7afc77fc63fc;
    inBuf[1931] = 256'h3efc01fcb4fb65fb14fbcffaa0fa7efa73fa7efa87fa91fa99fa88fa62fa2efa;
    inBuf[1932] = 256'he2f98ff943f9f9f8c2f8a5f894f896f8a7f8adf8adf8a8f883f84ff818f8cff7;
    inBuf[1933] = 256'h88f751f71df7fcf6f4f6ecf6eef6faf6f0f6dcf6c4f691f654f61ef6daf59df5;
    inBuf[1934] = 256'h79f553f53af536f527f51bf516f5f9f4d9f4bff48bf459f437f405f4def3cdf3;
    inBuf[1935] = 256'haff39af394f377f35df34cf31ef3f1f2d3f29ef273f25af22ff20ff204f2e1f1;
    inBuf[1936] = 256'hc4f1b6f18ff16bf156f128f1fff0eaf0c1f0a6f0a1f086f073f071f053f036f0;
    inBuf[1937] = 256'h21f0eeefc1efa4ef6def41ef2fef0beff5eef7eee1eed4eed6eeb5ee95ee80ee;
    inBuf[1938] = 256'h49ee17eefaedc6eda7eda8ed95ed91eda8eda0ed9ceda2ed7eed5aed40ed02ed;
    inBuf[1939] = 256'hcfecb6ec88ec72ec7eec74ec7bec9aec92ec8aec8dec63ec3aec22eceaebc3eb;
    inBuf[1940] = 256'hbbeb9feb9cebb6ebb3ebbcebd6ebc9ebbbebb7eb8ceb69eb5aeb31eb1eeb27eb;
    inBuf[1941] = 256'h19eb1deb39eb34eb37eb47eb2feb1eeb1feb00ebf2eafdeaeaeae9ea00ebf4ea;
    inBuf[1942] = 256'hf0ea00ebebeaddeae3eac7eabceacdeac4eaceeaf2eaf5ea02eb1eeb0feb05eb;
    inBuf[1943] = 256'h0aebe9ead6eae0ead4eae1ea0aeb17eb38eb69eb6feb77eb86eb64eb47eb3beb;
    inBuf[1944] = 256'h10ebfdea0feb12eb33eb75eb9debd2eb0eec19ec22ec2eec0aeceeebe7ebc9eb;
    inBuf[1945] = 256'hc6ebe9ebffeb30ec7beca4ecd2ec02ed00edf7ecefecbeec9aec94ec7eec87ec;
    inBuf[1946] = 256'hb7ecd9ec12ed64ed93edc0edf0edf3edf1edf5edd7edcbedd8edd3edeaed20ee;
    inBuf[1947] = 256'h41ee73eeb2eecbeee4eeffeef3eeefeef5eedeeedbeef1eef5ee10ef41ef5aef;
    inBuf[1948] = 256'h84efbdefd6eff8ef25f033f04bf070f07bf093f0b8f0c2f0d6f0f6f0fdf011f1;
    inBuf[1949] = 256'h31f13af154f182f19bf1bef1eaf1fdf118f237f23cf249f261f265f27cf2a8f2;
    inBuf[1950] = 256'hcaf201f34af380f3bff302f424f442f45df457f457f462f461f474f49df4bff4;
    inBuf[1951] = 256'hf7f43df570f5aaf5e3f5fcf513f62af62bf637f64ff661f68cf6caf602f74af7;
    inBuf[1952] = 256'h98f7cff704f834f849f85cf86ff876f88af8a6f8c2f8f1f829f958f990f9c7f9;
    inBuf[1953] = 256'hedf913fa33fa47fa62fa81faa0fad3fa0dfb43fb86fbc4fbf2fb1ffc42fc53fc;
    inBuf[1954] = 256'h64fc74fc85fca6fcd1fc02fd44fd8dfdcffd10fe41fe5efe6ffe71fe69fe69fe;
    inBuf[1955] = 256'h75fe91fec8fe14ff6fffd7ff37008900c700e300e300d200ae00880077007d00;
    inBuf[1956] = 256'ha600f4005c01d8015702c0020f033b0338031503e102a4027c0277029602e802;
    inBuf[1957] = 256'h6503f4038f041c057e05b705b90583053605dc04850459045f0494040805a405;
    inBuf[1958] = 256'h4706ea066c07b707d307b40761070707af0668065f068f06ed0685073308d708;
    inBuf[1959] = 256'h6f09d109ed09d9098f091a09ae0855081c0829087008e0088409310ac40a410b;
    inBuf[1960] = 256'h8b0b8f0b6c0b210bbb0a6b0a370a250a5a0abe0a3b0bda0b700cdb0c2d0d470d;
    inBuf[1961] = 256'h230de90c920c2c0cef0bd10bd20b180c810cf50c840dff0d4e0e8a0e950e6c0e;
    inBuf[1962] = 256'h420e080ec90db90dc30de00d340e960eef0e570fa10fc20fd90fc80f920f6d0f;
    inBuf[1963] = 256'h460f200f2a0f480f6f0fc00f11104d109510c010c610d110c710a810a410a110;
    inBuf[1964] = 256'h9b10bf10e81006113f116a117811921196117e117a116f115b116d1181118e11;
    inBuf[1965] = 256'hbf11e411f2111712281219121d121412f91100120412ff11231240124c127312;
    inBuf[1966] = 256'h89127f12831274124d1240122c121212221234123f1270129712a912d012df12;
    inBuf[1967] = 256'hcf12cd12b512871278126112431250125c1260128912a512a912c012bf129f12;
    inBuf[1968] = 256'h9512771247123a122b1218122f12471258128d12b312bf12de12e312c312b412;
    inBuf[1969] = 256'h92125a12421224120012081210120f1231124512421257125412321225120812;
    inBuf[1970] = 256'hd811cc11be11ac11c611e011f11120123f1246125c1254122d121612ea11aa11;
    inBuf[1971] = 256'h8b1167113e113e1140113f115e1170116c117c11751150113f111d11ec10de10;
    inBuf[1972] = 256'hcd10b910cd10e410f2101a1136113a11461134110211dc10a11055102910fd0f;
    inBuf[1973] = 256'hd00fcf0fd30fd40ff40f0710061011100110d60fbb0f8b0f4c0f2f0f150fff0e;
    inBuf[1974] = 256'h130f290f390f630f790f730f730f520f0e0fd40e880e320efd0dcc0da40dab0d;
    inBuf[1975] = 256'hb70dc10de70dfe0dfa0df70dd60d970d600d1b0dcf0ca50c860c710c870ca20c;
    inBuf[1976] = 256'hb80cdd0cee0cde0cc60c8d0c330cdd0b7e0b1f0be50abd0aa70abc0ada0af50a;
    inBuf[1977] = 256'h1a0b230b0c0be90aa40a460af1099809480921090f0912093a0960097c099909;
    inBuf[1978] = 256'h930964092409c6085708f6079b0754073b073707470772079607a907b3079907;
    inBuf[1979] = 256'h5e071407b3064c06fa05b6058b0585059005a905d005e605e605d605a7056005;
    inBuf[1980] = 256'h1105b90463042404f603dd03df03eb03fc030e041104ff03e003aa0363031b03;
    inBuf[1981] = 256'hd202910261023e02290221021e021b0217020502e901c30192015b012501f100;
    inBuf[1982] = 256'hc2009b007e006b005c004c003d0028000a00e8ffbdff8cff5aff23ffedfebffe;
    inBuf[1983] = 256'h91fe65fe45fe25fe07fef0fdd3fdb3fd96fd72fd4afd27fdfefcd5fcb4fc90fc;
    inBuf[1984] = 256'h6bfc4cfc2afc07fce9fbc1fb98fb72fb42fb11fbe6fab3fa83fa5cfa30fa08fa;
    inBuf[1985] = 256'he7f9bef995f976f94df924f903f9dbf8b7f89df87bf85cf846f825f804f8ecf7;
    inBuf[1986] = 256'hc6f79af773f73ff70cf7e3f6aef67ff65ef635f614f602f6e2f5c3f5aff58cf5;
    inBuf[1987] = 256'h67f54bf51cf5f0f4d1f4a4f47ef46cf450f43cf43af428f418f412f4f1f3ccf3;
    inBuf[1988] = 256'haef374f33bf311f3d7f2a7f290f271f263f26cf265f265f270f25bf241f22cf2;
    inBuf[1989] = 256'hf4f1bbf195f15df134f129f118f118f131f136f140f151f13cf11df101f1c2f0;
    inBuf[1990] = 256'h80f051f016f0f0efecefe4eff2ef1cf030f047f062f054f03df027f0edefb5ef;
    inBuf[1991] = 256'h8fef58ef39ef3def38ef4aef75ef85ef9aefb4efa1ef88ef73ef38ef06efebee;
    inBuf[1992] = 256'hbeeeaaeebaeebeeedaee0def23ef3fef5fef51ef40ef31effbeecceeb3ee88ee;
    inBuf[1993] = 256'h75ee80ee7dee92eebbeec7eedaeef4eee4eed4eecdeea3ee85ee7cee61ee5eee;
    inBuf[1994] = 256'h76ee7cee95eec1eecfeee1eef8eee8eeddeedceebbeea6eea4ee8dee87ee98ee;
    inBuf[1995] = 256'h93ee9ceeb5eeb3eebaeed0eec8eecbeedeeed6eedceef5eef6ee00ef18ef15ef;
    inBuf[1996] = 256'h1aef2def27ef2def44ef46ef56ef76ef7fef91efabefa8efabefb6efa4ef9bef;
    inBuf[1997] = 256'ha1ef95ef9defbcefcfeff5ef2bf04bf073f0a0f0a8f0b1f0bdf0acf0a3f0abf0;
    inBuf[1998] = 256'ha1f0adf0d2f0ebf015f152f176f19ff1cbf1d1f1d4f1d9f1bff1b0f1b4f1a7f1;
    inBuf[1999] = 256'hb2f1dcf1fdf132f27af2acf2e1f218f32af338f344f32ef31ef31ff311f31af3;
    inBuf[2000] = 256'h41f362f398f3e2f317f44ef484f495f49ef4a4f489f473f46cf45af462f487f4;
    inBuf[2001] = 256'haaf4e4f431f56cf5abf5e6f5fcf509f610f6f9f5eaf5e6f5daf5e5f50cf632f6;
    inBuf[2002] = 256'h6df6b6f6f0f62bf761f775f782f786f771f762f75cf751f75df77ff7a3f7dbf7;
    inBuf[2003] = 256'h1ef854f88ff8c4f8dcf8f2f801f9f8f8f5f8f8f8f5f807f92bf94bf97ff9bdf9;
    inBuf[2004] = 256'hedf923fa53fa6afa7dfa8afa84fa83fa88fa85fa94fab1facefafbfa30fb5bfb;
    inBuf[2005] = 256'h8bfbb6fbd1fbebfbfefb04fc11fc22fc31fc4cfc6ffc90fcb9fce4fc08fd2cfd;
    inBuf[2006] = 256'h4afd5efd74fd86fd95fda8fdbffdd7fdf7fd17fe35fe56fe72fe89fea2feb8fe;
    inBuf[2007] = 256'hccfee7fe05ff28ff50ff78ffa0ffcaffecff07001f002f003a00470055006800;
    inBuf[2008] = 256'h8600aa00d6000801370165019001ab01bd01c901cd01d101d801e201f9011e02;
    inBuf[2009] = 256'h48027c02b802ee022003490362037103760370036d036f0373038703ab03d603;
    inBuf[2010] = 256'h0c0447047e04b104d904ef04fd04fc04f004e704e104de04ee040c0533056905;
    inBuf[2011] = 256'ha205d7050b06300642064d064a063b06310626062206330650067406a906e206;
    inBuf[2012] = 256'h13074407660774077c0775075f07530749073f074d0765078007af07e1070708;
    inBuf[2013] = 256'h310850085b08660865085608520850084c085d0878089208bc08e70806092c09;
    inBuf[2014] = 256'h480951095c0960095409530952094b095809690976099609b709cc09ec09060a;
    inBuf[2015] = 256'h100a230a300a2f0a3b0a460a490a5c0a6f0a7a0a960aaf0abc0ad50ae90aef0a;
    inBuf[2016] = 256'h010b0e0b0f0b1e0b2c0b2f0b410b4f0b500b610b6d0b6e0b7f0b8e0b940bb00b;
    inBuf[2017] = 256'hca0bda0bfc0b190c250c3f0c4c0c470c4f0c4d0c3d0c440c4c0c4e0c6b0c890c;
    inBuf[2018] = 256'h9d0cc60ce60cef0c030d070df40cf10ce70cd00cd90ce70cf00c190d450d650d;
    inBuf[2019] = 256'h980dbb0dc30dd40dd30db70dac0d9b0d810d870d920d9a0dc20dea0d030e2d0e;
    inBuf[2020] = 256'h4a0e4e0e5c0e590e410e3d0e330e200e2b0e390e400e640e850e960ebb0ed20e;
    inBuf[2021] = 256'hd20ee00ee10ecf0ed00ec60eb10eb80ebb0eb40ec90edb0ee00efd0e110f150f;
    inBuf[2022] = 256'h2d0f370f2e0f3a0f390f270f2c0f270f160f1f0f220f1c0f310f3d0f3d0f550f;
    inBuf[2023] = 256'h600f570f630f5f0f480f460f3a0f1f0f200f1a0f0d0f200f2d0f2f0f4d0f620f;
    inBuf[2024] = 256'h640f780f7b0f690f670f550f320f270f150ffa0eff0e010ffc0e170f2b0f300f;
    inBuf[2025] = 256'h480f500f410f400f2c0f050ff30edb0ebb0ebc0ebe0ebf0edf0efa0e070f260f;
    inBuf[2026] = 256'h320f250f200f050fd50eb70e910e680e600e5b0e590e780e930ea40ec50ed20e;
    inBuf[2027] = 256'hc70ec20ea60e780e5b0e350e0c0e040eff0dfc0d190e300e3b0e560e5b0e490e;
    inBuf[2028] = 256'h3c0e190ee40dc10d950d660d570d4c0d410d550d650d6a0d7e0d820d710d680d;
    inBuf[2029] = 256'h4c0d1d0d000dda0cac0c9b0c890c730c780c790c6f0c750c6f0c580c4e0c340c;
    inBuf[2030] = 256'h0b0cf20bd10ba50b900b790b5c0b540b480b350b350b2d0b180b110bff0ae00a;
    inBuf[2031] = 256'hce0aaf0a820a640a3f0a110af609d609b409a709970983098109760961095709;
    inBuf[2032] = 256'h40091c09ff08d508a4088108590831081e080808f307ef07e107ce07c207a407;
    inBuf[2033] = 256'h7a0757072407eb06bd0689065a063e0621060a060506fb05ee05ea05d705b905;
    inBuf[2034] = 256'h9e0573053f051105d804a10478044c04290416040104ef03e703d403bb03a103;
    inBuf[2035] = 256'h760341030b03ca028c0257022402fe01eb01dd01db01e001de01d801c801a301;
    inBuf[2036] = 256'h71013101e100930049000200ceffabff95ff90ff91ff8eff8cff7aff53ff22ff;
    inBuf[2037] = 256'hdffe8efe41fef5fdb1fd86fd68fd59fd60fd67fd6bfd70fd5efd37fd06fdbcfc;
    inBuf[2038] = 256'h65fc12fcbafb6cfb38fb0dfbf5faf6faf5faf6fafcfaecfacbfaa2fa5ffa10fa;
    inBuf[2039] = 256'hc7f975f92bf9fbf8d1f8b9f8baf8b7f8b9f8c0f8aef88df866f820f8cff782f7;
    inBuf[2040] = 256'h28f7daf6a5f673f656f654f64ef651f65cf64cf634f618f6ddf59bf55ef511f5;
    inBuf[2041] = 256'hd0f4a7f479f460f45ef450f449f44cf431f411f4f1f3b3f376f343f3fef2c8f2;
    inBuf[2042] = 256'haaf280f268f267f253f248f247f22af20ff2fbf1ccf1a1f183f150f129f114f1;
    inBuf[2043] = 256'heaf0c9f0bbf095f076f067f03ff01ff010f0e9efccefc2ef9eef81ef75ef4def;
    inBuf[2044] = 256'h29ef15efe7eec2eeb2ee8cee74ee73ee5dee51ee58ee41ee2cee23eef7edcded;
    inBuf[2045] = 256'hb2ed7bed50ed3eed19ed09ed15ed0ded10ed27ed1eed16ed17edf1ecccecb7ec;
    inBuf[2046] = 256'h83ec5eec53ec34ec2cec41ec3eec48ec65ec5cec55ec57ec2fec0becf7ebc2eb;
    inBuf[2047] = 256'h9deb96eb79eb72eb8aeb86eb93ebb3ebacebaaebb4eb91eb74eb68eb38eb15eb;
    inBuf[2048] = 256'h0eebeeeae3eaf4eae7eaeaea07ebfeeaffea12ebfceaedeaf1eaceeab7eab7ea;
    inBuf[2049] = 256'h95ea87ea94ea84ea88eaa8eaa8eab6ead8ead4ead7eae6eacbeab8eab6ea8fea;
    inBuf[2050] = 256'h7aea80ea6eea74ea9aeaa7eac7eafbea0beb20eb3deb2deb20eb1febfaeae6ea;
    inBuf[2051] = 256'hedeadfeaecea1beb33eb60eb9febb7ebd4ebf5ebe7ebdbebdaebb5eba3ebaceb;
    inBuf[2052] = 256'ha2ebb8ebedeb0cec41ec88eca8ecccecf3ececece8ecedeccfecc2eccfecc9ec;
    inBuf[2053] = 256'hdfec12ed2fed60eda0edbceddcedffedf8edf4edf9ede0edd9edeaedeaed06ee;
    inBuf[2054] = 256'h3dee61ee96eed9eefcee21ef48ef49ef4def59ef49ef48ef5eef65ef83efb9ef;
    inBuf[2055] = 256'hddef11f052f076f09df0c9f0d6f0eaf008f110f127f153f172f1a3f1e4f113f2;
    inBuf[2056] = 256'h4df28ef2b4f2e0f210f327f347f371f38bf3b3f3e7f30ef442f47ef4a8f4daf4;
    inBuf[2057] = 256'h11f533f55ef58ff5b2f5dff516f640f674f6aff6dbf60bf73ef75ef784f7aff7;
    inBuf[2058] = 256'hcaf7eff71cf841f870f8a5f8cef8fdf82df94bf96df98ff9a3f9bdf9dff9fbf9;
    inBuf[2059] = 256'h24fa58fa86fabffafcfa2dfb5ffb8dfbaafbc7fbe2fbf4fb0dfc2bfc4afc76fc;
    inBuf[2060] = 256'haafcddfc17fd50fd7ffdadfdd5fdf0fd0bfe25fe3dfe5ffe89feb6fef1fe31ff;
    inBuf[2061] = 256'h71ffb4fff0ff2300510073008e00a900c100dd0003012f016401a001dd011a02;
    inBuf[2062] = 256'h54028302ac02d002e80200031d03390360039003c203fc0339046c049d04c704;
    inBuf[2063] = 256'he104f8040c0519052d05490567059405c705f4052806560674069006a306a706;
    inBuf[2064] = 256'hb006bd06c606e206080730076807a107cf070008280839084c08580857086608;
    inBuf[2065] = 256'h7b088e08ba08ef0820096209a109ce09010a2a0a3c0a580a700a7d0aa10acb0a;
    inBuf[2066] = 256'hf00a2f0b720bab0bf60b390c670ca10cd00cea0c130d380d4f0d7e0dad0dd10d;
    inBuf[2067] = 256'h0f0e4c0e790ebb0ef70e1e0f580f8a0fa40fd20ff80f0b103210521060108610;
    inBuf[2068] = 256'ha710b510dc10fd100c1132114f115711741187118211921199118a1194119911;
    inBuf[2069] = 256'h8d119e11ab11a811c011d111cd11e011e711d411d811cf11b211b011a8119011;
    inBuf[2070] = 256'h9911a2119b11b511c811c511dc11e811da11e211dd11c311c911ca11bc11d511;
    inBuf[2071] = 256'hed11f711241249125912811298129312a612a81293129f12a6129f12c212e412;
    inBuf[2072] = 256'hf7122e135a136d139a13b213ab13bd13be13a813b613bf13bc13e21304141514;
    inBuf[2073] = 256'h48146a146e148b1490147414731461143b143a14341423143c144d144d146c14;
    inBuf[2074] = 256'h79146a147214621438142b141214e813e713e213d213eb13fa13f5130c140f14;
    inBuf[2075] = 256'hf613f813e513bb13b413a5138c13a013b013b413de13fd13041424142d141b14;
    inBuf[2076] = 256'h24141e14061417142914331469149d14c2140615361548156e15781565157015;
    inBuf[2077] = 256'h6d155e157e15a115bd15051645166f16b016d416d016db16c9169b168b167516;
    inBuf[2078] = 256'h561668167e168a16bc16df16e316f416e216a71678163016d115951557151615;
    inBuf[2079] = 256'h0415f414da14df14cf14a0147d143914d31380131a13a61257120812ba119711;
    inBuf[2080] = 256'h711140112c110511c51096104e10f00fac0f5b0f010fcd0e980e610e500e390e;
    inBuf[2081] = 256'h180e150e020edf0dd20db40d850d6f0d4c0d200d130dfe0ce30ce90ce90ce10c;
    inBuf[2082] = 256'hf60c010d010d160d1b0d120d1b0d130dfd0cfb0cef0cdb0ce20ce30ce00cf70c;
    inBuf[2083] = 256'h050d0a0d220d270d1b0d1b0d080de30cca0ca40c780c610c420c220c1a0c050c;
    inBuf[2084] = 256'hea0be00bc70b9f0b820b500b110be10aa30a600a310af809bf099e0973094409;
    inBuf[2085] = 256'h2709fe08ce08a908750838080708ca07880757071c07e206be0695066c065806;
    inBuf[2086] = 256'h410629061d060706ee05de05c205a0058a056b054c053c052b05200525052805;
    inBuf[2087] = 256'h30053f0548054d0553054b053d0530051705fe04eb04d604c704c004ba04bc04;
    inBuf[2088] = 256'hc004bb04b604ad049804790450041b04e403aa036b033203fb02c50297026702;
    inBuf[2089] = 256'h33020202c7017c012f01d5006c00040094ff1fffb4fe4cfee7fd91fd3dfde8fc;
    inBuf[2090] = 256'h9ffc4efcf5fb9efb3cfbcefa64faf3f982f91cf9b6f858f80ff8c8f789f75bf7;
    inBuf[2091] = 256'h29f7f4f6c8f691f654f61df6d9f597f565f52ef502f5eef4dbf4d6f4e6f4f0f4;
    inBuf[2092] = 256'hfbf411f517f518f51cf50cf5fcf4f7f4e6f4e1f4f1f4fbf413f53ff55ff583f5;
    inBuf[2093] = 256'haff5c2f5cef5dbf5cef5bef5b5f59af589f58af57df57cf58cf588f588f591f5;
    inBuf[2094] = 256'h7df564f551f520f5ecf4c4f485f44bf423f4e8f3b2f38ff357f323f300f3c7f2;
    inBuf[2095] = 256'h8ef262f21ff2def1abf160f116f1dbf089f03df006f0bdef7def58ef24effcee;
    inBuf[2096] = 256'hebeec6eea7ee97ee6cee41ee23eeededbceda3ed7ced69ed73ed71ed82edabed;
    inBuf[2097] = 256'hbdedd3edf3edefedeaedeeedd1edbeedc1edb1edbbede4edfced29ee6bee8dee;
    inBuf[2098] = 256'hb3eee1eee1eedeeee4eec2eea8eea6ee88ee80ee98ee94eea0eec2eebaeeb2ee;
    inBuf[2099] = 256'hb2ee7fee46ee18eebded68ed2cedd2ec8dec69ec27ecf7ebe1eba4eb6beb40eb;
    inBuf[2100] = 256'he4ea86ea38eac0e953e901e994e83de80be8bde785e76ae72ce7f9e6d8e689e6;
    inBuf[2101] = 256'h41e60de6b5e56ce541e5fee4d6e4d2e4b7e4b6e4d4e4d3e4e2e407e507e515e5;
    inBuf[2102] = 256'h37e538e54be578e589e5b1e5f4e51ae656e6a9e6dbe61fe779e7ade7f2e74de8;
    inBuf[2103] = 256'h81e8c6e81de94ce989e9d9e901ea38ea83eaaaeae5ea37eb66eba6ebf7eb1dec;
    inBuf[2104] = 256'h50ec8eec97eca2ecb8eca0ec94ec9bec7fec79ec90ec87ec90ecafeca7eca3ec;
    inBuf[2105] = 256'ha7ec7aec4dec27ecd7eb94eb69eb23ebf6eae9eac7eabaeac6eab2eaa4ea9cea;
    inBuf[2106] = 256'h69ea39ea12eacbe993e973e942e92ee93de93fe95ae98ee9a7e9cce9fae901ea;
    inBuf[2107] = 256'h0bea20ea18ea20ea3fea4dea79eac6ea04eb5bebc8eb1aec77ecdbec18ed5bed;
    inBuf[2108] = 256'ha7edcfed06ee53ee8aeed9ee44ef98ef03f07ef0d8f03af19ff1d9f117f25bf2;
    inBuf[2109] = 256'h79f2a0f2d7f2f2f220f35ef382f3b5f3f2f310f435f45ff467f477f48af482f4;
    inBuf[2110] = 256'h88f495f487f489f495f48af489f490f47ff478f479f468f463f463f451f44df4;
    inBuf[2111] = 256'h4ef43bf433f430f41df416f41af418f426f444f461f48ef4c8f4fbf436f573f5;
    inBuf[2112] = 256'ha0f5d0f502f629f659f692f6ccf61bf778f7d7f748f8bff82bf99af903fa57fa;
    inBuf[2113] = 256'ha9faf8fa37fb80fbd5fb2bfc94fc09fd7efd01fe85fef8fe66ffc5ff0a004a00;
    inBuf[2114] = 256'h8100a600d100030133017001b401f40139027702a102c202d202cd02c102aa02;
    inBuf[2115] = 256'h8c02770265025502540257025a025f025a024a0231020a02d901a5016b013201;
    inBuf[2116] = 256'h0101d500b000940079006500510036001d000100dfffc3ffa8ff8dff80ff79ff;
    inBuf[2117] = 256'h73ff7aff87ff94ffaaffc0ffd3ffefff0f002b0054008400b200ed002b016201;
    inBuf[2118] = 256'ha401e90128027302c00208035e03bb0312047704e2044005a30507065a06b106;
    inBuf[2119] = 256'h06074f07a307f80742089c08ff085509b309130a5f0aae0af70a290b600b960b;
    inBuf[2120] = 256'hbc0beb0b1b0c410c790cb20cdd0c130d430d5e0d820d9d0da10db10dbb0db50d;
    inBuf[2121] = 256'hc30dcf0dcd0de40dfa0d010e1d0e330e380e530e640e640e7e0e900e950eba0e;
    inBuf[2122] = 256'hd90eea0e1e0f4d0f690fa30fd40ff10f2a1058107110a810d710f61039117411;
    inBuf[2123] = 256'h9d11ec1134126a12be12051335138013bf13ea1332146e149814e31421154915;
    inBuf[2124] = 256'h8f15c615e1150f16281625163516341622162a16241612161e161b1604160116;
    inBuf[2125] = 256'he815b21587154415eb14a5144e14f013af1365131613e2129d124a1201129b11;
    inBuf[2126] = 256'h1f11ac101d10850f040f770eef0d8b0d200db70c6b0c100cab0b560be30a640a;
    inBuf[2127] = 256'hfc097e090109a8084b08f707ce079f076f075f073d070d07f306c50688066906;
    inBuf[2128] = 256'h4206180618061906190642066a068806c206f306150750078207a707e9072908;
    inBuf[2129] = 256'h5e08b5080c095209b1090c0a530ab20a0e0b570bb60b150c660ccf0c380d8c0d;
    inBuf[2130] = 256'hf40d550e9a0eee0e3e0f760fbf0f0a1048109c10ef1035118f11df1112125412;
    inBuf[2131] = 256'h86129712b612cd12cf12ee121113291362139a13c413081439144a146e147a14;
    inBuf[2132] = 256'h65146a1467145314681480148f14cc14051528156a1596159f15bf15c515a915;
    inBuf[2133] = 256'hb015ae159d15be15e015f91545168a16bb160d1745175a178a179d179217a717;
    inBuf[2134] = 256'had17a317c517de17eb171e1841184e1875187f186a18681848180f18ed17ba17;
    inBuf[2135] = 256'h7b1758172c17f916e016b81683165e161e16ca157c1513159b142d14a2130d13;
    inBuf[2136] = 256'h8b12f9116611e4105210c10f3e0fa40e060e730dc50c0f0c640ba40ae5093309;
    inBuf[2137] = 256'h7208b90715076506c0052d058b04f1036703cb023102a40105016800dbff44ff;
    inBuf[2138] = 256'hb7fe3cfebafd46fdedfc91fc3ffc04fcc6fb8ffb69fb3bfb0dfbeefacbfaabfa;
    inBuf[2139] = 256'h9bfa8ffa8bfaa0fac0faeafa29fb71fbb8fb06fc4ffc8bfccafc06fd35fd6bfd;
    inBuf[2140] = 256'hacfdeffd4bfec0fe39ffc5ff6300f2007e010a027c02df023c038503d0032804;
    inBuf[2141] = 256'h7d04e5046605e805730606078607fd076708af08ed08240947097209a809e109;
    inBuf[2142] = 256'h310a8f0aec0a560bba0b040c4c0c810c970cab0cb40cb00cc10cd60ceb0c1c0d;
    inBuf[2143] = 256'h520d810dc30dfb0d1d0e470e5d0e5c0e6b0e700e650e720e7e0e840ea30ec00e;
    inBuf[2144] = 256'hd20ef80e130f1f0f390f470f440f4f0f4c0f3c0f370f240f080ffd0ee70ecb0e;
    inBuf[2145] = 256'hc00ead0e960e8f0e7d0e640e4e0e250ef20dbb0d6f0d1f0dce0c6c0c140cc40b;
    inBuf[2146] = 256'h670b150bc90a6c0a110aad092d09ac081c086e07c6061c066105b90417046e03;
    inBuf[2147] = 256'hdf025302b80129019200e0ff30ff71fe9afdccfcf6fb18fb50fa86f9bdf80ff8;
    inBuf[2148] = 256'h60f7abf60cf662f5aaf4fff346f381f2cdf115f15ef0bfef22ef90ee1aeea8ed;
    inBuf[2149] = 256'h3aeddfec81ec25ecd6eb7ceb29ebe5ea99ea5aea31ea09eaf3e9f1e9eee9fae9;
    inBuf[2150] = 256'h17ea2dea4fea7bea9fead3ea11eb46eb91ebeeeb45ecb0ec29ed98ed19eea4ee;
    inBuf[2151] = 256'h1defa6ef36f0b7f047f1daf15bf2eef288f30ff4a3f43af5bbf546f6d3f64af7;
    inBuf[2152] = 256'hcef755f8c8f848f9cbf93cfab9fa35fb99fb05fc6afcb1fcfefc48fd7afdb3fd;
    inBuf[2153] = 256'heefd1dfe57fe93febffef3fe23ff3fff5bff71ff72ff73ff72ff69ff6aff72ff;
    inBuf[2154] = 256'h77ff86ff98ffa3ffb1ffbaffafff9cff85ff63ff43ff27ff0cff00ff03ff08ff;
    inBuf[2155] = 256'h1aff32ff3dff41ff41ff2eff0effedfec0fe92fe72fe57fe48fe4efe50fe53fe;
    inBuf[2156] = 256'h5cfe53fe39fe1afedffd98fd57fd04fdb6fc80fc3ffc05fce7fbb6fb78fb47fb;
    inBuf[2157] = 256'hf9fa96fa38fabbf934f9c2f839f8b1f749f7d0f654f6f2f572f5e4f467f4c2f3;
    inBuf[2158] = 256'h10f373f2b5f1f1f04cf08fefd5ee3fee8fede1ec51ec9eebe6ea4cea95e9dde8;
    inBuf[2159] = 256'h47e898e7f0e669e6cce538e5c2e431e4a8e33ae3b0e22fe2cbe152e1ebe0a6e0;
    inBuf[2160] = 256'h52e014e0f5dfc4dfa8dfa7df8edf87df9adf97dfa9dfd6dff4df2ce081e0c9e0;
    inBuf[2161] = 256'h2fe1ace112e294e22be3a3e32ce4c6e448e5dee584e613e7c1e783e82ee9f5e9;
    inBuf[2162] = 256'hccea82eb48ec15edb9ed6aee1fefaaef48f0f5f07ff121f2d6f269f30ff4bcf4;
    inBuf[2163] = 256'h39f5bff541f68af6d5f623f743f770f7abf7c2f7eef72bf843f865f88ef888f8;
    inBuf[2164] = 256'h7df871f836f8fbf7cbf77ff73ff716f7dff6b5f69af66cf643f61af6d2f588f5;
    inBuf[2165] = 256'h3ef5e0f489f443f4fbf3caf3b0f394f387f38af381f378f372f35cf345f336f3;
    inBuf[2166] = 256'h21f319f326f339f361f39cf3d4f319f463f498f4d2f40ff534f560f598f5c3f5;
    inBuf[2167] = 256'h00f654f69bf6f0f655f7a2f7eff73ef866f88cf8b4f8b4f8b9f8cef8c5f8c8f8;
    inBuf[2168] = 256'he4f8e4f8eaf801f9f1f8daf8c6f882f836f8f2f785f716f7bbf645f6d7f580f5;
    inBuf[2169] = 256'h11f5a8f44ff4d3f355f3e1f246f2a4f10ff15df0abef10ef68eecded4bedbfec;
    inBuf[2170] = 256'h44ecddeb65ebf4ea8eea14eaa1e93ae9c4e85ee80fe8bfe788e76de755e758e7;
    inBuf[2171] = 256'h72e788e7afe7e3e70ce841e87fe8b5e8fee853e9a8e91deaa4ea2bebd2eb8aec;
    inBuf[2172] = 256'h38edfaedbeee71ef37f0f9f0a7f16bf232f3e5f3b3f48ff559f636f715f8ddf8;
    inBuf[2173] = 256'hb3f981fa2cfbdffb8bfc14fda7fd37fea9fe2affacff10007b00e20024016701;
    inBuf[2174] = 256'ha101b401c601d401c001ad019a016c0142011a01db009d0060000e00b8ff61ff;
    inBuf[2175] = 256'hfcfe94fe29feb3fd3efdcbfc53fce0fb6efbfdfa96fa36fad9f981f930f9e9f8;
    inBuf[2176] = 256'ha8f869f837f80bf8e2f7caf7bbf7b4f7c6f7e9f714f854f8a3f8f5f857f9c2f9;
    inBuf[2177] = 256'h2afa9ffa18fb8dfb13fca6fc36fdd8fd8dfe41ff0300d00096015e022903e503;
    inBuf[2178] = 256'h9b045405ff05a1064907ea0786082709c109500ade0a620bda0b480ca50cf30c;
    inBuf[2179] = 256'h3a0d6e0d920dad0db50dac0d9c0d830d5b0d280def0cb10c6a0c1d0ccc0b6d0b;
    inBuf[2180] = 256'h040b990a1b0a92090c097908dd074f07c0063306bc054505d004700407049803;
    inBuf[2181] = 256'h3b03d1025d0201029f013e010701da00b400ba00c700d5000701350157019401;
    inBuf[2182] = 256'hce01f9013f028d02da024c03ca034804eb0497053606e80699073808e2088a09;
    inBuf[2183] = 256'h230aca0a740b160cc70c7c0d250ed40e7e0f1510a8102b119b1108126412b012;
    inBuf[2184] = 256'hff1246137d13b513e413051420142b1424141614f413c2138e134a13f712a812;
    inBuf[2185] = 256'h4e12e911891119119e102a10a70f1b0f9d0e100e780df30c640cce0b500bc80a;
    inBuf[2186] = 256'h350abe094009ba085508e90773072607da0686065d0635060306ff05fd05ee05;
    inBuf[2187] = 256'h0d062b0637067306b106db0634079307e1075e08dc084509df097e0a030bb20b;
    inBuf[2188] = 256'h640cfc0cba0d790e1f0fe80fb31067113c121013cb13a21473152716f216b217;
    inBuf[2189] = 256'h5118ff18a019211aaf1a321b9c1b141c7c1cce1c351d8e1dcb1d141e491e611e;
    inBuf[2190] = 256'h811e891e721e641e401e031ed51d941d421d071db91c571c101cb41b411be41a;
    inBuf[2191] = 256'h6f1adf196719d9183518b31720177c1602167f15ef148e142014a5135513f212;
    inBuf[2192] = 256'h7b123112d41165112511db1087106c104b10221031103810301056106c106d10;
    inBuf[2193] = 256'h9110a1109f10c410de10f21038117d11bc1127128c12e1125113ac13e9132b14;
    inBuf[2194] = 256'h5414671488149a14a214c714e7140115311558156b1582157c1554152615dd14;
    inBuf[2195] = 256'h7a141b14b1134213e8128a122912d611761105119110fb0f4a0f980ec80de80c;
    inBuf[2196] = 256'h1b0c490b7b0ad2092c098c080f088a07ff068806f8055705cc042b048103fc02;
    inBuf[2197] = 256'h7502f201a4015d011d010d01fe00ee0002010a0107012301340137015d018001;
    inBuf[2198] = 256'h9f01e80137028602000384030404a7044b05e1058f063707c5076308f9087709;
    inBuf[2199] = 256'h080a9a0a1e0bbb0b610cfb0caa0d5d0efa0e9c0f3110a61017117411af11eb11;
    inBuf[2200] = 256'h24124e128712ca120c136013b81303144b147d14921493146c142514d5137213;
    inBuf[2201] = 256'h0713ab124f120112cd11951161113711f110911023108e0fe20e2e0e600d990c;
    inBuf[2202] = 256'heb0b3f0bab0a3d0acd09690913099f081a088e07d7060b06420567049603ea02;
    inBuf[2203] = 256'h4902c70171012501eb00bc0076002200c6ff43ffb2fe24fe8cfd03fd9bfc4afc;
    inBuf[2204] = 256'h1bfc10fc15fc2afc43fc4dfc4afc2cfcf3fbb2fb60fb04fbbafa7bfa4cfa3ffa;
    inBuf[2205] = 256'h40fa4dfa6dfa7ffa86fa8bfa6efa3bfa04fab1f956f90cf9b3f863f82df8edf7;
    inBuf[2206] = 256'hb4f78ef74df705f7c2f65df6e8f575f5e4f451f4cdf335f3a5f22ef2acf139f1;
    inBuf[2207] = 256'hdef074f010f0beef57efefee90ee19eea0ed2ceda6ec28ecc0eb56eb02ebccea;
    inBuf[2208] = 256'h99ea80ea84ea86ea95eaafeabceaceeae3eae6eaf3ea0feb25eb54eb9febf3eb;
    inBuf[2209] = 256'h64eceeec76ed0deeaaee2eefb3ef33f096f0fbf065f1c2f135f2bbf240f3e4f3;
    inBuf[2210] = 256'h99f43df5f1f5a3f62ef7b7f731f87cf8c9f816f945f985f9d8f91dfa7dfaf0fa;
    inBuf[2211] = 256'h49fba8fb05fc33fc52fc64fc44fc1afcedfba2fb62fb3dfb0dfbf4faf7faedfa;
    inBuf[2212] = 256'hecfaf5fadafab0fa80fa24fab9f953f9d2f850f8e8f77bf71ff7dff697f653f6;
    inBuf[2213] = 256'h1cf6c8f56af510f594f40cf48df3fcf273f20af29af13af102f1c2f084f05cf0;
    inBuf[2214] = 256'h21f0deefa4ef4defebee94ee29eec5ed78ed22eddcecb5ec81ec5dec54ec37ec;
    inBuf[2215] = 256'h1fec1becfbebddebd1ebaaeb88eb78eb4feb36eb39eb28eb29eb49eb54eb72eb;
    inBuf[2216] = 256'habebc4ebe4eb14ec1bec23ec38ec25ec18ec1dec06ec05ec22ec2cec4eec87ec;
    inBuf[2217] = 256'ha2ecccecffec02ed0aed16edf5ecddecd6ecb1eca4ecb3ecacecbdece3eceaec;
    inBuf[2218] = 256'hf8ec0bedf5ecddecc2ec86ec59ec3dec13ec05ec13ec1dec46ec82ecaaecdeec;
    inBuf[2219] = 256'h13ed2aed45ed5eed60ed71ed8eeda3edd5ed1cee63eec6ee37ef9bef0ef084f0;
    inBuf[2220] = 256'he7f056f1c5f124f293f20cf37bf302f497f423f5c5f56ef603f7a4f746f8cbf8;
    inBuf[2221] = 256'h55f9ddf948fab8fa28fb84fbedfb5afcb3fc1afd86fddafd38fe95fed4fe13ff;
    inBuf[2222] = 256'h49ff5eff73ff86ff7dff75ff70ff5eff56ff54ff41ff35ff2cff0dffe8fec0fe;
    inBuf[2223] = 256'h80fe36fee7fd89fd2cfdd6fc7bfc2dfcf0fbb3fb7bfb52fb29fbfdfad4faa8fa;
    inBuf[2224] = 256'h7afa4ffa20faf4f9d2f9b4f99bf98ff986f980f981f980f980f985f988f98af9;
    inBuf[2225] = 256'h92f999f9a6f9b9f9ccf9e9f90efa33fa5ffa90fabffaf3fa27fb53fb83fbb0fb;
    inBuf[2226] = 256'hcffbeffb0dfc1afc29fc3bfc42fc4dfc5dfc67fc79fc8efc98fca6fcb6fcb6fc;
    inBuf[2227] = 256'hb3fcaffca0fc8efc82fc71fc64fc5efc5afc5dfc63fc64fc66fc65fc59fc49fc;
    inBuf[2228] = 256'h38fc1ffc07fcf5fbe5fbddfbddfbe2fbeefbfafb07fc19fc28fc33fc44fc53fc;
    inBuf[2229] = 256'h63fc7efc9cfcc0fcf3fc27fd5efd9ffddbfd17fe59fe95fecdfe0bff44ff80ff;
    inBuf[2230] = 256'hc2fffdff40008f00d70025018101d90133029902fa025f03c80329048b04ef04;
    inBuf[2231] = 256'h44059905ef053a068606d80623077407ca071a086e08c208070946098109b009;
    inBuf[2232] = 256'hda09fe09190a390a5a0a760a960ab60ace0ae40af20aed0adc0ac10a990a680a;
    inBuf[2233] = 256'h2e0aee09b20974093409fa08ba0872082c08d8077c072507c0065506fa059b05;
    inBuf[2234] = 256'h3c05f004a0044c040b04c50377033603ec02980259021902d601ae0189016401;
    inBuf[2235] = 256'h5a01510144014c01530155016b0181019701c601f9012d027d02d10223038603;
    inBuf[2236] = 256'he40337049704ef0437058905da0520066d06bc06050752079907d50715085108;
    inBuf[2237] = 256'h7f08ad08d808f80818093109410950095a0955094d093c091b09fa08d4089f08;
    inBuf[2238] = 256'h6b083608f607b90779072e07e40694063b06e40589052a05da048b043a040104;
    inBuf[2239] = 256'hcf039c037c035b03370326031003ef02e202d502bf02c002c602ca02e6020403;
    inBuf[2240] = 256'h1f0353038b03b803f8033a047004b904060549059d05f6054506a10601075807;
    inBuf[2241] = 256'hbb071e087508d3082e097b09cc09170a510a8d0ac30ae90a110b360b500b6f0b;
    inBuf[2242] = 256'h8a0b9d0bb20bbd0bbc0bbc0bb30b9a0b800b5c0b2f0b080bdf0ab20a8c0a620a;
    inBuf[2243] = 256'h300a030ace098c094809fa08a1084b08ed078f074007f206a90672063906fe05;
    inBuf[2244] = 256'hce0592054e051205cc047c043904f803bc03950370034f0341032e0314030603;
    inBuf[2245] = 256'heb02c102a2027b024b022e02170204020b021b022e0258028302a402ce02f102;
    inBuf[2246] = 256'h070325033a0343035a0372038403a803d60302043b047404a804e70423055205;
    inBuf[2247] = 256'h8505b505d705fc052106450670069b06c406f506260753078307ac07cc07e907;
    inBuf[2248] = 256'hf807f807f407e707cf07b907a2078a07780768075607470733071807fc06d106;
    inBuf[2249] = 256'h9b0669063006f305c505960567054f053d05280521051605ff04f204db04b504;
    inBuf[2250] = 256'h99047a0454044304380430043f04530468049104ba04dc040c0539055d058f05;
    inBuf[2251] = 256'hbe05e705230662069e06e5062b076d07b407f10723085b088608a108be08d508;
    inBuf[2252] = 256'he308f308fe08060914091f0924092509200915090109df08b60883083f08f507;
    inBuf[2253] = 256'ha7074f07f4069d064006eb059b054205e80496043904d2036903f3027a020702;
    inBuf[2254] = 256'h8e011901b5005500fdffbdff81ff48ff21fffbfed1feaffe8afe63fe48fe2cfe;
    inBuf[2255] = 256'h14fe11fe14fe1bfe38fe5afe7ffeb3fee8fe17ff4eff83ffb1ffe5ff1c005300;
    inBuf[2256] = 256'h9400d7001c016b01bc0109025902a502e90227035d038803ad03c703d903ee03;
    inBuf[2257] = 256'h00040e041f042f043f0451045e04620461045b044b042f040c04e303b3037d03;
    inBuf[2258] = 256'h48031503e202b20285025a022d02fe01cb01920157011a01dd00a10067003500;
    inBuf[2259] = 256'h0f00edffcdffb9ffabff9aff8aff7bff69ff57ff42ff2eff24ff1dff1bff26ff;
    inBuf[2260] = 256'h37ff4dff6bff8affa7ffc7ffe3fff7ff0a001b002b0042005a0075009a00c500;
    inBuf[2261] = 256'hf5002c0163019901cf0101022d0251026c02830295029e02a602ae02b302b802;
    inBuf[2262] = 256'hbb02be02c402c202ba02b302a4028d02740250022702ff01ce019a016b013601;
    inBuf[2263] = 256'hff00cc008d0048000700bbff64ff0effaffe4afeedfd89fd22fdc7fc6dfc10fc;
    inBuf[2264] = 256'hbbfb61fb03fbadfa54faf4f99bf93ff9e3f897f84bf802f8c8f792f75ff73cf7;
    inBuf[2265] = 256'h1bf7f7f6def6c9f6b3f6a6f69bf690f68cf68cf691f69ff6adf6bff6d8f6f0f6;
    inBuf[2266] = 256'h10f73cf764f793f7cff70cf84df895f8d7f81df966f9a4f9e6f928fa5cfa95fa;
    inBuf[2267] = 256'hd4fa01fb32fb69fb8ffbb7fbe3fb01fc23fc47fc5afc73fc8efc93fc9bfca8fc;
    inBuf[2268] = 256'ha0fc99fc8ffc6cfc49fc28fceefbb7fb8bfb50fb16fbe8fab0fa7ffa54fa1afa;
    inBuf[2269] = 256'he2f9aff96df92bf9eef8a5f85ff81ff8d7f798f762f728f7f9f6d2f6a3f67ff6;
    inBuf[2270] = 256'h67f649f633f627f61bf61af620f622f631f643f64cf661f67df68ff6aaf6cef6;
    inBuf[2271] = 256'he9f60ff73ff769f79bf7d7f709f842f880f8b2f8e7f823f950f97ff9b2f9d6f9;
    inBuf[2272] = 256'hfaf924fa3cfa4ffa68fa73fa7dfa8bfa89fa8cfa98fa95fa94fa99fa8bfa7dfa;
    inBuf[2273] = 256'h75fa5afa39fa1cfaecf9b8f98cf94ef90ef9d7f892f84ef815f8ccf784f746f7;
    inBuf[2274] = 256'hfff6bef68df651f618f6ecf5baf58cf564f52df5f9f4c9f48df455f425f4f2f3;
    inBuf[2275] = 256'hccf3b6f3a0f39df3a9f3b0f3c2f3def3edf3fff312f416f420f42ef432f441f4;
    inBuf[2276] = 256'h5af46df48df4bbf4e4f416f54ff57ff5b9f5f6f528f662f6a1f6d4f612f754f7;
    inBuf[2277] = 256'h88f7c3f7fff729f859f889f8a6f8c6f8e8f8f8f812f932f947f968f990f9a9f9;
    inBuf[2278] = 256'hcff9fff91dfa40fa65fa78fa8bfa9afa94fa94fa95fa82fa76fa72fa67fa67fa;
    inBuf[2279] = 256'h70fa72fa81fa98faa2fab1fabefabbfabafab6faa1fa91fa81fa68fa56fa4cfa;
    inBuf[2280] = 256'h3efa3cfa40fa3dfa43fa4dfa4bfa50fa5dfa64fa73fa89fa9cfab9faddfafcfa;
    inBuf[2281] = 256'h1cfb39fb4bfb5dfb6cfb70fb75fb7afb7dfb8bfba3fbc1fbf0fb29fc62fca7fc;
    inBuf[2282] = 256'heffc2ffd70fdaafdd1fdf7fd18fe2afe39fe47fe4ffe62fe7cfe90feadfed4fe;
    inBuf[2283] = 256'hf6fe1dff4bff6cff87ffa3ffb8ffc2ffc4ffbeffb5ffa6ff90ff7dff6cff56ff;
    inBuf[2284] = 256'h42ff32ff1fff0cfffafee8fed7fec7feb6fea7fe9afe8dfe83fe7bfe71fe64fe;
    inBuf[2285] = 256'h52fe40fe2cfe12fef6fddbfdc1fdaefda3fda1fdb0fdcbfdedfd1bfe50fe84fe;
    inBuf[2286] = 256'hbbfef0fe1cff43ff65ff81ff9dffb5ffccffeeff180045007e00c3000d015d01;
    inBuf[2287] = 256'hb10106025c02ae02f8023f038303c003f503270457048104a504c604e7040105;
    inBuf[2288] = 256'h17052d0543055405680581059a05b805db05fa051b063b065406670671066b06;
    inBuf[2289] = 256'h5b063f061806f005c40593056f0553053c0539053e05420555056b0577058705;
    inBuf[2290] = 256'h8d05810578056805480530051805fd04f604f404f0040405200538055f058805;
    inBuf[2291] = 256'haa05d405fa0516063c065b066e068e06a806b706d106e606f00608071e072a07;
    inBuf[2292] = 256'h43075d0773079b07c607ee0726085f089208cf0805092c09520969096e097209;
    inBuf[2293] = 256'h68094f093c0925090909fc08f308ed08fc080e091d093e09570964097a098709;
    inBuf[2294] = 256'h81097e096f09500939091709e908ca08a60879085f08460827081d0812080208;
    inBuf[2295] = 256'h08080b0805081008120808080c080308e907dd07c807a4079307810769076807;
    inBuf[2296] = 256'h69076a078607a507c007f40727084e088608b608d60802092309330953096909;
    inBuf[2297] = 256'h71098b09a409b809e609150a400a870ad20a120b660bb60bf30b3a0c780ca30c;
    inBuf[2298] = 256'hd20cf00cfb0c100d1c0d190d240d290d230d2f0d3a0d3c0d4d0d5a0d600d760d;
    inBuf[2299] = 256'h820d830d8e0d890d720d650d450d100de10ca40c580c190cd00b800b470b0a0b;
    inBuf[2300] = 256'hc90aa20a7b0a4f0a380a1e0afa09e709cb09a3098b09670935091209e308a808;
    inBuf[2301] = 256'h800851081c080208e807cd07d307da07df0703082808450876089f08b608d808;
    inBuf[2302] = 256'hee08f508070910091109250939094c097709a109c709030a3b0a6b0aa80adb0a;
    inBuf[2303] = 256'h020b320b530b630b770b7b0b6e0b680b560b380b240b080be80ad60ac00aab0a;
    inBuf[2304] = 256'ha70a9d0a8f0a8d0a820a6b0a560a310afd09cc098c094109fb08a6084b08fe07;
    inBuf[2305] = 256'ha7074e070907c0067a064c061c06ef05da05c205a6059b058705680554053305;
    inBuf[2306] = 256'h0305df04b1047e045e043f041f04190419041a0431044c0465048e04b504d404;
    inBuf[2307] = 256'hfd04200539055b0578058e05ab05c105d305ec05000610062906450663068c06;
    inBuf[2308] = 256'hb906e6061a074a0773079b07b807c907d307cd07b907a30782075b0734070807;
    inBuf[2309] = 256'hdd06bb069b067c06630647062d061706f905d405ad057b053c05f504a1044304;
    inBuf[2310] = 256'hdd036c03fd0291022202be0163010d01c500840042000800d0ff8eff4eff0eff;
    inBuf[2311] = 256'hc4fe7bfe32fee0fd95fd4ffd04fdc1fc87fc4bfc13fce7fbbffb9ffb88fb7bfb;
    inBuf[2312] = 256'h77fb79fb83fb95fba8fbbafbcbfbd5fbddfbe1fbdcfbd8fbd9fbd9fbdefbeffb;
    inBuf[2313] = 256'h05fc21fc47fc70fc9dfccefcf9fc26fd50fd6bfd84fd9bfda4fda9fdacfda0fd;
    inBuf[2314] = 256'h93fd89fd74fd62fd56fd42fd33fd2efd20fd13fd0afdf4fcd9fcbbfc8dfc5afc;
    inBuf[2315] = 256'h22fcd6fb86fb38fbdafa7afa21fabbf95af905f9a8f852f80cf8c1f77ff74df7;
    inBuf[2316] = 256'h15f7dff6b6f680f643f609f6bff56cf51df5bff462f415f4c8f385f35af335f3;
    inBuf[2317] = 256'h21f324f322f327f33cf348f352f362f365f36bf37af37df389f3a2f3aef3c3f3;
    inBuf[2318] = 256'heaf300f41bf444f45af478f4a7f4c0f4e3f419f539f55ef591f5a8f5c4f5e8f5;
    inBuf[2319] = 256'hecf5eef5f8f5e3f5d2f5cff5aff596f592f574f55ef55df545f533f530f513f5;
    inBuf[2320] = 256'hf7f4e6f4b2f47cf44df4fcf3a8f35ff3f9f297f248f2e8f191f154f109f1cdf0;
    inBuf[2321] = 256'ha6f06ef03ef01ff0e6efaeef80ef3aeff8eec5ee7bee3bee0eeeceed98ed78ed;
    inBuf[2322] = 256'h45ed18ed00edd8ecbbecb6eca0ec96eca8ecacecbcece0ecefec02ed20ed24ed;
    inBuf[2323] = 256'h2aed3eed38ed3bed4fed52ed64ed8deda9edd8ed1cee4dee8aeed2eefdee2eef;
    inBuf[2324] = 256'h6aef87efaaefd6efe1eff6ef1bf027f03ff06bf07ef0a0f0d6f0f3f01bf153f1;
    inBuf[2325] = 256'h6df18af1b2f1b9f1c1f1d5f1caf1c4f1cef1c2f1c0f1ccf1bff1bff1cff1c4f1;
    inBuf[2326] = 256'hbff1c6f1b1f1a2f19df184f179f181f171f16ef17af16df165f166f14af12ef1;
    inBuf[2327] = 256'h17f1e4f0bbf0a3f07df06cf073f070f07ff0a6f0c0f0e0f009f11ef131f145f1;
    inBuf[2328] = 256'h3ff13ff147f13ef141f152f157f170f19cf1baf1e4f11df248f27df2bcf2e7f2;
    inBuf[2329] = 256'h1bf358f37ff3adf3e4f308f434f469f48af4b5f4eaf410f540f578f59af5c8f5;
    inBuf[2330] = 256'h02f624f651f688f6a9f6d5f60af728f74cf77af790f7a8f7c1f7c1f7c5f7cdf7;
    inBuf[2331] = 256'hc3f7c5f7d4f7d8f7ecf70ff829f854f887f8a5f8c5f8e5f8ecf8f1f8f1f8def8;
    inBuf[2332] = 256'hd0f8c8f8b7f8b5f8bff8c3f8d3f8eff802f91bf937f94bf966f982f996f9b2f9;
    inBuf[2333] = 256'hd2f9ecf910fa38fa55fa76fa97faaffaccfaeafafffa1cfb3ffb62fb8ffbc2fb;
    inBuf[2334] = 256'hf4fb2efc6bfca3fcdffc18fd4afd7ffdaffddbfd08fe2ffe53fe7efea5fec8fe;
    inBuf[2335] = 256'hf4fe24ff56ff90ffcdff10005c00a500ec00300169019a01c401e101fa011002;
    inBuf[2336] = 256'h1f0233024f026c029102bf02ee0224035d038d03be03ee031204360459047204;
    inBuf[2337] = 256'h8e04a704b604cb04dd04e304ef04fa04fc040605140520053d055d057905a405;
    inBuf[2338] = 256'hcf05ed05120630063b064d0659065206510651064a06510658065c0674068c06;
    inBuf[2339] = 256'h9c06bf06e60603072d07550774079f07c607df0700081808220835083f083f08;
    inBuf[2340] = 256'h5208650873089608bc08e1081a094e097709b109e4090a0a3d0a660a810aab0a;
    inBuf[2341] = 256'hcd0ae20a080b250b310b4c0b600b660b830b9e0bad0bd60b080c2f0c680ca10c;
    inBuf[2342] = 256'hcb0c030d2e0d400d560d5d0d4c0d470d390d1d0d180d170d110d240d350d3e0d;
    inBuf[2343] = 256'h640d850d970dbd0dd80de40d060e1e0e220e3a0e440e390e3e0e370e1d0e1b0e;
    inBuf[2344] = 256'h120efc0d050e110e150e3c0e670e860ebf0ef30e140f460f6a0f770f950fa70f;
    inBuf[2345] = 256'ha20fb50fc40fc30fdc0ff10ffc0f241047105c109010c110e1101b114a116111;
    inBuf[2346] = 256'h9011af11af11c311cb11b911bb11b511a011a611a8119e11b111be11bb11d011;
    inBuf[2347] = 256'hda11cf11da11d711c011c011b0118f1186116f1142112811fb10bd1093105810;
    inBuf[2348] = 256'h0e10e10fb00f7d0f6e0f5c0f460f4f0f500f400f430f320f090fee0ec10e7f0e;
    inBuf[2349] = 256'h530e1f0ee20dc20da00d7b0d780d730d650d750d800d7f0d960da50da70dba0d;
    inBuf[2350] = 256'hbf0db50dbd0db60d9b0d960d870d6b0d6a0d670d5a0d6d0d800d8b0db20dd40d;
    inBuf[2351] = 256'he50d070e1e0e200e300e320e1f0e180e050ee60dd70dbb0d940d830d660d410d;
    inBuf[2352] = 256'h370d2a0d140d190d190d0f0d190d170d060dff0ce30cb10c8c0c520c050cce0b;
    inBuf[2353] = 256'h8f0b480b1e0bf40ac90abc0aac0a930a930a880a6f0a6b0a5d0a3d0a2f0a180a;
    inBuf[2354] = 256'hf309da09b90991097809510922090909eb08ca08c108b808b208c608d508e208;
    inBuf[2355] = 256'h05091f0930094b09570957095f0955093f09370925090b09ff08ec08d608d608;
    inBuf[2356] = 256'hd608d508e708f90809092809430950095d095f094f0939091109de08aa086e08;
    inBuf[2357] = 256'h33080408d207a7079007790761075707440725070907e306ad0675063206e705;
    inBuf[2358] = 256'h9c054905f404a60452040004b7036d032503e802a90274024b021d02f401d301;
    inBuf[2359] = 256'haa0180015b012801f000bc007c003d000500c5ff8aff5dff2eff08fff4fee2fe;
    inBuf[2360] = 256'hd9fedefee2feedfe02ff12ff23ff39ff45ff4cff55ff54ff4cff44ff3aff32ff;
    inBuf[2361] = 256'h31ff33ff3cff4dff64ff82ffa3ffc2ffdffff7ff090016001800170013000500;
    inBuf[2362] = 256'hf5ffe8ffd3ffbcffa9ff8fff73ff5bff3dff20ff06ffe7fecbfeb8fe9dfe7ffe;
    inBuf[2363] = 256'h66fe43fe19feedfdb5fd75fd33fdeafc9dfc57fc12fcd2fb9ffb75fb53fb3efb;
    inBuf[2364] = 256'h2efb22fb1afb0ffb03fbf4fadcfabcfa9afa72fa48fa22fafef9dff9cbf9c1f9;
    inBuf[2365] = 256'hc2f9d0f9e5f901fa28fa4ffa77fa9dfab9fad3faecfaf8fa00fb0cfb0ffb15fb;
    inBuf[2366] = 256'h24fb29fb33fb48fb51fb5ffb77fb81fb8afba0fba7fbb0fbc6fbc9fbcafbd5fb;
    inBuf[2367] = 256'hcbfbbcfbb1fb8dfb64fb41fb07fbc9fa97fa56fa1afaeef9bbf98ff971f945f9;
    inBuf[2368] = 256'h1ef900f9cff89bf86ef82bf8e0f79bf744f7edf6a1f64cf600f6c4f581f547f5;
    inBuf[2369] = 256'h21f5f7f4d3f4bdf49ef481f46ff453f435f41ef4fdf3dff3c6f3a1f382f370f3;
    inBuf[2370] = 256'h55f341f33ff335f335f347f352f36af395f3b5f3dff318f446f476f4acf4cef4;
    inBuf[2371] = 256'hf1f416f522f530f545f545f54ff568f573f58af5b2f5d2f503f642f66df6a1f6;
    inBuf[2372] = 256'hdcf6fef620f740f741f743f747f730f71ef715f7f8f6e4f6dcf6c4f6baf6bdf6;
    inBuf[2373] = 256'hacf6a0f69cf683f66cf65bf632f60df6eff5baf58af566f531f503f5e1f4acf4;
    inBuf[2374] = 256'h7ff460f42ff404f4e9f3c1f3a1f390f376f363f35ef34df343f344f336f329f3;
    inBuf[2375] = 256'h26f316f308f304f3f6f2f2f2faf200f314f334f351f382f3bef3ecf322f462f4;
    inBuf[2376] = 256'h91f4c4f4fbf41ef544f570f58af5a7f5cff5ecf510f63ef663f68ef6c3f6eef6;
    inBuf[2377] = 256'h1ff758f780f7a8f7d3f7e7f7fbf712f812f812f816f806f8f8f7f2f7d7f7c2f7;
    inBuf[2378] = 256'hb9f79ef788f77cf75ef746f736f711f7f2f6dcf6aef681f65ff628f6f0f5c1f5;
    inBuf[2379] = 256'h82f547f517f5daf4a5f481f456f437f426f40bf4fdf3f9f3e4f3d5f3cdf3b3f3;
    inBuf[2380] = 256'h9ff393f375f35ef355f347f344f34ef352f369f38ef3acf3d7f30ef439f470f4;
    inBuf[2381] = 256'hadf4d9f40df546f56bf597f5c9f5e8f511f642f665f693f6cdf6faf631f775f7;
    inBuf[2382] = 256'habf7ecf733f869f8a6f8ebf81af94ef988f9abf9cff9f8f90cfa22fa39fa3cfa;
    inBuf[2383] = 256'h44fa4ffa49fa49fa53fa53fa5efa72fa7bfa8dfaa1faa7fab3fabdfaaefa9efa;
    inBuf[2384] = 256'h8dfa68fa44fa23faf5f9cff9b2f98ff979f971f962f95af95af950f94bf94af9;
    inBuf[2385] = 256'h3cf931f926f90ef9faf8e8f8cbf8b5f8a7f893f887f88bf88ef89bf8b0f8c6f8;
    inBuf[2386] = 256'he8f811f933f959f983f9a7f9ccf9eef906fa24fa44fa5cfa78fa96fab2fad8fa;
    inBuf[2387] = 256'h00fb25fb55fb8bfbbefbfcfb3efc79fcbdfc03fd3dfd79fdb1fdd9fdfefd1ffe;
    inBuf[2388] = 256'h2ffe3efe4cfe52fe5cfe6dfe7afe8bfea5febafed4fef1fe05ff18ff28ff2cff;
    inBuf[2389] = 256'h2cff29ff17ff04fff0fed2feb4fe98fe77fe5bfe43fe27fe0ffefcfde6fdd5fd;
    inBuf[2390] = 256'hc4fdaffd9efd8ffd7afd64fd4efd33fd18fdfdfce4fccdfcb6fca6fc9cfc93fc;
    inBuf[2391] = 256'h90fc93fc98fca9fcc2fcdafcf6fc18fd3bfd5cfd7dfd9afdb6fdd3fde9fdf9fd;
    inBuf[2392] = 256'h0cfe21fe39fe56fe7dfeaffee9fe28ff6cffbbff090051009900da000b013801;
    inBuf[2393] = 256'h5f0177018c01a301b501c901e001f9011a023c025c028402ac02cc02ef021103;
    inBuf[2394] = 256'h2a0341035403600369036a0365035f03520340032d031403fd02ea02d502c802;
    inBuf[2395] = 256'hbf02b402b302ba02bc02c002c502c502c502bf02b002a00287026a0254023b02;
    inBuf[2396] = 256'h200211020502fd0104020f0220023e025a0274029702b202c702e002ee02f402;
    inBuf[2397] = 256'hff02030302030c03170322033c035a037703a103d203ff03330468049904cd04;
    inBuf[2398] = 256'hfe042705520576059005ab05c005ce05df05ed05f105fe05100621063b065906;
    inBuf[2399] = 256'h7a06a606d006f606280752076c078a07a007a507aa07a4079007820772075a07;
    inBuf[2400] = 256'h4b073f07340738073b073e0750076007690779078207830785077b0768075d07;
    inBuf[2401] = 256'h460726071007f706db06cf06c106b306b706ba06b906c806d206d406e406f106;
    inBuf[2402] = 256'hef06f506fa06f806fd06f906ed06f206f306ee06f906000703071b0732074507;
    inBuf[2403] = 256'h6c079207af07db0701081d0844085f086c088408930893089f08a708a808bb08;
    inBuf[2404] = 256'hcd08db08fe08220941096b098f09ad09d609f609080a1f0a2e0a2e0a330a310a;
    inBuf[2405] = 256'h270a280a220a160a190a170a100a1d0a280a2d0a410a510a590a6c0a760a730a;
    inBuf[2406] = 256'h7b0a780a670a600a500a370a2a0a180a010afd09f409e709f009f309f109030a;
    inBuf[2407] = 256'h100a130a250a2f0a2e0a3b0a3d0a320a370a320a230a240a1c0a0d0a140a170a;
    inBuf[2408] = 256'h130a230a330a3d0a580a6d0a7b0a960aa60aaa0abb0ac00aba0ac10abe0ab10a;
    inBuf[2409] = 256'hb50ab40aab0aba0ac40ac90ae70a010b110b350b530b660b870b9e0ba40bb70b;
    inBuf[2410] = 256'hbf0bb90bbf0bba0bac0bb10bb00ba80bb70bc50bca0be40bfc0b0c0c2d0c460c;
    inBuf[2411] = 256'h530c700c840c8b0ca10ca90ca10caa0caa0c970c920c890c740c6e0c610c4b0c;
    inBuf[2412] = 256'h4d0c4b0c420c4c0c510c4c0c590c5b0c4f0c500c400c1c0c0b0cef0bc00ba30b;
    inBuf[2413] = 256'h800b530b3c0b200bfc0af00ae10ac70ac30ab80a9e0a950a800a5f0a500a320a;
    inBuf[2414] = 256'h060aee09d009a7099309790959094e093d092a092e092b0922092e0933093009;
    inBuf[2415] = 256'h410945093d0947094a0943094c094b094009440945093e094409480949095709;
    inBuf[2416] = 256'h62096d098909a109b309d109e809f6090a0a130a100a140a0b0af809ef09db09;
    inBuf[2417] = 256'hc309bc09b209a309a509a509a109a809a4099609940984096609510932090709;
    inBuf[2418] = 256'he308b9088808610832080108dd07b00781075f0731070107e006b7068c066c06;
    inBuf[2419] = 256'h44061b06fd05d405aa058c05620532051005e404b40492046c0444042b041304;
    inBuf[2420] = 256'hfa03ef03e703dd03dd03da03d403d403ce03bf03b703ae039e0394038f038b03;
    inBuf[2421] = 256'h91039903a403ba03d203ea0306041e04310442044f0457045e045c0457045804;
    inBuf[2422] = 256'h54044e044f044a0442043d0433042804230416040604f903e803d603c303ab03;
    inBuf[2423] = 256'h9203760350032903f902be0283024502fc01b50170012501dd00990055001800;
    inBuf[2424] = 256'hddffa1ff6aff30fff1feb3fe70fe26fedefd95fd48fdfffcb7fc6efc2bfceefb;
    inBuf[2425] = 256'hb6fb85fb57fb2dfb0afbe8fac8faaefa94fa77fa5ffa47fa2efa1cfa09faf5f9;
    inBuf[2426] = 256'heaf9e3f9dcf9dcf9def9e1f9ebf9f5f905fa1bfa2bfa3efa5bfa6ffa82fa9dfa;
    inBuf[2427] = 256'haefabbfad0fadafae0faeafaeafae7faebfae5fae2fae9fae6fae4faedfaebfa;
    inBuf[2428] = 256'he8faecfae0fad2fac8faabfa8bfa6efa3cfa09fae1f9a8f96df93df902f9ccf8;
    inBuf[2429] = 256'ha1f868f835f80ef8d9f7a7f77ff744f70cf7e2f6a4f663f630f6eff5aff57af5;
    inBuf[2430] = 256'h3bf500f5d5f4a0f46ff44df422f400f4edf3d1f3bff3b9f3a5f39af3a0f395f3;
    inBuf[2431] = 256'h8ef397f38ff38bf397f393f395f3a8f3abf3b6f3d1f3e1f3faf324f440f463f4;
    inBuf[2432] = 256'h92f4aef4cef4fcf414f52bf54bf557f568f582f587f595f5aef5b3f5c2f5dff5;
    inBuf[2433] = 256'he4f5f2f50cf60bf60ff620f616f60ef610f6f3f5d7f5c8f59ef576f55bf526f5;
    inBuf[2434] = 256'hf6f4d5f4a0f470f44ef419f4ecf3cff39bf36ff351f31bf3eaf2c8f28ff25af2;
    inBuf[2435] = 256'h31f2f2f1b9f191f155f11ef1f8f0c4f099f07ef056f03bf032f019f00bf00ff0;
    inBuf[2436] = 256'h05f000f00af004f006f013f011f015f025f027f035f051f05ef077f09ef0baf0;
    inBuf[2437] = 256'he2f019f13df16cf1a8f1cff1fcf134f257f282f2b6f2d2f2f6f225f33ff366f3;
    inBuf[2438] = 256'h98f3b1f3d8f30bf423f446f477f48df4adf4d9f4e7f4faf41bf521f52af53cf5;
    inBuf[2439] = 256'h35f534f53bf52bf523f523f50df504f507f5f2f4e9f4eef4dff4d7f4d9f4c9f4;
    inBuf[2440] = 256'hc0f4bef4a7f494f489f46ef45bf44df430f41df414f400f4fdf304f4fef307f4;
    inBuf[2441] = 256'h1cf421f431f44ef45cf472f48ff49ff4b5f4d5f4e8f405f52cf547f56cf599f5;
    inBuf[2442] = 256'hbdf5edf524f64df683f6c2f6f3f62ef771f7a7f7e7f72cf85ff899f8d8f809f9;
    inBuf[2443] = 256'h44f97ff9a9f9dcf914fa39fa68fa9cfac3faf1fa24fb48fb71fb9bfbb7fbd7fb;
    inBuf[2444] = 256'hf4fb02fc14fc26fc28fc2dfc36fc34fc37fc3efc3cfc3efc44fc43fc48fc4ffc;
    inBuf[2445] = 256'h4dfc4bfc4afc43fc3cfc34fc26fc1cfc11fcfffbf4fbeafbdbfbd2fbcefbc8fb;
    inBuf[2446] = 256'hc9fbcefbd1fbdcfbecfbfbfb0ffc23fc36fc51fc6bfc82fc9dfcb7fccefceafc;
    inBuf[2447] = 256'h06fd21fd41fd64fd87fdb4fde0fd0cfe40fe74fea7fedffe14ff47ff7cffadff;
    inBuf[2448] = 256'hd9ff080033005c008700ae00d400fd0026014e017a01a601d001f8011d024402;
    inBuf[2449] = 256'h69028802a902c802dd02f3020a031b032b033d03490356036603700379038503;
    inBuf[2450] = 256'h8d039903a803b203be03ce03d903e403f003f503fd030604030405040c040704;
    inBuf[2451] = 256'h06040d040f04150420042a043d045304610478049104a104b704cd04dc04f004;
    inBuf[2452] = 256'h01050a051e0530053d0557056e057c059805b805cd05ec050e0628064c067006;
    inBuf[2453] = 256'h8d06b306d706f30619073a0750076f078b079e07b607c807d307e907fc070808;
    inBuf[2454] = 256'h1f08340843085b086f087c089308a208a808b908c208c208cc08ce08c808d108;
    inBuf[2455] = 256'hd408cc08d408d808d008d408d408c808c908c608b308ab08a208900887087c08;
    inBuf[2456] = 256'h6b0867085d084d084a084208340835082e082108250821081708220823081c08;
    inBuf[2457] = 256'h2c083708360846084f084c08590861085c0867086d086a087708800881089408;
    inBuf[2458] = 256'ha408ad08c608d908e208fa080b091209260934093a094c0959095e0970097a09;
    inBuf[2459] = 256'h7d0990099a099909a409a7099e09a309a1099309950990097e097b0975096809;
    inBuf[2460] = 256'h66095f094e0948093e09290920091309fd08f108df08c708bf08b408a1089908;
    inBuf[2461] = 256'h8d087908710864084e0844083608210818080a08f807f307e907dd07e007da07;
    inBuf[2462] = 256'hce07d307d007c507c807c407b807be07bd07b707c307c907c707d607de07df07;
    inBuf[2463] = 256'hf007f807f80707080a080608100810080808120814080e08150814080d081208;
    inBuf[2464] = 256'h0d0800080008f707e807e207d407c407c007b1079f079c079107800778076607;
    inBuf[2465] = 256'h50074707350718070207e806c806b30695066f06550637061006f105cf05a905;
    inBuf[2466] = 256'h8c056a05440529050905e604d004b7049a04890476045f0451043e042a041e04;
    inBuf[2467] = 256'h0b04f403e903d903c403b903aa0398038f038303750371036a0361035f035903;
    inBuf[2468] = 256'h5303550353035003560359035a03620367036c0377037e0383038c038f039303;
    inBuf[2469] = 256'h9b039e039f03a403a2039d039c0395038a037f037203610350033a0323030e03;
    inBuf[2470] = 256'hf402dc02c702b002990284026c02510238021d020102e301c1019f017b015201;
    inBuf[2471] = 256'h2a010101d300a8007e0050002400faffcdffa3ff7bff50ff2aff08ffe3fec0fe;
    inBuf[2472] = 256'ha1fe82fe66fe4dfe32fe1afe06feeefddbfdccfdbefdb5fdadfda6fda5fda6fd;
    inBuf[2473] = 256'ha6fdabfdb4fdbafdc2fdcafdd0fdd8fde1fde5fde9fdeffdf4fdfcfd04fe0efe;
    inBuf[2474] = 256'h1bfe26fe31fe41fe4dfe56fe64fe70fe7bfe88fe8ffe93fe99fe9bfe9bfe9cfe;
    inBuf[2475] = 256'h97fe8ffe88fe79fe66fe54fe3bfe1ffe06fee6fdc5fdabfd89fd67fd4afd24fd;
    inBuf[2476] = 256'hfefcdefcb6fc8cfc67fc3afc0dfce8fbbbfb8dfb6afb43fb1efb02fbe5facafa;
    inBuf[2477] = 256'hb2fa94fa7afa63fa45fa28fa0ffaeff9d2f9bcf9a2f98ff980f96ef965f966f9;
    inBuf[2478] = 256'h60f960f96af970f97af98af996f9a9f9c0f9d3f9eff90efa26fa42fa60fa76fa;
    inBuf[2479] = 256'h92faaefabefad4faeefafbfa0afb1ffb2dfb3ffb53fb5dfb70fb85fb8afb95fb;
    inBuf[2480] = 256'ha7fba9fbacfbb4fbaefbacfbb0fba7fba2fba5fb99fb8ffb8ffb80fb70fb65fb;
    inBuf[2481] = 256'h4bfb30fb19fbf3faccfaabfa7efa52fa2cfafbf9ccf9a5f974f946f920f9f2f8;
    inBuf[2482] = 256'hc8f8a7f87ef859f83ef81df8fff7ecf7d5f7c2f7b3f79df78cf781f76df75bf7;
    inBuf[2483] = 256'h4ef73cf72cf725f71bf716f718f719f720f72df739f74cf761f771f789f7a3f7;
    inBuf[2484] = 256'hb5f7d0f7f0f709f82bf854f875f89df8ccf8f5f826f959f980f9adf9ddf900fa;
    inBuf[2485] = 256'h24fa4cfa68fa86faa4fab9fad3faecfaf9fa0afb1efb25fb30fb3efb3efb43fb;
    inBuf[2486] = 256'h4afb46fb47fb4dfb44fb40fb40fb37fb30fb2afb18fb09fbfafadffac7fab2fa;
    inBuf[2487] = 256'h92fa75fa5bfa38fa1bfa01fadff9c5f9aff98ff977f967f94df938f92bf919f9;
    inBuf[2488] = 256'h0df908f900f9fff803f906f912f922f932f94bf965f97cf99bf9bbf9d7f9fbf9;
    inBuf[2489] = 256'h1ffa3efa65fa8cfaacfad3fafbfa1cfb44fb6efb93fbc0fbedfb14fc44fc76fc;
    inBuf[2490] = 256'ha2fcd6fc0dfd3cfd6efda1fdccfdfafd26fe49fe70fe93fea9fec1fed9fee8fe;
    inBuf[2491] = 256'hf6fe02ff07ff0dff10ff0bff09ff04fff5fee9fedcfec8feb7fea5fe8dfe79fe;
    inBuf[2492] = 256'h67fe52fe40fe30fe1dfe0ffe01feeffde0fdd4fdc3fdb1fda0fd8efd7efd6afd;
    inBuf[2493] = 256'h55fd43fd32fd1ffd10fd01fdf3fce9fce0fcd9fcd8fcd9fcddfce6fcf0fcfffc;
    inBuf[2494] = 256'h14fd2bfd45fd62fd7ffd9efdc0fde2fd07fe2cfe4efe74fe9afebbfedefe05ff;
    inBuf[2495] = 256'h26ff48ff6eff91ffb5ffdbfffdff1f00430066008800ad00cd00ee0012013301;
    inBuf[2496] = 256'h520173019201b201d401f201120231024d026b0285029902ab02bb02c502cf02;
    inBuf[2497] = 256'hd502d402d402d402cd02c702c202bb02b502b002ab02aa02a802a402a302a002;
    inBuf[2498] = 256'h9c029f02a1029f02a402a702a602ad02b402b602be02c402c502cd02d302d302;
    inBuf[2499] = 256'hdd02e502e502ed02f802fd02070312031a032a033b0346035a03710382039c03;
    inBuf[2500] = 256'hb903d003f10314043004530476049504b804d804f1040d05280539054c055f05;
    inBuf[2501] = 256'h6a0573057c0583058a058e058e059005920591059105920590058e058c058805;
    inBuf[2502] = 256'h8705830580057e05790571056c05620556054c053d052a0519050305ea04d504;
    inBuf[2503] = 256'hbb04a0048a046f0453043c0421040304eb03d203b803a50392037f0372036503;
    inBuf[2504] = 256'h5b035a03560354035a035a0358035f035f0359035a0355034b0347033e033203;
    inBuf[2505] = 256'h2e0326031c031c031a03140317031803150319031c031d0327032d032e033a03;
    inBuf[2506] = 256'h45034b035a0367036f037f038b039203a103ab03ae03b803c003c203c803cd03;
    inBuf[2507] = 256'hcd03d303d403d203d803d803d403d903dc03dd03e603ed03f203020411041e04;
    inBuf[2508] = 256'h36044b045c0476048d049d04b504ca04d804ea04fa0402050f0519051e052705;
    inBuf[2509] = 256'h2e05300538053c053d054805500552055c0567056f057e058a059305a205ac05;
    inBuf[2510] = 256'hb305c005c805cc05d505da05db05e105e305e005e205e105dc05da05d205c505;
    inBuf[2511] = 256'hbb05ab05970585056d055405400527050f05fd04e804d404c804ba04ac04a304;
    inBuf[2512] = 256'h97048a048304770467045c044e043b0429041404ff03ea03cf03b20399037c03;
    inBuf[2513] = 256'h5d03410324030703ed02d102b602a1028c027702670257024602380228021b02;
    inBuf[2514] = 256'h0f02ff01f201e701da01cd01c101b301a50199018801760164014e0138012201;
    inBuf[2515] = 256'h0801ee00d400b8009f0087006d00580043002b0017000500f2ffe3ffd5ffc4ff;
    inBuf[2516] = 256'hb8ffaeffa0ff94ff88ff78ff69ff5aff45ff30ff19fffcfee0fec4fea3fe84fe;
    inBuf[2517] = 256'h69fe4cfe33fe1dfe08fef7fde9fdd9fdccfdc2fdb6fdaefda7fd9ffd98fd95fd;
    inBuf[2518] = 256'h93fd92fd96fd9cfda2fdadfdb8fdc3fdcefdd9fde1fdebfdf5fdfbfd02fe0bfe;
    inBuf[2519] = 256'h15fe1ffe2dfe3cfe4efe63fe78fe91feaffeccfeeafe0dff2eff50ff76ff9cff;
    inBuf[2520] = 256'hc1ffeaff120037005e008300a400c400e000f7000e01220130013f014e015901;
    inBuf[2521] = 256'h640171017c01870193019c01a601ae01b301b801bc01bb01b901b801b401af01;
    inBuf[2522] = 256'hab01a6019f0198018f01830176016701550141012a011101f700db00bd009f00;
    inBuf[2523] = 256'h81006200430025000600e8ffcbffaeff95ff7dff67ff54ff44ff36ff2bff22ff;
    inBuf[2524] = 256'h1bff14ff0cff02fff8feeafedbfecafeb7fea2fe8dfe77fe63fe50fe3dfe2dfe;
    inBuf[2525] = 256'h21fe12fe04fefbfdeefddffdd4fdc5fdb6fdaafd9afd8cfd82fd75fd67fd60fd;
    inBuf[2526] = 256'h53fd43fd3afd2afd15fd03fdeafccefcb4fc92fc6efc50fc2dfc06fce5fbbdfb;
    inBuf[2527] = 256'h94fb73fb4bfb1ffbf9facefaa1fa7dfa53fa29fa0afae8f9c5f9adf992f977f9;
    inBuf[2528] = 256'h62f94af92ef918f9fcf8ddf8c1f8a0f880f864f845f828f811f8f9f7e5f7d7f7;
    inBuf[2529] = 256'hc8f7c0f7bcf7b7f7b8f7bdf7bff7c9f7d7f7e4f7f9f711f828f848f868f886f8;
    inBuf[2530] = 256'haff8d8f8fbf828f957f980f9b1f9e3f911fa47fa7cfaaefae9fa23fb57fb95fb;
    inBuf[2531] = 256'hd2fb08fc47fc85fcbdfcfffc42fd80fdc6fd0bfe4cfe96feddfe1eff65ffa9ff;
    inBuf[2532] = 256'he4ff22005d009000c500f4001d0148016f019001b601d601f2010f0229023e02;
    inBuf[2533] = 256'h54026802780289029602a302b102bc02c702d402dd02e702f002f502fa02fd02;
    inBuf[2534] = 256'hfa02f902f602ed02e602de02d202c802bf02b202a8029d028f02830276026402;
    inBuf[2535] = 256'h550248023702270219020c020002f601ef01e901e301df01dd01d701d201ca01;
    inBuf[2536] = 256'hbf01b301a4018f017b01640147012c010e01ec00cd00ab00840061003a000f00;
    inBuf[2537] = 256'he9ffbdff8bff61ff31fffafecbfe97fe5dfe2bfef4fdb6fd81fd45fd02fdc9fc;
    inBuf[2538] = 256'h89fc41fc02fcbefb72fb30fbe9fa9bfa57fa0efac2f980f938f9eff8b1f86ef8;
    inBuf[2539] = 256'h2bf8f2f7b7f77cf74bf719f7ebf6c4f69cf67af660f643f62df61ef60df602f6;
    inBuf[2540] = 256'hfcf5f4f5f2f5f5f5f4f5fcf508f60ff622f638f64bf66af68df6aef6dcf60df7;
    inBuf[2541] = 256'h3cf77bf7b9f7f5f741f88cf8d2f827f97cf9cbf927fa80fad5fa36fb94fbebfb;
    inBuf[2542] = 256'h51fcb2fc0dfd74fdd7fd33fe9cfefffe5dffc6ff27008400ec004b01a5010a02;
    inBuf[2543] = 256'h6602be0220037b03d20331048704dd043a058c05de0534067e06c80615075507;
    inBuf[2544] = 256'h9507d6070b08410876089f08cc08f80818093c09600979099609b209c309db09;
    inBuf[2545] = 256'hf009fa090d0a1c0a210a2e0a380a390a420a460a420a430a3d0a300a290a180a;
    inBuf[2546] = 256'h000aed09d209b209960973094c092a090009d508ae087e084d082008e807af07;
    inBuf[2547] = 256'h78073607f506b6066c062506e10591054705fe04aa045c040f04b4035e030703;
    inBuf[2548] = 256'ha3024402e20174010d01a3002e00c3ff57ffe1fe76fe0afe96fd2cfdc1fc4ffc;
    inBuf[2549] = 256'he8fb7efb0efbabfa45fadaf97bf91af9b6f85ef802f8a5f753f7fcf6a5f659f6;
    inBuf[2550] = 256'h07f6b7f573f529f5e4f4abf46ef438f40df4dff3b9f39ef37ef367f35bf349f3;
    inBuf[2551] = 256'h41f341f33df345f353f35df376f394f3adf3d6f303f42af461f49bf4d0f413f5;
    inBuf[2552] = 256'h57f597f5e6f534f67ef6d8f631f786f7ebf74df8adf81df989f9f4f970fae6fa;
    inBuf[2553] = 256'h5cfbe4fb65fce6fc78fd02fe8bfe23ffb0ff3c00d5005f01ea01810208039103;
    inBuf[2554] = 256'h2604ac043505cb055306de067407fa078508170998091c0aa60a1e0b980b170c;
    inBuf[2555] = 256'h840cf50c6a0dcd0d360ea10efa0e590fb70f04105410a210de101d1157118011;
    inBuf[2556] = 256'had11d311e911051217121b122512241216120c12f711d611ba1191115e113311;
    inBuf[2557] = 256'hf810b7107e103610e80fa20f4b0fef0e980e300ec30d5b0ddf0c610ce80b5d0b;
    inBuf[2558] = 256'hd20a4e0abb092a09a1080a087807ed065406c1053405980401047103d2023902;
    inBuf[2559] = 256'ha60107016f00ddff40ffaefe20fe8afdfefc77fce7fb63fbe1fa59fadcf95ff9;
    inBuf[2560] = 256'hdcf865f8ebf770f700f78ff61df6b7f550f5eaf492f437f4e0f398f34bf304f3;
    inBuf[2561] = 256'hccf28ef256f22bf2faf1cff1aef186f165f14ef12ef117f109f1f4f0e9f0e9f0;
    inBuf[2562] = 256'he3f0e7f0f6f000f117f135f14ff177f1a4f1ccf103f23ef275f2b9f202f348f3;
    inBuf[2563] = 256'h9cf3f1f346f4aaf40df570f5e3f553f6c4f644f7c1f740f8cef856f9e1f97bfa;
    inBuf[2564] = 256'h0dfba2fb47fce0fc7dfd29fec9fe6dff1f00c4006f012902d40287034804fa04;
    inBuf[2565] = 256'hb20577062a07e207a3085109020ab80a590bfe0ba70c3a0dd20d6e0ef60e830f;
    inBuf[2566] = 256'h131091101311961106127a12ea124613a613fd1340148614c214eb1416153715;
    inBuf[2567] = 256'h47155b1562155b155a1549152b151215e914b41483144014f213a9134c13e612;
    inBuf[2568] = 256'h87121212961123119a100d10890ff20e580ec90d270d860cf00b460ba00a060a;
    inBuf[2569] = 256'h5909af0810085f07b2060f065905a90403044c039c02f80143019900faff4fff;
    inBuf[2570] = 256'haffe1afe7bfde9fc60fccdfb49fbcbfa43fac9f954f9d6f866f8f9f786f71ff7;
    inBuf[2571] = 256'hbbf653f6f9f5a0f544f5f9f4adf45ff421f4e1f3a1f36ef337f300f3d4f2a3f2;
    inBuf[2572] = 256'h72f24ef221f2f6f1daf1b5f194f182f16af158f154f14bf14af155f159f165f1;
    inBuf[2573] = 256'h7bf189f19ef1bbf1d0f1ebf10df228f24df277f29cf2ccf203f335f375f3bbf3;
    inBuf[2574] = 256'hfdf34df4a0f4f1f44ff5aef50bf676f6def645f7baf72cf89ef81df997f913fa;
    inBuf[2575] = 256'h9efa21fba6fb3afcc5fc52fdeefd80fe14ffb6ff4b00e30087011d02b5025803;
    inBuf[2576] = 256'hec0381042005af053f06d8066207ef07830807098f091c0a990a190b9d0b0f0c;
    inBuf[2577] = 256'h830cf60c580db90d170e640eb20efa0e310f6a0f9d0fc20fe90f0a101e103710;
    inBuf[2578] = 256'h47104b105410511043103a1023100110e30fb60f7f0f4c0f090fc00e7c0e290e;
    inBuf[2579] = 256'hd00d7f0d200dbe0c620cf70b8b0b270bb20a3b0acb094a09c9084e08c3073807;
    inBuf[2580] = 256'hb506230695050f057c04ee036a03db025302d2014601c2004400baff3affbefe;
    inBuf[2581] = 256'h36feb7fd3cfdb7fc3bfcc2fb41fbcbfa57fadcf96ef901f98ef828f8c3f75af7;
    inBuf[2582] = 256'hfff6a2f643f6f1f59bf543f5f9f4aaf458f414f4caf37ef341f3fcf2b8f283f2;
    inBuf[2583] = 256'h49f211f2e7f1b7f18bf16ff14cf12bf118f1fcf0e6f0daf0c4f0b4f0aef09ef0;
    inBuf[2584] = 256'h96f099f092f094f0a3f0abf0bef0dcf0f2f016f142f166f198f1d2f101f23bf2;
    inBuf[2585] = 256'h7bf2b2f2f5f23af377f3c1f30df451f4a5f4faf447f5a7f508f663f6cef639f7;
    inBuf[2586] = 256'h9df711f882f8edf867f9daf946fabffa33fb9efb17fc8afcf7fc71fde5fd54fe;
    inBuf[2587] = 256'hcffe43ffb4ff3100a50014018d01fc016702d8024003a3030b046a04c6042605;
    inBuf[2588] = 256'h7b05cf0527067606c30614075d07a507ef0730087208b508ef08280960098f09;
    inBuf[2589] = 256'hbd09e709080a290a460a5a0a6d0a7a0a810a890a8d0a8c0a8c0a870a7e0a780a;
    inBuf[2590] = 256'h6b0a5b0a4c0a330a170afc09d409aa0980094a091209db08990857081608cc07;
    inBuf[2591] = 256'h83073d07ed069f065206fa05a7055105f00492043304c8036203f80283021602;
    inBuf[2592] = 256'ha6012d01bc004900ceff5effeafe6ffefffd8cfd12fda4fc31fcb5fb46fbd5fa;
    inBuf[2593] = 256'h5afaebf97af903f998f828f8b6f752f7e9f67ef623f6c5f565f512f5bef46bf4;
    inBuf[2594] = 256'h24f4d8f390f354f312f3d3f2a1f269f234f20cf2ddf1b4f198f176f15cf14ef1;
    inBuf[2595] = 256'h39f12ef12ff129f12cf13af140f151f16bf17af194f1b5f1ccf1eff119f238f2;
    inBuf[2596] = 256'h62f294f2bcf2f0f22cf35ef39cf3e1f31df466f4b3f4f5f444f597f5dcf52ef6;
    inBuf[2597] = 256'h82f6c9f61bf770f7b9f70cf862f8aef805f95df9aff90afa66fabbfa19fb76fb;
    inBuf[2598] = 256'hcefb2dfc88fcdefc3bfd93fde8fd43fe98feebfe46ff9cfff1ff4c00a300fc00;
    inBuf[2599] = 256'h5a01b3010d026c02c4021e037c03cf0324047f04d00421057405c0050e065d06;
    inBuf[2600] = 256'ha406ee0639077d07c307080847088a08ca08040940097909aa09dd090d0a340a;
    inBuf[2601] = 256'h5e0a820a9e0aba0acf0ade0aef0af90afd0a030b020bfc0af60ae90adb0acc0a;
    inBuf[2602] = 256'hb20a960a7a0a500a250af909be0983094809fe08b6086f081a08c80779071d07;
    inBuf[2603] = 256'hc60670060e06b3055805ef048b042904b8034c03e2026d02fd018d0111019d00;
    inBuf[2604] = 256'h2d00b5ff43ffd5fe5efef1fd88fd19fdb2fc4efce5fb86fb2dfbcdfa74fa21fa;
    inBuf[2605] = 256'hc9f979f92df9e1f89cf859f818f8e0f7a9f775f74af724f701f7e4f6c8f6b2f6;
    inBuf[2606] = 256'ha4f695f68af686f680f67ff686f68af693f6a3f6b1f6c7f6e3f6fcf61df745f7;
    inBuf[2607] = 256'h6af797f7c8f7f7f72df867f89df8d9f817f951f991f9d1f90cfa4efa8ffacafa;
    inBuf[2608] = 256'h0dfb50fb8efbd3fb18fc5bfca5fcedfc36fd86fdd3fd1efe6ffebefe0dff5eff;
    inBuf[2609] = 256'habfff9ff48009100de002f017801c60117026002b00204034f03a103f5033e04;
    inBuf[2610] = 256'h8d04df0425057305c00501064c069906d7061d076607a507ed0736087408ba08;
    inBuf[2611] = 256'h00093c098109c509fe093d0a7c0ab00aea0a1f0b4a0b7b0ba70bc70bef0b120c;
    inBuf[2612] = 256'h2b0c490c610c700c870c970ca00cb00cb90cba0cc20cc10cb90cb60ca80c960c;
    inBuf[2613] = 256'h8a0c6e0c4c0c300c080cdc0bb30b7b0b430b120bd20a900a540a090abf097c09;
    inBuf[2614] = 256'h2809d40885082708c80770070a07a5064506d9056f050c059d043104ce036303;
    inBuf[2615] = 256'hfc029a023102cc016c010601a2004600e5ff83ff27ffc8fe6afe10feb7fd63fd;
    inBuf[2616] = 256'h12fdbffc73fc2dfce8fba9fb71fb3dfb0cfbe1fabafa99fa7dfa65fa50fa3efa;
    inBuf[2617] = 256'h30fa25fa1ffa1efa1efa22fa2bfa36fa45fa5bfa70fa89faabfaccfaedfa19fb;
    inBuf[2618] = 256'h43fb6bfb9cfbcdfbfcfb33fc67fc9cfcd8fc11fd4bfd8efdccfd0cfe55fe96fe;
    inBuf[2619] = 256'hd9fe27ff6dffb2ff000047008c00d8001b015c01a101df011b025b029302c902;
    inBuf[2620] = 256'h020334036903a103d10306043f046d04a104da0408053a056f059805c705f705;
    inBuf[2621] = 256'h1a0642066c068b06ab06cd06e806070725073c07590775078907a207ba07cc07;
    inBuf[2622] = 256'he307f6070208140822082a0838084308470852085b085e0867086c086d087408;
    inBuf[2623] = 256'h7608720874087108680865085a0849083d0829081008fb07de07bb079d077607;
    inBuf[2624] = 256'h4d072807fa06cb06a20670063e061106db05a50573053805fc04c2047e043904;
    inBuf[2625] = 256'hf403a60359030c03b4025f020c02b1015601fe00a0004500e9ff89ff2dffd0fe;
    inBuf[2626] = 256'h6ffe14feb6fd54fdf8fc9cfc3efce7fb8dfb36fbe6fa93fa40faf9f9b3f96bf9;
    inBuf[2627] = 256'h2cf9eef8b2f87df847f815f8eaf7bef796f773f750f732f71af701f7eff6e4f6;
    inBuf[2628] = 256'hd6f6d3f6d8f6ddf6ecf602f717f736f75cf782f7aef7e0f711f847f881f8bbf8;
    inBuf[2629] = 256'hfaf838f978f9c0f907fa4cfa9afae6fa30fb83fbd3fb22fc7afccefc1ffd76fd;
    inBuf[2630] = 256'hcbfd1efe76fec9fe1bff73ffc1ff10006500b100fa004b019401d90127026a02;
    inBuf[2631] = 256'ha802ed022b036603a403d90309043a0462048704ae04cc04e504000514052405;
    inBuf[2632] = 256'h36054805570562056a0576057f0584058c05920592058f058b0584057b056d05;
    inBuf[2633] = 256'h5e0550053c0522050a05ef04d304b704970478045b0438041504f403cf03ab03;
    inBuf[2634] = 256'h8903660341031b03f202cc02a7027e0256022e020002d701b101830155012a01;
    inBuf[2635] = 256'hfd00d200a4006f003f000e00d5ffa1ff6bff2ffff5febafe7afe3dfefdfdbafd;
    inBuf[2636] = 256'h7dfd3efdfbfcbffc7efc3cfc02fcc4fb82fb49fb0cfbcafa8ffa4efa0cfad0f9;
    inBuf[2637] = 256'h8cf945f909f9c7f883f847f806f8c2f788f74cf713f7e0f6a7f674f64bf61cf6;
    inBuf[2638] = 256'hf0f5cdf5a7f586f56df54ff537f526f50ff502f5fdf4f2f4eff4f2f4f0f4f8f4;
    inBuf[2639] = 256'h08f512f526f540f554f56ff592f5b2f5daf506f62ef660f696f6c7f603f744f7;
    inBuf[2640] = 256'h81f7c8f711f859f8abf8fdf84bf9a4f9fef952fab0fa0cfb62fbc3fb1efc73fc;
    inBuf[2641] = 256'hd4fc30fd82fdddfd36fe86fedffe32ff7dffd3ff24006b00ba00050147019101;
    inBuf[2642] = 256'hd701130253028f02c602ff0231035b038703af03d003f0030c04230439044904;
    inBuf[2643] = 256'h53045d04620463046404600456044704370424040e04f703db03bb039e038003;
    inBuf[2644] = 256'h5b0337031003e702c1029d02720247021c02ed01c1019301620135010701d100;
    inBuf[2645] = 256'h9e006e0038000500d2ff9fff6fff3eff0bffddfeaffe7efe54fe2afefffdd8fd;
    inBuf[2646] = 256'hb3fd8cfd6cfd4afd23fd04fde7fcc6fca9fc8dfc6efc52fc36fc17fcfefbe4fb;
    inBuf[2647] = 256'hc9fbb3fb9afb7efb68fb4ffb37fb24fb0cfbf4fae3facafab2faa2fa8dfa76fa;
    inBuf[2648] = 256'h69fa54fa3ffa35fa23fa0efa06fafaf9e7f9dbf9cdf9bff9b6f9a8f999f991f9;
    inBuf[2649] = 256'h83f976f96ef961f955f950f947f940f93df939f939f93df93ef944f94ff956f9;
    inBuf[2650] = 256'h63f975f983f995f9abf9bef9d7f9f3f90afa27fa49fa64fa85faadfad0faf7fa;
    inBuf[2651] = 256'h23fb4dfb7afbaafbdafb0cfc41fc75fcadfce6fc1bfd57fd94fdcffd0efe4cfe;
    inBuf[2652] = 256'h87fec9fe0cff49ff8bffcbff070047008900c800090145017e01bb01f5012a02;
    inBuf[2653] = 256'h62029502c402f50223034c0374039903bd03e103030422043f04590473048a04;
    inBuf[2654] = 256'h9c04b004c004c904d304dc04e004e104de04d804d304c804ba04af04a1048c04;
    inBuf[2655] = 256'h79046504500439041e040504ef03d203b4039703770359033e031b03f902dc02;
    inBuf[2656] = 256'hba0298027a02570237021e020002e001c601aa018f0179015e01460134011e01;
    inBuf[2657] = 256'h0501f400e200cc00bc00ae009f00920086007b0073006c006600630060006000;
    inBuf[2658] = 256'h62006400660069006c0073007c00820088008e0093009c00a800b000b700c000;
    inBuf[2659] = 256'hc900d400e000eb00f800060112011e012901340140014c0154015e0168016f01;
    inBuf[2660] = 256'h74017c01830188018d019101960199019c019e01a001a101a201a501a501a101;
    inBuf[2661] = 256'h9e019a01960192018d0185017f0176016d0167015e01550151014b0143013c01;
    inBuf[2662] = 256'h36012f012b01260122011f011901130112010f010a0109010801040106010a01;
    inBuf[2663] = 256'h0a010a010e0116011e0124012b01350140014a015801670173017f018d019b01;
    inBuf[2664] = 256'hab01bd01cc01dc01ee01ff0115022a023a0250026a0280029802b002c402dc02;
    inBuf[2665] = 256'hf8020f03230338034c036303780388039c03b003c003d303e403f10304041604;
    inBuf[2666] = 256'h2204340441044a045a0467046c047804820486048f04960496049b04a104a004;
    inBuf[2667] = 256'ha304a604a604a904a904a504a704a804a304a704a7049f049e049c0496049704;
    inBuf[2668] = 256'h94048c048e048e0488048c048d0488048f04970498049f04a404a704b904c404;
    inBuf[2669] = 256'hc404d304e304e804f60401050705180525052c053e054c055405660576058005;
    inBuf[2670] = 256'h9305a505b005c005cd05d905eb05f405fa050a06130617061f0621061d062106;
    inBuf[2671] = 256'h21061d061d0613060306fc05ee05da05cb05b7059b058105630542052005f904;
    inBuf[2672] = 256'hd204aa04780448041d04e703b00380034a030f03d8029b025f022502e401a401;
    inBuf[2673] = 256'h67012201df009c0053000e00cdff84ff3ffffdfeb7fe76fe36fef2fdb8fd80fd;
    inBuf[2674] = 256'h42fd0efddefca8fc78fc4efc22fcfcfbdafbb6fb9afb80fb64fb51fb44fb33fb;
    inBuf[2675] = 256'h26fb20fb1cfb1cfb20fb27fb31fb3ffb51fb64fb79fb93fbaffbcefbedfb0ffc;
    inBuf[2676] = 256'h38fc62fc88fcb6fceafc19fd4dfd89fdbefdf6fd39fe76feb1fef2fe2dff6aff;
    inBuf[2677] = 256'hadffe8ff240064009d00d700150146017801b501ec011c0251028202b302e602;
    inBuf[2678] = 256'h12033f036f039703bd03eb0310043104560473048b04aa04c704dd04f1040505;
    inBuf[2679] = 256'h1b052c053805470553055e056a05730577058105860585058805880584058605;
    inBuf[2680] = 256'h85057f057d05770571056f056a056505630559054f054e0547053c0534052605;
    inBuf[2681] = 256'h19050d05f704e304d304ba04a1048b046d044f0435041204f203d403ad038903;
    inBuf[2682] = 256'h66033c031603ed02bb028c025d022702f201bb017c0140010101bc0079003200;
    inBuf[2683] = 256'he8ffa0ff50fffefeb5fe63fe0bfebcfd64fd09fdb7fc5ffc01fcaffb56fbf7fa;
    inBuf[2684] = 256'h9efa43fae9f99af943f9ebf8a0f850f8fef7b9f770f726f7e8f6a7f664f62df6;
    inBuf[2685] = 256'hf6f5c0f591f560f534f512f5edf4cef4bbf4a3f491f48cf488f489f493f49df4;
    inBuf[2686] = 256'hadf4c9f4e6f409f531f55af58ff5c6f5faf53af67df6bef60bf75af7a5f7fcf7;
    inBuf[2687] = 256'h52f8a6f809f96bf9c6f92efa95faf8fa64fbcefb36fca8fc14fd7afdeafd56fe;
    inBuf[2688] = 256'hbcfe2aff92fff5ff5f00c10020018601e20139029902ed023a038f03da031904;
    inBuf[2689] = 256'h5e049b04cf0409053d0564058b05af05cc05e805ff050f0620062c0632063706;
    inBuf[2690] = 256'h3a0636062d06240616060406f105da05bb059d057f0556052d050605d504a404;
    inBuf[2691] = 256'h750440040a04d6039c0361032703e802ad0274023202f201b60173013401f600;
    inBuf[2692] = 256'hb0006f003200edffaeff70ff2bffedfeb0fe6cfe2efef1fdadfd70fd2ffde9fc;
    inBuf[2693] = 256'habfc6cfc27fce8fba4fb60fb25fbe3fa9ffa62fa21fae1f9a8f966f926f9f1f8;
    inBuf[2694] = 256'hb2f873f83ff803f8caf796f756f71df7edf6aff675f648f610f6d9f5abf574f5;
    inBuf[2695] = 256'h42f51bf5e9f4bcf49af46ff44bf430f40ef4f0f3dbf3c2f3b0f3a4f393f38cf3;
    inBuf[2696] = 256'h8bf384f387f391f399f3a9f3baf3caf3e9f30bf426f44ff47cf4a3f4d7f410f5;
    inBuf[2697] = 256'h45f586f5c9f506f652f6a2f6ecf642f79bf7f0f753f8b5f813f97ff9e9f950fa;
    inBuf[2698] = 256'hc3fa34fba1fb17fc8cfcfcfc75fde8fd58fecffe3fffabff1f008b00f4006301;
    inBuf[2699] = 256'hc9012a029402f5024d03ab0302045104a304f00435057b05ba05f00526065a06;
    inBuf[2700] = 256'h8506ac06ce06e706fd0612071f072507290725071a070e07fa06e106c706a506;
    inBuf[2701] = 256'h7c0652062406f005bb057e053d05fd04b80470042a04dd038a033b03ea029302;
    inBuf[2702] = 256'h4002ea018f013801de0081002900ceff6eff16ffb9fe5afe04feaafd4efdfafc;
    inBuf[2703] = 256'ha3fc4afcfdfbaffb5cfb13fbc9fa81fa42fafef9baf982f945f90af9dbf8a7f8;
    inBuf[2704] = 256'h73f849f81af8eff7cff7a8f785f76df74bf72ef71ef706f7f1f6e5f6d2f6c3f6;
    inBuf[2705] = 256'hbdf6b0f6a9f6aaf6a1f6a1f6a9f6a5f6a8f6b4f6b6f6bff6d3f6dff6edf600f7;
    inBuf[2706] = 256'h0ff725f73cf74ef76af785f799f7b9f7d9f7eff711f835f851f876f89ef8bff8;
    inBuf[2707] = 256'heaf815f93cf96cf99df9caf9fff933fa63fa9dfad6fa0bfb4afb86fbc0fb02fc;
    inBuf[2708] = 256'h3efc7bfcc3fc05fd44fd8cfdccfd0dfe5bfea1fee2fe30ff78ffbdff0c005400;
    inBuf[2709] = 256'h9900e6002c016f01bb01010244028c02d002110355039403d10310044b048604;
    inBuf[2710] = 256'hc204f60429055c058a05b805e00504062b064e06670682069c06af06c106d106;
    inBuf[2711] = 256'hdc06e706eb06ec06ed06ea06e506df06d106c106b2069c0683066a064b062b06;
    inBuf[2712] = 256'h0c06e405ba059305650538050d05db04a70475043f040904d5039c0366033303;
    inBuf[2713] = 256'hf902c0028a024f021502e201ac01740141010c01d800a700750046001a00eaff;
    inBuf[2714] = 256'hbfff9cff73ff4bff2aff08ffe9fed2feb6fe9bfe89fe74fe5ffe55fe49fe3dfe;
    inBuf[2715] = 256'h3afe36fe31fe36fe39fe3afe44fe53fe5dfe6dfe7ffe90fea4febbfed3feeefe;
    inBuf[2716] = 256'h09ff23ff45ff65ff82ffa5ffcbffedff14003e0062008900b600df0007013201;
    inBuf[2717] = 256'h5c018a01b701dc010502320259028002ab02d102f7021e03410365038903a903;
    inBuf[2718] = 256'hc903e70301042204400455046e0488049a04b004c504d404e804fb0404051205;
    inBuf[2719] = 256'h1f05260532053d05410548054b054b05500552054f05530553054b054a054805;
         
    encBuf[0] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[1] = 256'h0008000800080008000800080008000800080008000800080008000800080008;    
    encBuf[2] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[3] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[4] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[5] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[6] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[7] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[8] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[9] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[10] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[11] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[12] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[13] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[14] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[15] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[16] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[17] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[18] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[19] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[20] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[21] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[22] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[23] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[24] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[25] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[26] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[27] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[28] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[29] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[30] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[31] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[32] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[33] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[34] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[35] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[36] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[37] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[38] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[39] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[40] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[41] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[42] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[43] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[44] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[45] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[46] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[47] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[48] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[49] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[50] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[51] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[52] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[53] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[54] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[55] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[56] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[57] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[58] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[59] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[60] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[61] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[62] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[63] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[64] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[65] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[66] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[67] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[68] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[69] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[70] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[71] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[72] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[73] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[74] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[75] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[76] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[77] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[78] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[79] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[80] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[81] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[82] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[83] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[84] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[85] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[86] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[87] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[88] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[89] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[90] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[91] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[92] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[93] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[94] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[95] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[96] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[97] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[98] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[99] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[100] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[101] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[102] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[103] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[104] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[105] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[106] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[107] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[108] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[109] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[110] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[111] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[112] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[113] = 256'h0008000800080008000800080008000800080009010800080008000800080008;
    encBuf[114] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[115] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[116] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[117] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[118] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[119] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[120] = 256'h0008000800080008000800080008000800080008080000080008000800080008;
    encBuf[121] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[122] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[123] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[124] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[125] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[126] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[127] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[128] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[129] = 256'h0008000800080000080800080009010800080008080000080008080801080008;
    encBuf[130] = 256'h0008000800090108000800080008000901080008000800090108080801080008;
    encBuf[131] = 256'h0009010800080008000800080008000800080000080800000900000800080008;
    encBuf[132] = 256'h0008000800080008000808080100090000080800000009000008080000080008;
    encBuf[133] = 256'h0008000800080008080000080008000800080800000800000900000800080008;
    encBuf[134] = 256'h0008000800080008000800080008000800080008000808080100080900000008;
    encBuf[135] = 256'h0008000901080008000800090100080800080008000800080008000800080000;
    encBuf[136] = 256'h0908010808000008000800080008000800090100080800080009010008080801;
    encBuf[137] = 256'h0808000800080000090000080008000800080008000800080008000800000900;
    encBuf[138] = 256'h0008000800080008000800080008080000080008000900000008000800080008;
    encBuf[139] = 256'h0008000808000008000800080000090000080008000800000908010808080108;
    encBuf[140] = 256'h0008000800090100090000080008000800080008000800080008000800080008;
    encBuf[141] = 256'h0008000800090108000800080008000800080008000800080008000800080008;
    encBuf[142] = 256'h0008000800080008080000080008000800080008000800080008000008080008;
    encBuf[143] = 256'h0008000800000900000009080108000800080008000808080108000800080008;
    encBuf[144] = 256'h0008000008080008000800080008000800080008000901080009010800090108;
    encBuf[145] = 256'h0008000800080009010008080800000800080000090000080800000009010908;
    encBuf[146] = 256'h0108000800080008080000080008000800090000000800080008000800080808;
    encBuf[147] = 256'h0100090000080008080801000900000900000008000800080008000800080008;
    encBuf[148] = 256'h0008000901080008000800080008000009000008000800080008000800080008;
    encBuf[149] = 256'h0800000800000808000800080008000009000008000800080008000800080008;
    encBuf[150] = 256'h0008000800080808010009080008010800080008000800080008000800080008;
    encBuf[151] = 256'h0008000800080008000800080008000800080009000000080800000800080008;
    encBuf[152] = 256'h0008000800080008000800080008000800090100080800080008000800080000;
    encBuf[153] = 256'h0808000800080008000800080008000800080008000800080008000800080008;
    encBuf[154] = 256'h0008000008080800000800080008000800080008000800080008000800080008;
    encBuf[155] = 256'h0008000800080008000009000008000800080008000800080008000900000009;
    encBuf[156] = 256'h0000000800080008000901080008000008080008000800080008000009000009;
    encBuf[157] = 256'h0000000800080008000800080008000800080008000800090108080801000908;
    encBuf[158] = 256'h0108000800080008000800080000090800000008000800090000000800000900;
    encBuf[159] = 256'h0008000800080008000800080008000901080008000800080008000800080008;
    encBuf[160] = 256'h0000090000080008000800080008000800080000090000080008000009000009;
    encBuf[161] = 256'h0108000800080008080801090100090000080808000800000008000009080100;
    encBuf[162] = 256'h0908010800080008000009080108000800080008000900000008000008080009;
    encBuf[163] = 256'h0108080000080008000901000900000008080800000009000009000000080008;
    encBuf[164] = 256'h0008000800080008000901000908010800080008000800080000090000080008;
    encBuf[165] = 256'h0008000800080008000800090000000800080808010800090000000800080008;
    encBuf[166] = 256'h00080000090800080908030603090f0b02010c0a03030103020c0e0801010200;
    encBuf[167] = 256'h0809000001040401090e0c0205080f09000109020400090001080b0908000109;
    encBuf[168] = 256'h0b090101090e0d0902000c0207030801020d0e0802010a0a0901010200000009;
    encBuf[169] = 256'h0901040403090f0d01020103040a0d01030b0f0a02020100080900000808090b;
    encBuf[170] = 256'h0c0808000706090802090e00040a0b0707070108000808080000080000080808;
    encBuf[171] = 256'h09090908090801000900000a0c0a0a0a0005030008090a010202080102000407;
    encBuf[172] = 256'h0603030208090800080305030402000801000a0b090b0c0004010800090d0b0b;
    encBuf[173] = 256'h0c0d09090a0900080b0b0b0f0d090908000100000001000001080a0802020607;
    encBuf[174] = 256'h0302030401000108080002040404020108080b0c0908080000090b0c0c0b0b0a;
    encBuf[175] = 256'h0b0c0b0b0c0b0b0c0e0b0c0a0801010108090b0d090801020304020101010203;
    encBuf[176] = 256'h030203020304030200000800040702080b0f0f0c0b0a080808080a0c0c0c0b0b;
    encBuf[177] = 256'h0a09080809080909090a0a0c0c0a090104040201000a09010406030403010000;
    encBuf[178] = 256'h020404030201000909090a0c0d0d0c0b0a0a090a0c0d0c0b0c0a090909090b0a;
    encBuf[179] = 256'h0c0b0a0b0a0c0a0a0a0908080a0c0c0b0a000206040304020202020305030403;
    encBuf[180] = 256'h0301000809090908090a0c0d0b0c0b0a0a0a0b0b0b0b0c0c0d0d0c0b0c090a08;
    encBuf[181] = 256'h090a0c0b0b0b0a0a0a0b0c0b0908020404030201000808000405040503020201;
    encBuf[182] = 256'h080a0c0b0a09010202080a0f0b0b0c09080809090b0d0d0b0b0a080001080a0f;
    encBuf[183] = 256'h0c0c0b0a090102050302080a0c0c0a0902050403030108090b0a080103050303;
    encBuf[184] = 256'h0301080a0d0b0b0b0a0009090d0e0c0a0b090008080b0d0d0b0a0a0800010101;
    encBuf[185] = 256'h01080c0d0a0b0902030603030101080001010305040404020203000101020404;
    encBuf[186] = 256'h020100090b0b0b09080a0a0a0e0b0b0e0c0b0d0b09080801080a0c0c0b0a0909;
    encBuf[187] = 256'h000a0a090b080201050402030503040401030303050502030301000008090008;
    encBuf[188] = 256'h00030405030201080b0a08090103090d0d0e0b0a0a0b0a0d0b0b0a0900080000;
    encBuf[189] = 256'h0a08040406030302030304040302030102040403050201000800010100010909;
    encBuf[190] = 256'h010107040201000b0b0a0a0a090f0b0c0c090909090a0c0b0a09000203050403;
    encBuf[191] = 256'h0404030402020304030503020100000103050403030201080808090809090908;
    encBuf[192] = 256'h000101090f0c0e0c0a0909000808080b0c0b0a0a080808010800000104060405;
    encBuf[193] = 256'h04030403030303030502020302020204040304030200000a090a0a0a0a0a0909;
    encBuf[194] = 256'h080100080d0f0d0c0b0b0b080003040302080a0c0e0b0a0a0801040504030302;
    encBuf[195] = 256'h0100000001040405030402000008080800010202010009090801020503020108;
    encBuf[196] = 256'h0b0c0c0b0900020302090f0d0c0a090003060302020000090a08010207050404;
    encBuf[197] = 256'h0201000a0b0c0a08010303040200080a0b0c0a0b09080003040203040101080b;
    encBuf[198] = 256'h0c0b0d0901010404010201000202030503030504040503030301000008010403;
    encBuf[199] = 256'h03040108090b0d0b0c0a08000102010a0d0e0c0b0a0909090900080900090b0b;
    encBuf[200] = 256'h0f0b0a0908000009080808060503040108080a0a010406050303040200000a0a;
    encBuf[201] = 256'h09090104030303000908090900090d0a0c0a000000000b0f0a0c0b0a0b0b0b0d;
    encBuf[202] = 256'h0a09000002090c0c0d0c090a0900080a08090a090a0c090b0b01020204000a08;
    encBuf[203] = 256'h0a0903090e0c0d0c08010406030201090b0b0c09010203060200010909080908;
    encBuf[204] = 256'h010102040100030101050200010b0f0d0c0d0a0a0900000101090e0c0e0b0a09;
    encBuf[205] = 256'h0901010101080b0c0c0c0a090901010001090b0c0c0b08080002010101020205;
    encBuf[206] = 256'h0304040202020202030303040303040201090c0c0b0b0a08080800090c0b0d0c;
    encBuf[207] = 256'h0b0c0b0b0c0b0d0c0a0b0a09080a0c0d0d0c0a0a0900000100090b0d0b0a0a09;
    encBuf[208] = 256'h080102030201090c0d0b0901030503010a0c0c0a09000103040100090b0c0b09;
    encBuf[209] = 256'h00060505030202000a0a0a090307030302000a0c0b09000205020208090a0a09;
    encBuf[210] = 256'h09080a0c0b0d0d0b0b0e0b0b0b0a080000090f0d0c0b0a090003020100090b0c;
    encBuf[211] = 256'h0b0a090102060403030200080909010504040402020201030203040201000000;
    encBuf[212] = 256'h0101010100090a0b0f0d0c0c0a090800030101090e0c0b0c090900020201080a;
    encBuf[213] = 256'h0f0b0c0a09080103030201000a0a0a0a01030505030201010908090900000800;
    encBuf[214] = 256'h080d0c0b0d09080801010a0b0c0e09000307050202010809090a010205040302;
    encBuf[215] = 256'h01000a0b0a0803070503030200080a090a0908000800090c0c0e0c0b0b090801;
    encBuf[216] = 256'h00000b0f0c0c0a09080001080a0b0c0c09090801010304040303020008000307;
    encBuf[217] = 256'h0504020301000000000100010101030503030308090a0c0a0102050303020008;
    encBuf[218] = 256'h0a0d0e0c0c0c0a0909000008080a0b0b0b0b0b0900030605030402010008090a;
    encBuf[219] = 256'h0a09090002060304040108090c0b0a09020504040201080a0b0d0b0b09000305;
    encBuf[220] = 256'h040101000a0b0a0b08020506040302020008090a080102050303020201000202;
    encBuf[221] = 256'h04020201090a0c0a0a000101000d0f0f0d0b0c0a090900010201080a0c0c0b0b;
    encBuf[222] = 256'h0901030504020000090a09080204050402020208000002040604030201000808;
    encBuf[223] = 256'h010204040202080b0b0d0a0a09080008090a0c0d0b0c0b0908020403010a0d0d;
    encBuf[224] = 256'h0b0b080003030200090b0d09080307040303030000090800030505030301080a;
    encBuf[225] = 256'h0c0b0a0a080202040100090c0b0c090900000800090800020503030101090a0c;
    encBuf[226] = 256'h0d0b0900070604040200000a0a09010305050202010809090a0a090a09000801;
    encBuf[227] = 256'h010a0c0f0c0c0a0a09080808080a0a0a0b0a0a09080801030505040403030302;
    encBuf[228] = 256'h02020101020102030405060303030100090a090306050403020208090c0e0b0c;
    encBuf[229] = 256'h0b0a090100000a0d0e0c0a0a090000000001000202020008090a080103060200;
    encBuf[230] = 256'h080a00020504030008080803070603030200000a09090800000100090d0d0d0c;
    encBuf[231] = 256'h0b0c0a0a080800090a0c0c0a0a09080101010201000101010304040304020302;
    encBuf[232] = 256'h02010305060305030202010809090908010201090f0d0b0c0a0909090a0b0d0b;
    encBuf[233] = 256'h0c0a0a0b0a0a0a0b090909080909080003070404040203030204020303040102;
    encBuf[234] = 256'h030103040304030101090b0e0b0d0a0a0a0a090a0c0d0d0b0d0b0a0a090a090a;
    encBuf[235] = 256'h0a090a08080809090b0a01050604030302010303030503020202020505040303;
    encBuf[236] = 256'h020100000001020101080a0b0e0b0d0c0c0d0b0c0b0b0a0b0a0b0b0c0b0a0b0a;
    encBuf[237] = 256'h0909000204060304030101000908090000020304040402030200000809000204;
    encBuf[238] = 256'h07050304010100090b0b0d0c0b0b0c0a0909080809090b0a0901040603020100;
    encBuf[239] = 256'h080a090a09080a000909090b0f0e0c0c0c0a0a09000203040202010100080809;
    encBuf[240] = 256'h0a0a090802060603050302030101000000030305030401020808090b0f0b0d0b;
    encBuf[241] = 256'h0c0c0b0b0c0b0b0a0b0a0909090a0900000204030200090a0b0b080207050504;
    encBuf[242] = 256'h040303030100080a090901030504030101080a0c0d0d0b0d0b0b0c0a0a0a0909;
    encBuf[243] = 256'h0a080a090b0a0c0b0c0a0a080205060404040303030303020100080909090003;
    encBuf[244] = 256'h0505020200090c0c0c0c0a0b0b0a0a090908090b0d0c0c0a0b0a09090a0b0c0c;
    encBuf[245] = 256'h0b0b09010206040304020202020102040404050303020201080a0a0c0b0c0a0a;
    encBuf[246] = 256'h0a0a090909090b0b0d0b0b09000206030202090b0d0d0b0b0a0a090002030403;
    encBuf[247] = 256'h01080c0d0b0a0804060404030202010100000808080908080001030403030304;
    encBuf[248] = 256'h04030201080b0c0b080106040301000808010606040403020101010205030502;
    encBuf[249] = 256'h01000909090a0908080909090001040303000809080407070304030201000a0c;
    encBuf[250] = 256'h0c0c0a0a0a0909090a0b0b0b090a0a0c0f0d0c0b0a090001010100080a0b0908;
    encBuf[251] = 256'h0800090a0b090307070703020202020101020101000a0b0c0b09010307030202;
    encBuf[252] = 256'h08090b0b0b0a0a080909010407050404020108090c0b0b0b0b09090001020503;
    encBuf[253] = 256'h040402000008090808020102030101020108020b0d0c0f0e0b0d0c0a0b090801;
    encBuf[254] = 256'h04050305020101000809080908080801010305040304030201080809090b0a0c;
    encBuf[255] = 256'h0b0c0a0a000405050301010a0c0d0c0c0b0b0a0a080003040302080a0f0d0c0b;
    encBuf[256] = 256'h0d0a0a0b09090a0a090b00010407040304010000000003050603050302030302;
    encBuf[257] = 256'h020108090a0a08010506050303040100080a0c0c0d0b0b0c0a0b0a0a090b0c0c;
    encBuf[258] = 256'h0c0c0b0c0a0b0909080001030305030403020303020303050305030502030303;
    encBuf[259] = 256'h02010008090b0c0c0c0b0b0b0b0a0b0b0c0d0b0d0c0b0b0b0c0a0b0909080102;
    encBuf[260] = 256'h0203030301010800000204050504030503030303030301010100080101020303;
    encBuf[261] = 256'h0302000a0c0e0d0c0c0c0c0b0c0b0b0c090a0809000800080809090800010404;
    encBuf[262] = 256'h060305040303040202020101010001010000000a0a0b0c0c0b0c0c0c0c0c0b0c;
    encBuf[263] = 256'h0b0b0a0b0a09090801010102000000090908020406050303030100000a090800;
    encBuf[264] = 256'h020703050503040302040304040403040304020201010809080a090909090b0d;
    encBuf[265] = 256'h0d0c0d0b0d0b0b0b0c0a09090900080001000101030404050304030305020303;
    encBuf[266] = 256'h0303020202010000090a0a0c0b0b0d0b0c0b0c0c0b0c0b0b0c0a0a0a0a080800;
    encBuf[267] = 256'h00020103020203020203030303030403040203020108090c0d0c0b0c0b0a0a00;
    encBuf[268] = 256'h01040504040203030202010101020204040303030100090d0d0d0c0c0c0b0c0b;
    encBuf[269] = 256'h0b0a0b0a0a090a090a0808000103040504040403040403030304020202020101;
    encBuf[270] = 256'h01000808090a0a0c0b0c0c0b0c0c0b0b0d0a0b0a090a08090800080100000108;
    encBuf[271] = 256'h000000020505040403030402030303030503030303020201020201030101000b;
    encBuf[272] = 256'h0e0e0c0c0c0c0b0c0b0b0b0c0a0a0a0b0b0c0b0c0b0a09080001020304040304;
    encBuf[273] = 256'h0305030204020202020203030203010100080a0b0c0e0c0c0b0c0b0c0a09090a;
    encBuf[274] = 256'h09090b0a0c0b0b0c0a0b0a0b0a09080002020401020000080101050504040403;
    encBuf[275] = 256'h03050304030403030202020100000809090a0b0c0c0b0d0c0c0d0b0d0b0b0b0c;
    encBuf[276] = 256'h0a0a08090800010102030305020403030404040403040302030302010100080a;
    encBuf[277] = 256'h0b0e0b0c0b0c0a0c0a0c0a0c0b0b0b0c0b0a0909080001020402030303030204;
    encBuf[278] = 256'h030305040201020808090b0c0909010405040503020303020404050604040404;
    encBuf[279] = 256'h03030303010000090a0a0a0b0a0a0c0b0e0c0c0d0b0c0b0b0b0a0a0800000201;
    encBuf[280] = 256'h03030303050403050303050302040302030302020000080a0b0c0c0b0c0b0b0b;
    encBuf[281] = 256'h0b0c0b0b0c0c0b0b0b0b0b0a090801010204020303020201000a090c0c0a0b0b;
    encBuf[282] = 256'h0909090000080000090b0b0c0a00040707050403040203030101010008090909;
    encBuf[283] = 256'h0909090a0a0d0c0d0d0b0d0c0a0c0a0a0a090a08080000020203050204030303;
    encBuf[284] = 256'h05030304040302030303020108080b0c0c0c0b0b0b0a0b0a0a0a0a0a0b0b0c0b;
    encBuf[285] = 256'h090901030505040304030302010009090a0c0b0c0b0b0b0c0a09080801020103;
    encBuf[286] = 256'h02030405040404030403040304020101080a0d0c0d0b0c0a0b0b0b0b0c0b0b0b;
    encBuf[287] = 256'h0c0b0c0a09090801020404040203030203030402030202010108090a0a0c0c0b;
    encBuf[288] = 256'h0d0b0d0b0c0c0a0b0b0a0b0b0a0a090800010201020001010203050203010008;
    encBuf[289] = 256'h090b0a090e0b0e0d0c0a0b090001040403030402040403040402030202020101;
    encBuf[290] = 256'h010109090b0d0c0c0b0d0b0b0d0b0b0b0b0b0a090a0900000105040404040304;
    encBuf[291] = 256'h0203020202020303050203020101090a0c0d0c0c0b0d0a0b0a09090909090a0a;
    encBuf[292] = 256'h09090908010001020204060305030201080a0d0c0b0d0b0b0b0b0a0a09010204;
    encBuf[293] = 256'h0404020303020405040704040503050303040201010008090a0a0b0a0a0a0b0c;
    encBuf[294] = 256'h0d0c0d0b0d0b0b0b0a0a09080002020304020303030404030503040303040303;
    encBuf[295] = 256'h0302020200090a0c0b0d0b0c0a0a0b0a0a0a0a0b0c0b0c0a0b0a0a0908010203;
    encBuf[296] = 256'h0304030200000a0d0b0e0c0b0b0c0a0b09090801020203030303030404040504;
    encBuf[297] = 256'h04040403020303020000090b0c0c0b0b0b0b0c0b0b0c0b0d0b0c0b0c0b0b0b0a;
    encBuf[298] = 256'h0a08000203050305030402030203020302030305030503050203020100090a0c;
    encBuf[299] = 256'h0b0c0b0b0a0a09090908090b0b0e0c0c0b0a0a08000305030402020200000809;
    encBuf[300] = 256'h0a0b0c0b0a080206050403030303020302020203020102030304030501080c0e;
    encBuf[301] = 256'h0d0d0b0c0b0b0b0b0b0b0a0a0a090909090a0b0b0b0802070504040303030402;
    encBuf[302] = 256'h020202010109090a0a0b0a090a090c0d0d0b0d0b0b0b0c0a0b0a0b0909010104;
    encBuf[303] = 256'h02030100090b0b0c090a0a090a0b090801050304010a0e0c0c0a080205040503;
    encBuf[304] = 256'h020302030202010108090a090908010201090c0f0d0b0c0b0c0a0a0b0a0b0a09;
    encBuf[305] = 256'h000205040403040302030302030303030303040402020208090c0e0b0c0c0a09;
    encBuf[306] = 256'h0909080909090b09090a0808090b0b0c0c0a0a0901030404050201000b0e0d0c;
    encBuf[307] = 256'h0d0a0b0c0a090909080900000801040306050403040304050306040305030402;
    encBuf[308] = 256'h02020008080a0b0a0b0b0b0a0b0d0b0e0c0c0b0c0b0b0b0a0800020203040303;
    encBuf[309] = 256'h03030304040304030404020402020302010000090b0b0d0c0b0b0b0a0b0a0909;
    encBuf[310] = 256'h090a0a0c0b0c0b0b090901010203020100090b0c0d0e0b0d0b0c0c0a0a0a0808;
    encBuf[311] = 256'h01020305030403030303030303050404030403020200080b0c0c0b0d0a0b0b0b;
    encBuf[312] = 256'h0c0a0b0a0b0b0b0c0b0b0c0a0b09090801020405040404020303010101080800;
    encBuf[313] = 256'h000102030305030201000a0c0d0c0b0a0b080801020303030503030404020101;
    encBuf[314] = 256'h0000010104030402000a0c0d0d0c0b0c0c0b0c0b0a0908010102020203020403;
    encBuf[315] = 256'h0504030304020302040204020201090a0d0c0b0c0a0b0a0a0a0b0a0a0a09090b;
    encBuf[316] = 256'h0d0c0c0b0a0901020403030108090b0c0b0b0b0d0c0c0b0c0a0a090000000008;
    encBuf[317] = 256'h000103050504020302020203050404020300080b0d0c0c0b0b0b0b0c0b0c0b0b;
    encBuf[318] = 256'h0b0a090909090a090802060504040302030302030303020208090c0b0b0a0a08;
    encBuf[319] = 256'h080a0c0d0c0c0b0b09090908080808010305050403030201000000000000080a;
    encBuf[320] = 256'h0c0b0d0a090a08090c0c0b0e0a090002050403030303040303040301000a0d0c;
    encBuf[321] = 256'h0b0c0a090a090a0b0e0c0c0c0c0a0c0a0a0a0a09080800010202030305040504;
    encBuf[322] = 256'h040403050204030404040304030202010009090b0c0b0b0b0b0c0b0c0c0c0c0b;
    encBuf[323] = 256'h0c0b0b0b0a090801030403040303030402040303030403030303040302020200;
    encBuf[324] = 256'h090a0d0c0b0c0c0a0a0a090808000108090a0c0b0c0b0909000008080a0c0c0c;
    encBuf[325] = 256'h0c0b0c0b0c0b0c0b0a0b0a080002040504040304030303020202020303040402;
    encBuf[326] = 256'h0200080b0d0c0c0b0c0b0b0b0b0a0b0b0b0a0a0a0a0a0a0a0909000203050404;
    encBuf[327] = 256'h04040305030303020100080a0909080203060403030303020200000008000205;
    encBuf[328] = 256'h06040404020108090b0d0c0a0b0a0b0a0a0a09090908090a0c0b0d0a0a000306;
    encBuf[329] = 256'h0503040303030402030402010100090909090908090a0c0d0c0c0b0c0b0b0c0b;
    encBuf[330] = 256'h0b0b0b09000203050202010808090a0808080008090808010303080e0f0e0c0b;
    encBuf[331] = 256'h0b0a09080000020202040302040200080a0d0a0b0a080800000a0e0d0b0d0b0a;
    encBuf[332] = 256'h0a0a0b0b0c0c0a09080103040302030202040305030203030305040404030202;
    encBuf[333] = 256'h080a0c0d0b0b0a09080808080a09090900010108090c0a090107040503020201;
    encBuf[334] = 256'h0101020304030108090b0a0a020505030301080b0e0a0b0b0a0a0b0a0b090203;
    encBuf[335] = 256'h06040100080d0b0c0a09080000080b0d0d0c0b0b0a0909080a0d0c0b0c0a090b;
    encBuf[336] = 256'h090a0d0b0a0c0908090001080002040506050305040304050404040403030402;
    encBuf[337] = 256'h02000009090a0b0b0b0b0c0c0b0c0c0c0c0b0c0a0b0a09080002020403030304;
    encBuf[338] = 256'h020304020402030303020402030302030100090a0d0c0b0d0b0a0b0a0a080000;
    encBuf[339] = 256'h0000090b0c0d0a0b0b0a0a0a0b0c0d0b0d0b0b0c0b0b0c0b0b0b0b0a08000404;
    encBuf[340] = 256'h05040403040402030202010101010102010108090b0f0c0c0b0b0c0a0b0b0a0a;
    encBuf[341] = 256'h0a0a0809000000000000010102030402010100000203050503030200080b0909;
    encBuf[342] = 256'h0006050404040204030304030201000808080000020302000a0f0c0d0b0c0b0c;
    encBuf[343] = 256'h0b0b0c0a0b0a0a09080000010202030504050304040203040203020302010009;
    encBuf[344] = 256'h0c0b0d0c0b0a0b0b0b0a0b0b0b0b0b0b0b0c0b0b0a0a00020504040201000808;
    encBuf[345] = 256'h09090a0b0c0c0d0b0c0b0b0a0909000008000908000003070403040303040202;
    encBuf[346] = 256'h01000a0d0e0c0b0c0b0a0b0b0b0c0c0a0b0b0a09090909090008010404050403;
    encBuf[347] = 256'h03030302040202030101080909080002060202030100010800010808090f0d0b;
    encBuf[348] = 256'h0d0b0a0b0b090a0a090908020306050303030203050306040304030203020100;
    encBuf[349] = 256'h080b0b0d0b0c0a0a090809080809090a0d0b0b0c0a0900030604050403030302;
    encBuf[350] = 256'h00000a0b0c0c0b0c0b0b0b0b0c0b0b0d0c0c0b0c0b0b0a090001030603040304;
    encBuf[351] = 256'h02040302040305030603060304040302020101080a0a0b0b0c0b0b0b0c0b0c0c;
    encBuf[352] = 256'h0c0c0b0c0b0a0a09080101040303030402030303040303030403030304030304;
    encBuf[353] = 256'h0302010108090c0c0b0d0a0a0a09080001000009090c0d0b0d0b0b0c0b0b0c0b;
    encBuf[354] = 256'h0b0c0b0a0a0a0a0b0b0a0b0a0900020706030603040304020201010000000808;
    encBuf[355] = 256'h080808090a0b0c0c0c0b0b0b0b0b0b0a0a090800010203030302000c0c0e0c0b;
    encBuf[356] = 256'h0d0b0c0a0b0a0909000100010008080102060604050503050303030302020008;
    encBuf[357] = 256'h090a0a0b0b0b0b0b0a0b0d0d0c0b0c0b0a0a0908000101020203010200080a0a;
    encBuf[358] = 256'h0d0b0b0c0b0b0b09010307060304030303020000000801010305030403020100;
    encBuf[359] = 256'h0a0c0c0c0c0c0b0c0b0c0a0b0c0a0b0a0a0a0a0a090809080a0b0a0a01040704;
    encBuf[360] = 256'h03040202010009090a0a0a0a080002020202080809090b090b0c0a0b0c0b0d0f;
    encBuf[361] = 256'h0d0c0c0b0c0b0a0c0a0b0c0b0c0a090800010304040304020303020402040304;
    encBuf[362] = 256'h03040202020008090b0b0c0b0b0b0b0c0c0b0b0b0c0b0a0c0a0b0a0a09080003;
    encBuf[363] = 256'h04040404020303030403020100080b0c0b0a0a00010001020104060405040203;
    encBuf[364] = 256'h02000100000103040402010a0e0d0d0b0c0b0b0a0a0b0b0b0b0b0b0b0a0b0e0b;
    encBuf[365] = 256'h0c0c0a0909000204050403050305030305030304040305040304030302010009;
    encBuf[366] = 256'h0b0c0c0c0a0b0a0b0a0b0c0b0d0b0b0c0b0a0a09000203060304020303020202;
    encBuf[367] = 256'h0203030203030201030202040203020100090a0c0b0b0b0a0803040603020208;
    encBuf[368] = 256'h0c0e0c0d0c0b0c0b0c0b0c0c0a0b0b0a0a0a0809000000020204040404040304;
    encBuf[369] = 256'h040303030202010008090a0b0c0a0c0a0c0b0b0c0a0b0a090908000001010302;
    encBuf[370] = 256'h04030304020108090c0d0c0d0b0d0b0b0b0c0a09090801010304030404040304;
    encBuf[371] = 256'h030403030402020101010808080809090a0b0b0d0d0b0c0c0b0b0b0b0a0a0800;
    encBuf[372] = 256'h020202030303040203030503040402030202010000000809090b0e0c0b0b0c0a;
    encBuf[373] = 256'h08080002030402020200080a0e0c0d0c0b0b0b0a0b0a0b0d0a0b0c0a0a0a090a;
    encBuf[374] = 256'h090000030603050303030402020201000108080809090a0c0c0c0c0b0c0b0d0b;
    encBuf[375] = 256'h0c0b0c0b0b0b0d0b0a0c0a090a0909090909090a080808000008010001040101;
    encBuf[376] = 256'h010a09010407070503050203040202030202010001000000080b0d0d0e0b0b0d;
    encBuf[377] = 256'h0a0b0a0b0a0a0a080802040404050304030203030201000809090a0a0b0c0b0c;
    encBuf[378] = 256'h0b0a0b0b0b0a0a090304060404030403030302020100090a0c0c0b0d0a0a0a09;
    encBuf[379] = 256'h09080a0b0c0d0b0b0b09090808080a0a0a0a0a00090d0d0c0d0b0b0a08010305;
    encBuf[380] = 256'h040403040402050404050504040403040303010100090a0b0c0b0b0b0b0b0c0c;
    encBuf[381] = 256'h0c0c0b0d0a0b0a09090001020403040303030203020303030303020101010102;
    encBuf[382] = 256'h04030503030101090909090002050404020200080b0c0e0b0d0c0b0c0b0b0c0c;
    encBuf[383] = 256'h0b0c0b0b0c0a0908080001020201020303060403040304020302020101080909;
    encBuf[384] = 256'h0b0c0b0c0b0b0c0a0a0a090002040603050302020100090a0a0c0c0b0b0d0b0c;
    encBuf[385] = 256'h0b0c0b0c0b0b0b0b090900020404040304030404040304020302020000080a0a;
    encBuf[386] = 256'h0b0c0b0c0b0b0c0b0c0b0a0c0a0a09080104050404030303020100000009080a;
    encBuf[387] = 256'h0b0c0c0c0b0b0a0b0a0a090908000203070403040303030203010100080b0e0c;
    encBuf[388] = 256'h0c0c0b0b0a0a0b0a0a0b0b0a0b090001040404030503030303030100090a0a0c;
    encBuf[389] = 256'h0b0c0b0c0c0c0b0c0c0a090a0800000101020203040304030304020100090a0d;
    encBuf[390] = 256'h0d0c0c0c0b0b0c0a090a0a0a0a0a090800040405030502030304030203020101;
    encBuf[391] = 256'h08080a0c0b0d0c0b0c0b0b0b0a0a080800020303040503040303040201000808;
    encBuf[392] = 256'h09090908090a0d0d0c0c0a0b0a0a090908090001030504040305030303030302;
    encBuf[393] = 256'h01080a0c0c0b0b0a0a0b0b0c0d0c0b0b0b0a0900010201010000000102040303;
    encBuf[394] = 256'h01010a0d0d0c0d0c0c0c0c0a0b0a0a0800010103030503040403040403060405;
    encBuf[395] = 256'h04040403040202020808090b0c0b0a0b0a0a090b0b0e0b0d0b0c0a0a0a080002;
    encBuf[396] = 256'h0305030303020301020102020202010102020305030404030203010000090a0a;
    encBuf[397] = 256'h09080104030402010a0d0d0d0c0b0b0c0b0b0b0d0b0c0c0b0c0b0a0a0a090808;
    encBuf[398] = 256'h08000101020404040303040303030302010008090908090008090a0d0c0c0b0a;
    encBuf[399] = 256'h0901050504040203010108090b0d0b0d0b0c0b0c0a0b0b0b0c0a0b0a0a000104;
    encBuf[400] = 256'h040403040303040304030403030302010009090b0c0c0a0b0a0b0a0b0a0a0a0b;
    encBuf[401] = 256'h0b0a0a080205060403040202000008080909080909090b0d0b0b0c0a09080103;
    encBuf[402] = 256'h060405030403030202010008080a0a0b0e0b0e0b0c0c0b0a0b0c0a0b0a0b0a0a;
    encBuf[403] = 256'h090800010101010202060305030303010108080a0b0b0c0c0b0b0c0b0c0a090a;
    encBuf[404] = 256'h080000000108080008000200080a0f0c0d0c0b0c0c0c0b0d0b0b0c0b0b0a0a08;
    encBuf[405] = 256'h0800020204040204030403040304030304020201010108000809080909090900;
    encBuf[406] = 256'h01000101090a0c0d0c090a09000101030101010002050305030208090d0b0a09;
    encBuf[407] = 256'h0802000a0d0f0d0b0b0a010505040402030202020102030100080c0b0c0d0a0b;
    encBuf[408] = 256'h0b0c0b0c0a0a090801010202010008000803060405030200090c0f0a0a0a0908;
    encBuf[409] = 256'h090a0d0d0c0b0a0b090000020202030204040605050604040404030303020100;
    encBuf[410] = 256'h090a0c0b0b0b0a0b0a0a0b0d0c0c0c0b0a0b0908000204040304030202010100;
    encBuf[411] = 256'h0800080808080008000002030404030302020102030404050403030402020008;
    encBuf[412] = 256'h0b0d0c0c0b0c0b0c0b0b0c0b0c0b0c0a0b0a0a0a080900080001020306030404;
    encBuf[413] = 256'h0202020001080008090808000001020204020103010003050505040304030201;
    encBuf[414] = 256'h08090c0d0c0b0c0b0c0b0a0b0b0b0b0a0a0a0901020405040403040203020303;
    encBuf[415] = 256'h04030303020200080b0c0d0b0b0a0a0900020303050202010101030705050403;
    encBuf[416] = 256'h04020100090b0d0c0b0b0c0a090a090a09090909080001020404050404030203;
    encBuf[417] = 256'h010108090b0b0c0d0b0b0d0b0b0b0b0909000203040303040202010200000809;
    encBuf[418] = 256'h0a0b0e0c0b0e0b0d0b0b0c0a0a09090800000100020203040404030303030301;
    encBuf[419] = 256'h0008090b0c0b0d0a0b0c0a0b0b0b0b0a0b0c0a0b0a0901020404030303010001;
    encBuf[420] = 256'h0001020008080b0b080903060202020a0a090c01050307030202030101030203;
    encBuf[421] = 256'h040101020808010900050205050202010a0e0d0d0c0c0c0b0b0b0b0a0a0a0908;
    encBuf[422] = 256'h0801010203030404010203010303010102090a0a0f0b090c0a00000506040305;
    encBuf[423] = 256'h030203010000090b0b0c0c0c0c0c0b0d0c0b0b0c0a0a09090900000800010001;
    encBuf[424] = 256'h0202050404040403060405040404040403040202020008090a0b0c0b0a0a0b0a;
    encBuf[425] = 256'h0a0b0d0b0d0b0c0a0a080001040305030303010108080a0a0a0b090909080100;
    encBuf[426] = 256'h0203040404030403030503030404020303020108090b0e0c0b0d0b0b0b0c0b0b;
    encBuf[427] = 256'h0c0b0c0a0b0b0b0a0a09080800010102020201030203030201010a0b0e0b0b0a;
    encBuf[428] = 256'h0908010104030404040405030504030503040203020108090a0d0c0b0c0b0b0a;
    encBuf[429] = 256'h0b0b0b0b0b0a0a08000306040404040303020302010008000908090809090a09;
    encBuf[430] = 256'h0a09090800020406040403040302020202020202030100090d0d0c0c0b0b0a0a;
    encBuf[431] = 256'h09080001030404040304030303040304020301000b0d0d0d0b0c0c0a0b0b0b0a;
    encBuf[432] = 256'h0b0b0b0b0a0b0a0909090801010203030201010808090809090b0c0c0b0c0909;
    encBuf[433] = 256'h080101010201080c0d0d0c0b0a0a0908010000090a0b0c090900080a0d0d0c0c;
    encBuf[434] = 256'h0b0a0b0c0b0d0d0d0b0c0b0b0a0a090900000304050404030304030304030504;
    encBuf[435] = 256'h0203030201010100010101020000080b0b0c0d0b0b0d0b0b0b0b0a0b0a080901;
    encBuf[436] = 256'h030604050303050202020208080a0d0c0b0d0b0b0c0c0b0b0c0b0a0908000203;
    encBuf[437] = 256'h03050302030101000a090a0a09010205050302000a0f0c0d0b0c090900010203;
    encBuf[438] = 256'h0202090b0e0d0b0c0b0b0a0a090808000808090a0a0a08010407050504050405;
    encBuf[439] = 256'h0305040304030203020108090b0c0c0a0b0a090a090a0a0c0b0c0b0b0a090103;
    encBuf[440] = 256'h0604040303020108090b0d0b0b0b0a0908010304040304030303040302040303;
    encBuf[441] = 256'h0304020201000a0c0c0c0c0c0b0a0b0b0a0a0a0a090a0a0b0c0b0c0a0b0a0909;
    encBuf[442] = 256'h0900000800080a0a0c0e0b0d0b0c0b0b090a0800020305040203030303030403;
    encBuf[443] = 256'h0404040304040304020100090b0e0b0c0b0b0b09090000010001080008080002;
    encBuf[444] = 256'h05050404030303020000090b0a0c0a0b0a0b0b0b0b0a09000306040503040303;
    encBuf[445] = 256'h02020108000900000103030301090d0e0c0c0b0a090002040504030302030101;
    encBuf[446] = 256'h000100010008090b0e0d0c0c0c0b0c0c0b0b0b0b0c0a090a0908080801000000;
    encBuf[447] = 256'h08090a0b0d0b0c0b0b0b0b0b0c0c0b0b0d0a0b0a080001030503050303030202;
    encBuf[448] = 256'h0109090a0b0a0808000108090a0d0b0b0e0b0d0d0c0b0c0b0b0b0c0b0c0a0b0a;
    encBuf[449] = 256'h0908000103010203040405020303010101080801090801000106030505020203;
    encBuf[450] = 256'h030403010102090002010406030403040203020100090b0c0c0a080801020108;
    encBuf[451] = 256'h090d0d0d0d0b0c0c0a090900010101080b0c0c0c0a0808020503050402030201;
    encBuf[452] = 256'h010009090a0a0b090b0a0a0c0b0c0c0b0c0a0b090a09090908090a0a0c0c0b0d;
    encBuf[453] = 256'h0b0b0c0a09080103030404030306030406030504050404040404030403030202;
    encBuf[454] = 256'h0100090a0b0c0c0a0a0a0909090a0b0c0c0b0b0b0a0003050504030203000809;
    encBuf[455] = 256'h0b0e0b0b0b0a09080203060403030302030102010101020203020301080b0f0d;
    encBuf[456] = 256'h0b0d0c0a0b0a090a080800080008090b0c0b0d0b0a0b0a0b0b0b0b0c0a0a0909;
    encBuf[457] = 256'h0900090a0a0d0b0b0b0a0103050502010009090a090800020406040504040402;
    encBuf[458] = 256'h030101090a0c0c0b0c0a0a090000020202020008080800030704040402030302;
    encBuf[459] = 256'h00080a0c0c0c0b0b0a090908000808090800000103040302030108080a0b0901;
    encBuf[460] = 256'h03070503030200080a0c0b0b0a09010407040404030302030303040304020201;
    encBuf[461] = 256'h090a0c0e0b0e0b0c0c0b0b0c0a0b0a0a0a0a0908080808090a0b0b0d0b0b0a0a;
    encBuf[462] = 256'h0a090908090b0b0e0b0a09000206050304040304030302030201000000010102;
    encBuf[463] = 256'h040101080e0c0d0c0c0b0b0b0a0b0a090b0a0a0a0b0a0a090908000102050503;
    encBuf[464] = 256'h0503010100080002030704040403030303020203010303050304020201000000;
    encBuf[465] = 256'h080001090b0c0f0b0c0d0a0b0a0a09000103020404020202030204010008090a;
    encBuf[466] = 256'h0b0c0b0c0c0b0b0b0a09090a0b0e0c0a0a080305050402020000090a0a0a0a0a;
    encBuf[467] = 256'h0a0a0d0b0b0d0a090908000b0c0e0d0d0b0d0b0a0b0808010403040302020100;
    encBuf[468] = 256'h0809080103040604030304020403040503050403050303030402010008080a0b;
    encBuf[469] = 256'h0b0b0c0c0a0a0b0a0b0a090800020306040503040303040202010108090a0b0b;
    encBuf[470] = 256'h0a0a08010102030100090a0a0908040405040304030303040108000a0c0b0d0b;
    encBuf[471] = 256'h0b0c0c0b0b0e0c0b0d0b0c0b0a0a090900000202030304030303020303010108;
    encBuf[472] = 256'h0b0d0e0d0b0c0c0b0b0b0a0a0a080000020304050303050202020000080b0c0b;
    encBuf[473] = 256'h0d0c0a0b0b0a0a0908000102030503050404030403030202010000080a0a0c0c;
    encBuf[474] = 256'h0b0b0c0b0a0a0a0a0b090909080808000001040303050101080a0c0b0e0c0b0b;
    encBuf[475] = 256'h0c0b0a0900010205030403030404040404030402020200090a0c0e0b0d0b0c0a;
    encBuf[476] = 256'h0b0a0a0909090a0a0a0c0b0a0b09090808090a0c0b0d0b0b0b0b0b0d0a0a0b09;
    encBuf[477] = 256'h0900020405050404040203030201020202020100090a0e0b0d0b0c0c0a0b0c0a;
    encBuf[478] = 256'h0a0b090a0a0a0a0a0b0a0a0801040505040203020101090a0a0c0a0908020404;
    encBuf[479] = 256'h04030302010008000102060305030403030201000b0c0d0c0a0b090a09090b0b;
    encBuf[480] = 256'h0d0b0c0a0b090a0800010306040404030204020202020202020008090a0b0c0c;
    encBuf[481] = 256'h0a0c0b0a0c0b0a0b0b090a09080a0c0b0f0b0c0c0b0b0b0c0a0a0b0a0c0b0a0c;
    encBuf[482] = 256'h0c0a0a0a0908090108010205040603030303010200000100010202020208090b;
    encBuf[483] = 256'h0f0c0c0b0b0a0802060504050304030302030101000808080802020203010000;
    encBuf[484] = 256'h0801060505040403040303040304040203030203020102020102010201010000;
    encBuf[485] = 256'h090a0b0b0d080003070503050303030402020102010200010008090c0e0c0c0c;
    encBuf[486] = 256'h0b0b0b0a0a0a09090801020306030303020101090b0d0d0d0c0c0b0d0b0b0a0a;
    encBuf[487] = 256'h0a0808080008080008000102020200080a0c0b0c0c0a0b0b0b0b0b0c0c0c0c0b;
    encBuf[488] = 256'h0b0b090103050403020201000809090c0b0d0b0b0b0a080809090b0d0c0b0a00;
    encBuf[489] = 256'h040505030403020100080909090002040404010108090a080105060304040102;
    encBuf[490] = 256'h00080a0a0a0b090900010202040200080e0d0d0c0c0b0a0a0a090a0a0c0b0b0b;
    encBuf[491] = 256'h0a0a080102030503030403010201000a0a0e0c0b0d0a0b090800020306020402;
    encBuf[492] = 256'h030203010202000008090a090b080800010108090d0f0c0c0c0b0b0b0a090801;
    encBuf[493] = 256'h0204030300080a0d0c0a0c0a0a0b0c0b0d0b0909010204030303050304040302;
    encBuf[494] = 256'h020009090a0a0c0b0e0b0c0b0b0b090909090809090000010002020307060404;
    encBuf[495] = 256'h0304040201020008080a0c0a0c0b0c0b0d0b0d0c0a0b0b0b0909010103040203;
    encBuf[496] = 256'h0200010001020503030302000a0d0c0c0b0b0a0a0b0c0b0c0c0b0a0b09080004;
    encBuf[497] = 256'h0604040403030202010202020404030305020303030202020100010305050404;
    encBuf[498] = 256'h04030302040103030304040303050204030204020202010100080909080a0001;
    encBuf[499] = 256'h04060403040303030303040402040203020301020109090a0d0a0a0b08090901;
    encBuf[500] = 256'h0100030108000b0f0d0c0b0a0909010200020a0e0c0d0c0b0c0b0a0b0c0b0b0d;
    encBuf[501] = 256'h0a0a0b08090908090a0c0c0b0c0b0c0b0b0b0b0c0b0a0b0a0a0b0d0a0b0b0909;
    encBuf[502] = 256'h0901000801000001090c0c0f0c0a0b0b08080002010008090c0b0e0c0b0c0b0b;
    encBuf[503] = 256'h0a0900010405030402020000080a0a0a0a0a0a090908080809090c0c0d0c0c0b;
    encBuf[504] = 256'h0d0b0a0900030505040202020100000102030504030302020109090d0c0d0c0b;
    encBuf[505] = 256'h0c0b0c0a0b0a0a0a090a0909090a0b0d0c0c0b0c0a0b09090801020502030300;
    encBuf[506] = 256'h080a0d0b0c0b0a090808000809080b0a080005060403030208090e0b0d0b0b0b;
    encBuf[507] = 256'h0a0908000001090c0c0d0b09080205050305010200080a0a0c0c0a0a09000002;
    encBuf[508] = 256'h020208080c0c0c0b0b0a0a0800010206030403040204010202020101090a0a0d;
    encBuf[509] = 256'h0a0808010403020308090b0f0b0a0a09020206050203030008090c0c0a0a0901;
    encBuf[510] = 256'h0306040301010b0c0d0d0a0b0a08000002030302020108080809000908000c0c;
    encBuf[511] = 256'h0c0e0c0b0c0b0a0b0b0b0a0b090b090808020204050504040403030302010008;
    encBuf[512] = 256'h0800000305030503020201080808000307060403040304020202030203040302;
    encBuf[513] = 256'h0403030403030303020100080809080002020404030504040405030403040302;
    encBuf[514] = 256'h0101000808080900000800090c0c0c0b0c09090003050404030203010108090a;
    encBuf[515] = 256'h0c0b0b0c0b0a0b0a0b0d0d0b0c0c0b0a0b090a0a0a0a0c0a0c0b0a0a0a090909;
    encBuf[516] = 256'h090a0c0b0e0c0a0c0a0a0b0b0a0b0c0a0c0a0a0b09090801020202000c0f0d0c;
    encBuf[517] = 256'h0c0a0a09080102030301080a0d0c0b0a0900020404030302080a0e0d0c0b0b0b;
    encBuf[518] = 256'h0a09080801010101030303040201090c0c0c0a08010504050202080b0f0c0d0b;
    encBuf[519] = 256'h0c0a0a08010404050303030200090b0c0c0b090900010304030201080b0d0c0b;
    encBuf[520] = 256'h0a0a080205040403030200090b0e0b0c0a0a0800010402040201010809090b0b;
    encBuf[521] = 256'h0b0b09080001020301010008080003070404040302030100090a0c0c0c0b0b0b;
    encBuf[522] = 256'h0a09080800000808080800010303050200000b0e0b0e0c0b0b0c0a0b09090808;
    encBuf[523] = 256'h0000000101030504050304030304020201010108090809080102050403040303;
    encBuf[524] = 256'h03020203010100080808000207040305020200000a090a080103060404020201;
    encBuf[525] = 256'h00080a09080003060504040402030202010008090b0b0d0c0b0c0c0b0a0a0900;
    encBuf[526] = 256'h0103050203020101010001010002040305050404030402020101080800010205;
    encBuf[527] = 256'h050304040204020302040202030303030303020102000801010002020001080b;
    encBuf[528] = 256'h010203070707040302040202010108080808080100040403050302020109090b;
    encBuf[529] = 256'h0d090908040405040302020108080b0d0a0c0b0a0b0c090a0a09090a0a0b0e0a;
    encBuf[530] = 256'h0c0c0a0a0b0a0a0a090a09000909080b0e0b0e0c0b0b0c0a0b0a09090a090c0c;
    encBuf[531] = 256'h0b0d0c0a0b0b090a080000020200080a0f0d0c0c0b0c0b0b0b0b0b0b0a090908;
    encBuf[532] = 256'h08090a0b0e0b0d0a0c0a090a0a090a09090908080002020304010000090a080a;
    encBuf[533] = 256'h090a0f0e0c0c0b0b0b0a09090a090b0d0a0c0b0a0c0b0c0b0c0a0b0800020505;
    encBuf[534] = 256'h0404030304020202010000080b0a0b0b0a080104040303030001000801030505;
    encBuf[535] = 256'h050304030301000a0d0c0d0a0b0a090808000009090a0d0c0b0b0b0808020503;
    encBuf[536] = 256'h0503020303020305020403010201090a0c0d0b0b0c0b0a0b0b0b0d0a0a090802;
    encBuf[537] = 256'h03040401090c0f0c0c0b0c0a0a0a09080801080000090b0c0d0b0a0908030405;
    encBuf[538] = 256'h040303020201010000000000020102050101020001010101040800000c0a090a;
    encBuf[539] = 256'h00030102020b0b0b0f0d0a0c0b0a0d09080a0000080103030706030404030403;
    encBuf[540] = 256'h0304020303030303040202030203030304030102010001010307040405030304;
    encBuf[541] = 256'h0303040203020302030302020202040306040404030402030203030204030403;
    encBuf[542] = 256'h0503030503040402020100000a0b0b0d0a0a0909000000020000010001020504;
    encBuf[543] = 256'h040402030008090c0d0a0b0b0a0a0a0a0a0c0a0a0b0b0b0b0001040704030402;
    encBuf[544] = 256'h00000a0b0c0b0c0b0a0b0a0b0b0c0d0c0c0c0b0c0a0a090909080a0b0c0b0a09;
    encBuf[545] = 256'h09000100090a0e0b0c0c0a0a090800000101080a0c0e0c0b0b0b0b0b09090800;
    encBuf[546] = 256'h020202040100080b0d0b0e0c0b0c0c0b0c0c0b0c0c0a0b0a0908000001010100;
    encBuf[547] = 256'h00010203040301080a0d0c0b0b0a090001030503030201080a0d0b0b0c0a0909;
    encBuf[548] = 256'h0908080801090a0a0f0b0a090104040303080808000507030303090b0e0c0a09;
    encBuf[549] = 256'h0105050404030303030102000808080801020404030300080d0c0d0c0a0b0b0b;
    encBuf[550] = 256'h0a09080001030304030302010100000808010406050505030303030108090a0b;
    encBuf[551] = 256'h0b0a0a0808010203040202020201020103050404050305020200080c0c0d0c0b;
    encBuf[552] = 256'h0b0c090a090800080000090a0a0c0b0b0a090000020304040403040302040203;
    encBuf[553] = 256'h04040303030108090b0a0a00030504030300090d0d0d0c0b0b0c0a090909090a;
    encBuf[554] = 256'h0b0b0c0a0a09000003060306030402020100080a090808020301020101030707;
    encBuf[555] = 256'h0405030303030202010102020304020403040404030502020202010000000001;
    encBuf[556] = 256'h0002030204040204030403040203040204030405030305030202020008080a0a;
    encBuf[557] = 256'h0b0c090a0800020104020008090c0b0c0c0a0a0a0001010302080a0f0e0c0c0c;
    encBuf[558] = 256'h0a0b0b0a0909000000010809080b0a09000003040204020101090c0c0e0c0b0c;
    encBuf[559] = 256'h0b0b0b0d0c0c0c0b0b0c090a09090a0b0b0d0b0b0a0b0a0a0b0a0b0b0b0c0c0b;
    encBuf[560] = 256'h0c0b0c0b0b0b0b0b0b0a090908090b0c0c0b0a000406030301090e0d0b0d0a0a;
    encBuf[561] = 256'h0a0809090a0b0c0c0c0b0b0a0b0a090801020304050202030001080808000908;
    encBuf[562] = 256'h090e0c0c0c0b09090802020201080a0c0c0b080903060405030402030100090a;
    encBuf[563] = 256'h0b0b0c0a090908000a0a0b0e0b0a0b0900000002080104030706030504030302;
    encBuf[564] = 256'h0208080a0b0a0c0a080900020100000c0d0c0d0c0b0b0c090909090909090909;
    encBuf[565] = 256'h0100020300090a0f0b0b0b0b080a0a000a09020808020d0d0b0e0a0102070603;
    encBuf[566] = 256'h040303010100090a0a0908090800090b0b0f0b0a0b0c0a0d0b0b0b0b09080206;
    encBuf[567] = 256'h0305040202020101000808090908010405050304030302010800080001040404;
    encBuf[568] = 256'h0304030302030302040203040305040305020301010100000002040304020100;
    encBuf[569] = 256'h090a0a0a00030704040402020301010101020203040403050403040402030202;
    encBuf[570] = 256'h010100010101020303050402040304030302020109090b0c0a090a0801020505;
    encBuf[571] = 256'h0304040103010808090b0b0d0b0c0b0b0b0b0b09090b0a0c0c0a0a0a02040406;
    encBuf[572] = 256'h030101080b0c0c0c090900010108090c0f0b0c0b0b0b0c0a0b0c0a0c0a0b0a0b;
    encBuf[573] = 256'h0a09090002030703040303010208090a0b0b0a0b0a080c0c0c0e0c0a0c0a0a09;
    encBuf[574] = 256'h090800000808090b0e0b0c0a0a080103040301000b0f0c0d0b0b0c0a0b0b0a0a;
    encBuf[575] = 256'h0a0a090908080809090b0b0c0a09080801080b0c0f0b0b0b0a00000203010809;
    encBuf[576] = 256'h0d0b0a0b09000909080e0b0c0c0b0b0d0c0c0c0c0b0b0c090909010002020101;
    encBuf[577] = 256'h0009090909000504050503020200090a0d0b0a0a090002030603050302030301;
    encBuf[578] = 256'h010009090000030703040401010108090808000200090a0f0f0b0c0b0a0a0800;
    encBuf[579] = 256'h010103010201000001010104030406020303020100090b0a0c09020306050202;
    encBuf[580] = 256'h010a0b0d0d0b0a0b0a0a0a0b0b0d0b0c0c0b0a0b090100020301080a0f0b0a0b;
    encBuf[581] = 256'h0003050504020300080a0b0c0b0a080206040402030202000000090001000203;
    encBuf[582] = 256'h0404030203020001090901000407050306020303020203010203020305020504;
    encBuf[583] = 256'h0304050305030303030202010001020204050304040204020204020303040303;
    encBuf[584] = 256'h030203030203020102000808080a000000070403050402030202020301040402;
    encBuf[585] = 256'h05020203010000080a08090a000009030201050108000b0f0c0c0d0a0a0b0b0b;
    encBuf[586] = 256'h0d0a0c0b0c0b0d0b0b0d0a0c0a0b0a0b0a0a0a090a0b0a0b0d0b0c0b0b0b0908;
    encBuf[587] = 256'h0001030101080b0f0d0c0c0b0c0a0b0a0b0a0a0c0a0c0c0a0b0b0a0a0a090908;
    encBuf[588] = 256'h0909090a0d0c0b0e0b0b0c0b0b0c0a0b0a0b0b0b0b0a0a0a0808010201030304;
    encBuf[589] = 256'h05030504020302000a0a0f0c0b0c0b0a0a0a09080a090d0c0b0d0b0a0b090000;
    encBuf[590] = 256'h00020808090d0b0b0c0b0a0909080800010808000a09080a0904020607020403;
    encBuf[591] = 256'h030204010204020404020201080b0b0e0a090900020101010b0c0c0e0a090900;
    encBuf[592] = 256'h030305050202020101010101020202050203040204030203030201020808010a;
    encBuf[593] = 256'h09010903070405050203040001080a0b0b0c0a090801030302020b0e0c0e0b0a;
    encBuf[594] = 256'h0b090800000208080b0f0c0b0c0b0909000200010109090a0b0a020206050202;
    encBuf[595] = 256'h02080a0a0e0a0a0b09090a09090c0c0b0d0b0b0c0a0a0a08000800010808090a;
    encBuf[596] = 256'h0804060705030503020201000008000304050404020303020202010203040403;
    encBuf[597] = 256'h0404020304030403050303030403030304030403030303030403030304020302;
    encBuf[598] = 256'h0201020103050504040304030303030303050304040204020202030102020202;
    encBuf[599] = 256'h020103020003030305040104030102020001000a080b0f0a0b0e0b0b0d0b0b0c;
    encBuf[600] = 256'h0b0b0d0a0b0c0b0a0c0a0b0b0b0c0c090a0b08090900090b0a0e0c0b0b0d0a0a;
    encBuf[601] = 256'h0a0a0a0b0b0d0c0b0c0c0a0b0b0b0b0c0a0a0b0b0b0c0b0c0b0c0b0c0b0c0a0b;
    encBuf[602] = 256'h0b0a090a09000908080a0a090b0b080a0801000205020202090c0d0f0b0c0c0b;
    encBuf[603] = 256'h0a0b0a090800010102020002000908080900000103030103080d0d0e0d0c0b0c;
    encBuf[604] = 256'h0a0b09080002040403040201010809090a0900020307030204010000090b0c0c;
    encBuf[605] = 256'h0c0a0a0801010202090d0e0e0b0c0b0a090900000000080a0a0a0b0a00080103;
    encBuf[606] = 256'h0405040202040203040201020909090a0a000103070202020009080d0c0b0d0b;
    encBuf[607] = 256'h0a0a090101010408090a0f0b0b0c0a08000803000800090b0203060705020302;
    encBuf[608] = 256'h02010008020204070304040202030000000a0a090b0a00090a010a0d0a0e0c0b;
    encBuf[609] = 256'h0c0c090b0a080a09090c0a0a0c09080800020008090f0b0c0d09090901040204;
    encBuf[610] = 256'h030101000b0a0c0d09090800030205030304010108090b090a08060505050304;
    encBuf[611] = 256'h0302020101010002030405040303050202030202030202040302050304040303;
    encBuf[612] = 256'h0403020302010302020304030504020403020303020202010201020403040503;
    encBuf[613] = 256'h0204010100000900080803010305010101090a0a0e0b0a0c0a0a0c0b0b0e0c0a;
    encBuf[614] = 256'h0c0b0a0c0a0b0b0c0b0e0a0b0d0a0b0b0c0a0a0b0a0c0a0b0d0a0b0c0b0a0b0b;
    encBuf[615] = 256'h0a0c0b0b0c0b0b0c0b0b0d0a0a0b0b0a0c0a0a0c0a0b0c0b0b0c0b0a0b0a0a0c;
    encBuf[616] = 256'h0a0a0c0b0a0b090909010008080a0d0b0c0c090909080008000909080a0b0a0c;
    encBuf[617] = 256'h0a090b0803020507020303000800090804030705020304020001000001010304;
    encBuf[618] = 256'h020402080a0a0f0b0a0b0a00000102000a080f0b0a0c0a080a09010a0a090d0c;
    encBuf[619] = 256'h090d0b0a0c0c0b0c0b0b0b0b0a0b0a090c0c0a0d0b0a0b0a0008000401010308;
    encBuf[620] = 256'h00000909000a0804000607020404020202000000090002020605030403020302;
    encBuf[621] = 256'h0002020204050304030303040303050203030001080a09000004060303050101;
    encBuf[622] = 256'h0108000800010304040402030302020302040303040304030502020302030208;
    encBuf[623] = 256'h08080b0b0c0c0b090908020304040100080b0b0c0b08020506030201080c0c0d;
    encBuf[624] = 256'h0c0a0b0909090808090801010207030405030404030404020402030203030304;
    encBuf[625] = 256'h0403050203040201020202030305050204020302020203030305040204030204;
    encBuf[626] = 256'h0303050303040302030203030404030502030302030201030402040302040101;
    encBuf[627] = 256'h02020104030205020101000a000909020302050209000c0e0a0b0c0a0a0b090b;
    encBuf[628] = 256'h0e0a0b0d0a0b0c0b0b0d0b0b0c0b0b0c0a0b0b0b0d0b0b0d0b0b0b0d0a0b0b0b;
    encBuf[629] = 256'h0d0b0c0b0b0c0b0a0b0c0b0b0c0b0c0b0b0b0b0b0c0b0b0c0b0b0a0c0a0a0a0b;
    encBuf[630] = 256'h0a0d0a0b0c0b0a0a0908090808090b0c0c0a0c09080801030303040108080a0a;
    encBuf[631] = 256'h0a0b090008020502030502020401030201020300040602060403030502020201;
    encBuf[632] = 256'h02040204040204030204030202030101010909090b09000003060102080b0d0d;
    encBuf[633] = 256'h0c0b0b0a0a080808080b0c0c0c0c0a0c0a0a0b0c0a0b0a0a0908010101000b0e;
    encBuf[634] = 256'h0c0d0b0a0a080303040301080b0f0c0a0c0a090909080909090a0a080a0a090d;
    encBuf[635] = 256'h0c0b0e0a090800030204030008090c0908000306030303010102000307020304;
    encBuf[636] = 256'h0101010900030207050303040201000000010102040202020008010002050202;
    encBuf[637] = 256'h030800010005070504040202020000090a090800020403040302010108080008;
    encBuf[638] = 256'h0003040603040403030402010008090a0c0b0d0a0a0900020404040302020100;
    encBuf[639] = 256'h0103040706040305020303010202010303040503040304030303030303040303;
    encBuf[640] = 256'h0403050204020302030302040103030304030303030203050204040203020101;
    encBuf[641] = 256'h000800020207040304030202000000080001020103000b0b0f0d0b0c0c0a0c0b;
    encBuf[642] = 256'h0b0c0b0b0c0b0b0c0c0b0c0c0b0b0b0b0b0b0a0c0b0c0c0b0b0d0b0a0b0a0b0a;
    encBuf[643] = 256'h0b0b0c0c0b0c0b0c0b0c0b0b0b0b0b0c0a0b0c0b0c0b0b0d0a0b0b0a0a0a0a0a;
    encBuf[644] = 256'h0a0b0b0b0b0c0b0b0b0d0a0c0a0a0b0a090900010002020100080c0b0b0c0804;
    encBuf[645] = 256'h0406050303030203010101040307040304030304030202030202030102030102;
    encBuf[646] = 256'h050205040203030200010900000103060303030201000908000901020801010a;
    encBuf[647] = 256'h0a080d0b0a0f0d0a0c0b0a0c0a090b0c0b0e0c0b0d0a0b0a09090909090b0d0c;
    encBuf[648] = 256'h0b0c0a0b0a0a0a0b0b0c0c0a0a09000808000a0b0b0d0b000105060403030202;
    encBuf[649] = 256'h0000080808010203060403030302020208000101050603040402020101000000;
    encBuf[650] = 256'h0305050404020302020101000203040403030402010101010101010202010101;
    encBuf[651] = 256'h02050403060203010100080809080001020202030303060304020208090c0b0b;
    encBuf[652] = 256'h0a0104050402010a0c0e0b0c0a08000203030304020205040404040303030304;
    encBuf[653] = 256'h0304050402040202020101010203050404030302030202030502030402020401;
    encBuf[654] = 256'h0403030504020303020102000303050504020403010301010201010304020502;
    encBuf[655] = 256'h0204020202030001080909090b000000050208000c0e0b0d0c0a0b0a0a090b09;
    encBuf[656] = 256'h0b0c0a0c0d0a0b0d0a0c0a0b0b0a0a0b0b0b0d0d0b0c0c0b0c0b0a0a0a0b0b0c;
    encBuf[657] = 256'h0b0d0c0b0b0b0c0a0a0a0b0a0b0c0b0c0b0a0b0c0a0b0b0b0b0c0a0a0b0b0b0c;
    encBuf[658] = 256'h0c0b0b0c0b0b0a0b0b0a0b0b0a0b0b0b0d0c0b0d0b0b0a0a0000010402030200;
    encBuf[659] = 256'h0800090005030705030305020202020102010303030405030403030403010202;
    encBuf[660] = 256'h0002020104030403040203030202030204030305040204040203040202020100;
    encBuf[661] = 256'h010800010800010800000909080c0b0a0f0d0b0d0c0a0b0a0908000100090b0f;
    encBuf[662] = 256'h0e0b0b0b09080003020301080a0c0c0b0a0a08020101030000000909090d0b0c;
    encBuf[663] = 256'h0d0c0a0b09090800010808090a0a080903060204050104030405030402020100;
    encBuf[664] = 256'h00080103060503030300090c0b0c0a0102070303030208090b0b090206050404;
    encBuf[665] = 256'h0202010108080800020305040403020202020101010204030503030202010000;
    encBuf[666] = 256'h0900000205030303020000000407050404030402010100010205030603030202;
    encBuf[667] = 256'h0100080001020504030302010808090900030406030202010800080802050405;
    encBuf[668] = 256'h0402040202020202030503050304030302030108000000020403050201000a0d;
    encBuf[669] = 256'h0b0c0b080001030200090d0f0b0b0a0908000201000a0d0d0c0b0a0a08080108;
    encBuf[670] = 256'h080a0e0c0c0c0a0a0a09090a090b0d0c0b0d0b0a0b0b0a0a0b0a0c0c0b0d0b0a;
    encBuf[671] = 256'h0b0a0a09090a0c0b0c0c0b0b0b090a09080a0b0e0c0c0b0b0b0a090808080b0c;
    encBuf[672] = 256'h0d0c0b0c0a090808010100080a0c0c0b0c0908000303040301080a0c0c0a0900;
    encBuf[673] = 256'h0503050402010009090a0909010304040201080a0c0a0b090102040502010108;
    encBuf[674] = 256'h0800010407040304030203010101010304030503030203010200080808090900;
    encBuf[675] = 256'h080104010202090b0a0f0a080901040203030202030305070204030301020909;
    encBuf[676] = 256'h090b0a080800010a0c0d0e0b0c0c0b0b0e0b0c0b0b0b0a090008080a0d0c0c0c;
    encBuf[677] = 256'h0b0a080103040404020100080808080003040405020302020001090800080002;
    encBuf[678] = 256'h0204030203020202040305040204010100080802030705040304030201000000;
    encBuf[679] = 256'h0002040504030402030100010002030306030303020201030206040304040202;
    encBuf[680] = 256'h0101010303050603040304020201020100020304040402030302000009080909;
    encBuf[681] = 256'h01030307040103010808090a0801010604040304020201010201020404020502;
    encBuf[682] = 256'h0203020102020103030003000b090d0e0a0a0b09090b090a0e0a0b0d0a0a0a01;
    encBuf[683] = 256'h010105030204020001080a08090a020302070200000c0f0b0d0b0b0c0a09090a;
    encBuf[684] = 256'h090a0d0b0e0c0a0c0b0a0b0a09090909090b0c0c0c0b0b0c090a090008010108;
    encBuf[685] = 256'h08080c0c0c0c0b0b0c0a0a0a0a090a0b0d0d0c0c0b0c0b0a0b0a090908090a0a;
    encBuf[686] = 256'h0c0b0c0c0a0b0a0a0a0908080800000001090c0b0e0b0b0c0908000203020001;
    encBuf[687] = 256'h0a0d0a0d0b0a0a0a0a0a0a080900040203050108090d0c090900070306030303;
    encBuf[688] = 256'h030100010900000802020303050203040000080b0e0b0e0a0908010305040302;
    encBuf[689] = 256'h02000808000801040405030303040102020201020808080b0c09090802000008;
    encBuf[690] = 256'h0f0e0b0e0b0b0c0a09090a090a0b0b0c0b090908010800010800020002050001;
    encBuf[691] = 256'h010a0900090207020304080b0f0d0b0c0a09000103040101090c0c0c0c0a0908;
    encBuf[692] = 256'h0103040503030402010201000102030605030404020302010000080000000103;
    encBuf[693] = 256'h0304030303030304030302020000080106050505030403030302010101020205;
    encBuf[694] = 256'h040403030402020302020303020303020202030504040404030303020108090b;
    encBuf[695] = 256'h0c0b0a0801060403050200000a0c0b0c0b090002050304020108090b0d0a0b0a;
    encBuf[696] = 256'h09080808000900090901080901090c0a0d0c0808010604040304010208080909;
    encBuf[697] = 256'h0b080908020202040300000a0e0b0e0c0a0c0a0b0a0b0b0b0b0c0b0c0b0c0b0b;
    encBuf[698] = 256'h0c0c0b0c0c0a0a0a090800010008080c0c0d0b0c0b0b0b090a08090a0b0d0d0c;
    encBuf[699] = 256'h0d0b0c0c0b0b0a0b0b0a0b090b0b0d0b0e0a0c0a0a0a0a09080000000008090c;
    encBuf[700] = 256'h0b0d0c0b0b0b09090800010000090c0b0f0b0a0c0a090908010801010800010a;
    encBuf[701] = 256'h0a0a0f0b0a0b0a08080206020204020103000102090002090206020605030404;
    encBuf[702] = 256'h0201020808090a08000104050304040203020101000a0a0a0c09010105060304;
    encBuf[703] = 256'h0302020109090a0b0801030704030403020202010008090a0a0c080102070503;
    encBuf[704] = 256'h030402010809090b0a0a000104060203030100080b0c0b0c0b0a0b0900080202;
    encBuf[705] = 256'h0008090f0b0b0c0a0909000809090a0b0a020606050403030200000908080206;
    encBuf[706] = 256'h050404040202010101000808000001010403050303020301080a0a0d0a090802;
    encBuf[707] = 256'h0504050402030302010200000101040404050304040202020108000000020305;
    encBuf[708] = 256'h0403030502020203020303020203010302020406020503030502010101080800;
    encBuf[709] = 256'h0901030307050304030103010808090b080808040504040302020208080a0c09;
    encBuf[710] = 256'h0a0a010202070402040200000a0c0b0c0b0a0808040203040108090b0e0a0b0b;
    encBuf[711] = 256'h0a090902010004010000090e0b0c0d0a0a0a080801010108090d0d0a0c0a0a08;
    encBuf[712] = 256'h0908080a0a0d0c0c0b0b0a0a0a090b0c0b0d0c0b0c0c0a0b0b0a0a0a09080800;
    encBuf[713] = 256'h0a0c0c0d0c0b0c0b09090001010101090a0c0e0c0b0b0c0a090908080800090a;
    encBuf[714] = 256'h0c0e0c0b0d0b0b0b0a09090908090a0b0e0c0b0c0a0b0a0a0908080808080808;
    encBuf[715] = 256'h090a0b0b0e0b0b0b0c0a090900080101000a0c0f0d0b0c0b0b0a090102020501;
    encBuf[716] = 256'h00000b0c0b0d0a09090003020305020203000102080000090005020705030305;
    encBuf[717] = 256'h02010108090a0b090800020602040302020109090a0c0a080903070304040101;
    encBuf[718] = 256'h00090a0b0d0a080801030202020808090c09090a0a080b0a0009020703050301;
    encBuf[719] = 256'h090a0f0b0c0a09010206030302010a0c0b0d0a0800020404030201080a0c0c0b;
    encBuf[720] = 256'h0b0a0001030602030108090b0e0b0a0900020504050203020100000908010103;
    encBuf[721] = 256'h0704040303030202000808080001040503050302020000080809080102040603;
    encBuf[722] = 256'h0403030302020301020404040504030303030201010101020405030402020100;
    encBuf[723] = 256'h09090908010204030202000909090a0801000303000301040704040502020101;
    encBuf[724] = 256'h0900080005040404030102080a0a0c0c0a0a0a080800000109090d0e0c0c0c0b;
    encBuf[725] = 256'h0a0a000003040201000c0d0c0c0b0a090802010302000a0c0d0c0b0c0a090808;
    encBuf[726] = 256'h0008000009090c0c0c0b0c0a0b0909080800080a0b0d0c0c0b0a0a0908080909;
    encBuf[727] = 256'h0b0d0c0b0c0b0b0a0b090a0b0b0d0d0b0c0c0b0c0b0a0a0900010001080b0d0e;
    encBuf[728] = 256'h0c0a0b0a09000102030202090c0b0f0c0a0b0a0a08000102030400080b0f0c0b;
    encBuf[729] = 256'h0d0a0909000101020308090a0e0b0b0c0a08090102030305020102090a0c0c0b;
    encBuf[730] = 256'h0a09000303050301090a0f0b0a0b0801000203080a0b0f0a0800020702030201;
    encBuf[731] = 256'h08090b0900010604040303020202010304020303010203020506040305020201;
    encBuf[732] = 256'h0009090a08010205050203030302020002020102030306050404040303030100;
    encBuf[733] = 256'h090b0a08000505040402010108090a0808020404040303020201010102030304;
    encBuf[734] = 256'h0403030403050302020200080808020505040403030100090809000305050502;
    encBuf[735] = 256'h0302020101000202020503030503030404020303020301000101010405030503;
    encBuf[736] = 256'h0202010800000a00080901010006030404030202000a080a0b01040507030203;
    encBuf[737] = 256'h020000080a08080903010002000a020208070009090d0e0a0b0a080008040009;
    encBuf[738] = 256'h080c0d0a0b0b08080901090d090a0c000100040108080b0f0a09090201000309;
    encBuf[739] = 256'h0e0b0d0c09090900000a0a0d0e0a0b0a090808000009090b0e0a090a00080802;
    encBuf[740] = 256'h080a00000007040204000a0a0e0b0a090003050202000c0b0e0c090a08080108;
    encBuf[741] = 256'h000a0b0c0c0b09080900090c0c0c0c0a0a0900000000090b0c0d0c0b0b0b0a0c;
    encBuf[742] = 256'h0b0c0b0c0a0b0a0a0c0b0c0e0b0c0b0b0a0a09090808090b0b0d0c0a0b0c0b0b;
    encBuf[743] = 256'h0c0c0a0b0a090900090a0d0d0d0c0b0c0a0a09080008080a0b0c0d0b0c0b0b0a;
    encBuf[744] = 256'h0a0a090909000809080a0b0b0d0c0a0909010203060203020008080a0c0a0c0b;
    encBuf[745] = 256'h0b0b0b080800050100000e0c0b0e0a090a080101020300010209080108010508;
    encBuf[746] = 256'h01020a01050106040203030000080b09080b08020a08000d0902000407010201;
    encBuf[747] = 256'h090b0b0e09010307070304030302020201020203050304050204020203010008;
    encBuf[748] = 256'h090b0a090a000202040201090c0e0b0c0b0a08080202030101090a0b0c090800;
    encBuf[749] = 256'h0307030403040302020100090908000407040305020100090b0d0b0a08000405;
    encBuf[750] = 256'h030403020101080800000205040404030402030203010008090a090a08010205;
    encBuf[751] = 256'h04020200090c0c0d0b0b0a090000020203030402010100080808000405060403;
    encBuf[752] = 256'h04040202020102010001010808090a0b0a090003040402090d0e0d0c0b0b0a09;
    encBuf[753] = 256'h000103040202020008090a0b0b0c0a090002060403040200090d0d0c0b0c0b0a;
    encBuf[754] = 256'h09000000010108090b0d0c0b0c0a0a0908020305030403020000090908000204;
    encBuf[755] = 256'h06030502020101010808080a0a0b0d0d0b0c0c0a0b0a0b0a0c0c0b0c0b0b0c0a;
    encBuf[756] = 256'h0b0a0a0b0a090801030404040201000a0a0b0b0901060505030303010108090b;
    encBuf[757] = 256'h0b0b0b090002050503040201080b0e0c0b0b0a0801030404030100090b0b0b0b;
    encBuf[758] = 256'h090001020300080a0f0b0c0d0b0b0d0b0b0c0b0b0a0b0a0c0b0c0b0c0a090800;
    encBuf[759] = 256'h0203040101000a08080105050504040303030303030202000008000003060504;
    encBuf[760] = 256'h04030200090b0f0b0b0b0a0001030503020208090c0c0b0c0909010204040402;
    encBuf[761] = 256'h03020000090a0a0b0900010306030402030202000008090c0b0d0b0908020605;
    encBuf[762] = 256'h0403030202080a0a0b0a00030705040303030302010100000000000102030306;
    encBuf[763] = 256'h0303040202000a0b0d0c0c0a0b090800040404040303020100090a0a08010407;
    encBuf[764] = 256'h050403040203010008080a0909080104050305020200080a0c0d0a0b0a090801;
    encBuf[765] = 256'h02030101080b0d0c0c0a0a0901010203040101010801000002020101080b0b0e;
    encBuf[766] = 256'h0c09090901030204020a0b0f0e0b0b0c09090002030404020200080b0a0d0b09;
    encBuf[767] = 256'h08080305040403030300080a0d0d0b0c0b090908010001000a0d0d0d0b0c0a0b;
    encBuf[768] = 256'h090900000100010009080a0b090a09020202060201020102030203040109090e;
    encBuf[769] = 256'h0e0b0d0b0b0a0a08000001080b0e0d0c0c0b0b0a0a090800020202010208080b;
    encBuf[770] = 256'h0c0c0b0b0b080003070403040101090b0f0b0d0b0a0b09080001010108090e0c;
    encBuf[771] = 256'h0c0b0c0a0a0900010103030200080a0c0c0b0b0a09000102020301080a0e0d0c;
    encBuf[772] = 256'h0b0b0d0a0a0a0a0a0b0b0c0c0b0c0b090a0a09090a0b0c0c0a0a090004040604;
    encBuf[773] = 256'h0303030201010809080800030704040303030201090a0c0c0b0a090002040503;
    encBuf[774] = 256'h040101080a0b0e0b0b0b0a00010405030302000a0b0f0b0c0a0a080002040203;
    encBuf[775] = 256'h02000a0c0c0d0a0b0909000203050303020000090a0a0a000204060403030302;
    encBuf[776] = 256'h01010808080808010800000a0a080a09030102030e0d0d0f0b0b0d0b0a0a0800;
    encBuf[777] = 256'h00010208090c0e0c0b0d0a090900010302030200080b0d0b0b0b090802050403;
    encBuf[778] = 256'h05030203010100090a090a0003060605030304010100090a0a0a090801040503;
    encBuf[779] = 256'h030501010008090a0a0b0909010204060304040202020000090b0b0c0a090005;
    encBuf[780] = 256'h05040502020208090c0c0b0a0a000205050303030200090b0b0d0a0908020306;
    encBuf[781] = 256'h040303030200080a0b0e0a0a090802040404020200090b0d0c0c0b0a0a090001;
    encBuf[782] = 256'h02020202080a0d0c0c0c0a09090002030404030202010008090a0b0a09000206;
    encBuf[783] = 256'h05040403030200090b0d0c0a0a09000203040202080b0d0d0b0b0a0a08000101;
    encBuf[784] = 256'h010108080a0b0a09090000090a0d0d0d0b0c0a08000203050202090b0f0c0b0b;
    encBuf[785] = 256'h0a08010306030402020008090909090001020404040404030304020100090b0c;
    encBuf[786] = 256'h0c0b0908010306030201080b0f0b0d0b0a0b090800010203020100090c0c0c0b;
    encBuf[787] = 256'h0b0b0900030405040302020100090b0c0c0b0a09010306040403020200090b0c;
    encBuf[788] = 256'h0b0b0a08010405040303020200000a0a0c0b0b0b0a0003060504030301000a0c;
    encBuf[789] = 256'h0d0c0b0b0a09000103030301080b0d0d0c0b0b0a080801030306020303010101;
    encBuf[790] = 256'h0809090a0900000307050404030402020100090c0b0b0a090104060305020200;
    encBuf[791] = 256'h090a0d0b0c0b0a090001030305020200090b0d0c0b0b0a090003050403030201;
    encBuf[792] = 256'h090a0c0c0b0c0909000204040403020201000a0b0d0b0a090002050503030301;
    encBuf[793] = 256'h00090b0d0b0b0a0800020404040303020100090b0c0c0b0a0a08020306030302;
    encBuf[794] = 256'h00090c0c0d0a0b0a09080102040403020101090a0c0c0b0a0908020403040202;
    encBuf[795] = 256'h010009080808080009000808030505060303040100090b0d0b0c0b0908090100;
    encBuf[796] = 256'h01010201010108090c0f0c0b0b0b0900040503040301010a0c0d0c0b0b0a0a08;
    encBuf[797] = 256'h00020404020301090a0e0c0b0b0b090002050304020200080a0b0d0c0b0a0a08;
    encBuf[798] = 256'h0002050404020300080a0d0c0b0b0a08000203030300090c0d0c0b0c0a0b090a;
    encBuf[799] = 256'h09090002030405030202000a0b0c0c0b09000306040304030200090a0c0d0b0b;
    encBuf[800] = 256'h0a08000204030302080b0e0c0c0b0c090a09080808080808000800080a0d0c0d;
    encBuf[801] = 256'h0b0b090801040504020201080b0b0d0b0a09000204040302030100080a0a0a0a;
    encBuf[802] = 256'h0908020405040303030302000008090a0c0b0b0b0908030706030302000a0d0d;
    encBuf[803] = 256'h0c0b0b09090102030201080b0e0c0a0a09080102030202020001000000000000;
    encBuf[804] = 256'h0001000002040101010000010107050305030101080a0a0b0b08000304040100;
    encBuf[805] = 256'h000b0b090a09080a080a0c0a00020507030302010a0d0d0c0c0b0b0b0b0a090a;
    encBuf[806] = 256'h08080908090b0e0d0c0c0b0b0900020405020200080b0d0c0a0a090001030403;
    encBuf[807] = 256'h0201010808000101030403040303040202030201020008090c0e0c0d0c0b0b0a;
    encBuf[808] = 256'h090001040302020a0c0e0c0b0a0a00020404030201000b0c0c0b0b0909010203;
    encBuf[809] = 256'h05030304030202010008000800030405040201010a0d0b0e0c0a0c0a090a0808;
    encBuf[810] = 256'h0801010000080a0c0b0d0a090802040303020a0d0e0c0b0a0b08010104030202;
    encBuf[811] = 256'h00080a090a010304060402020208090b0d0c0a0b0b090b0908090a00090a0101;
    encBuf[812] = 256'h04060304020109090d0b0a0a0004030304080a0f0e0b0b0b0a00020504030402;
    encBuf[813] = 256'h0108090b0b0b0a080304050403020100090a0d0b0a0a08020404050203030100;
    encBuf[814] = 256'h0808090809000202040502020302020202020302020303070403050403040303;
    encBuf[815] = 256'h04010101000a090909090800030403040201090b0f0c0b0c0b09000203060303;
    encBuf[816] = 256'h030201080a0b0a0a000306060404020303010100080900000105030603030303;
    encBuf[817] = 256'h0100080a0a0b09080101040302020108090b0b09000007030205020102000801;
    encBuf[818] = 256'h0800030604050302030109090b0b08020407050304020100080a0a0b0a080003;
    encBuf[819] = 256'h050402030200080a0d0a0a0a08030307040203020001080b09090a0001010301;
    encBuf[820] = 256'h0801080b05040406030303030008090b09000007040305020101090c0c0b0c0a;
    encBuf[821] = 256'h090803040405020201000a0a0c0c090a0801020205010009090d0b0c0b090909;
    encBuf[822] = 256'h01020305040203030000080a0b0b0b09000206030302010b0b0d0d0a0a0a0802;
    encBuf[823] = 256'h0103030103030900080a08000c0a0d0e0a0c0d0a0a0b08010004030201080c0b;
    encBuf[824] = 256'h0e0b090800050403030200090c0d0b0b0b090801020208080b0c0c0b0b080002;
    encBuf[825] = 256'h0404020300080a0b0d0808010405030302090b0f0d0b0b0b0a00030504040201;
    encBuf[826] = 256'h08090b0d0b0b0b08010304040301000b0c0e0c0b0a0b08000103050302010009;
    encBuf[827] = 256'h0b0d0b0a0900010305020101090a0b0d0b0c0a0a0a090a080801000203060202;
    encBuf[828] = 256'h00090d0c0c0b0c0a09080800020000090b0f0d0c0a0b0a08080101030201080a;
    encBuf[829] = 256'h0d0d0c0b0a0b0a0a0a09090b0a090a0b0a0b0d0d0b0c0b0a0900010404030201;
    encBuf[830] = 256'h08090b0d0b0b0a090808000008090a0b080a0a090a0d0b0d0b0b0c0b08080800;
    encBuf[831] = 256'h0108090c0d0c0c0d0b0a0b090000010301010a0e0c0c0b0b0a0801020102000a;
    encBuf[832] = 256'h0b0f0c0a09090101020400080a0b0e0b0b0901020504020202090c0c0c0b0a0b;
    encBuf[833] = 256'h09020204040200090d0c0c0c0a0a090801010202080a0b0f0b0c0b0a08090001;
    encBuf[834] = 256'h0008010909090b0b090909000000010b0a090c0b0a0c0a090a0a010a0b080d0b;
    encBuf[835] = 256'h0a0c0a01000205020203080b090f0a0b0c0a080b0a090a09010908010b0b0b0f;
    encBuf[836] = 256'h0b080a090002050502020308080a0d0b0b0b0900080205020404000102080800;
    encBuf[837] = 256'h0900020106050204030202000808090b0b090a08030204070203040302030202;
    encBuf[838] = 256'h0200090201030703040503020108080a0d0c0a0a0a0800020504030302020009;
    encBuf[839] = 256'h0c0b0b0b00030607030304020108090a0b0b0908010505040304020202000808;
    encBuf[840] = 256'h090000020504040303020100090a0a0a0a080104040303030303020405040402;
    encBuf[841] = 256'h030301000009090808020403030301080c0d0d0a0a0900020604040402020201;
    encBuf[842] = 256'h08080808000104040402020100080a0908010604050303040201000808010000;
    encBuf[843] = 256'h030503030201080c0d0b0c0c0909000104050303020208090a0b0b0802040604;
    encBuf[844] = 256'h03020108090b0d0a0b0a08080002020202000000080802030106010100090b09;
    encBuf[845] = 256'h0d0b000205060403040100090b0c0a09000406040403020200090a0b0d090908;
    encBuf[846] = 256'h02030404030100080a0b0d0b0a090902040403040301000909090b0b09090008;
    encBuf[847] = 256'h09090a0d0a0b0b08090a00090f0b0d0c0a0a090203060403020200090a0d0d0a;
    encBuf[848] = 256'h0a09000104040403030100090c0b0c0b0901020504030302000a0c0c0d0a0b09;
    encBuf[849] = 256'h090800020102010100090b0e0b0b0d090908000103030201000a0d0d0c0b0c0a;
    encBuf[850] = 256'h09080801030403040200000b0d0c0b0a0a08000203040200090a0d0c0a0a0900;
    encBuf[851] = 256'h010204010102010800080a000a0b0b0e0b0a0c0a080900010008020201010000;
    encBuf[852] = 256'h000c0a0b0e0a0b090a090a0a0c0d0c0a0d0a0a0a090a080908090a0900020101;
    encBuf[853] = 256'h0801080b0b0c0d0c0a0b090b09080802040404040201080b0e0c0b0b09010405;
    encBuf[854] = 256'h040202000a0c0d0c0c0a0a0900020303040300090b0e0b0c0b0a080002030503;
    encBuf[855] = 256'h0200090c0c0c0b0b0a09080102020201010808090a0a0b0c0b0b0c0a08020604;
    encBuf[856] = 256'h04040201080a0d0d0b0b0b0b080102040404020200090c0d0b0b0a0908020403;
    encBuf[857] = 256'h040201080b0e0c0b0b0a09000103040303030202010008090a090b0b08010106;
    encBuf[858] = 256'h03030200090d0f0c0b0b0c0b0a080003050403030301080a0d0d0a0b09080103;
    encBuf[859] = 256'h05030301000a0c0c0b09090104040404020201000009090a0909090008000808;
    encBuf[860] = 256'h0a0a0d0a0a0a01020307040202010808080a00040405030301000a0c0d0b0a0a;
    encBuf[861] = 256'h0a0808080101000203020402010201090b0a0c0a090803060304030000000a0a;
    encBuf[862] = 256'h090d0b0b0b00010207070303030201090b0c0b0d09090001040403040101000a;
    encBuf[863] = 256'h0b0e0b0c0a0a080205040403030208090c0c0b0b0a0001030603020101090a0c;
    encBuf[864] = 256'h0c0b0b090900010204040202030108000b0d0b0c0b0a08000104040403040202;
    encBuf[865] = 256'h00090c0d0b0b0a0802070403040201000a0b0c0c0b090802030503040100080a;
    encBuf[866] = 256'h0b0b0c0a090801020304030201080a0d0b0c0a09090102030302020100010202;
    encBuf[867] = 256'h030301080c0d0c0b0c090802040404020008090b0c0a09000101030201030301;
    encBuf[868] = 256'h01080a0c0e0b0b0b0909010305030202020009000204030303010c0e0c0c0b0a;
    encBuf[869] = 256'h080003030401080a0d0d0b0b0a09080103050404020201080b0d0c0c0a0a0a00;
    encBuf[870] = 256'h000303040201090c0c0b0c0a090800010001010202030403080a0f0e0b0c0b0a;
    encBuf[871] = 256'h090002050303030201090b0d0b0c0a09000105030504020201080a0d0c0c0a0a;
    encBuf[872] = 256'h080102040402010109090b0c0b0a0a080103050403030201090b0e0b0c0a0a08;
    encBuf[873] = 256'h0001050203010008090a09080003040301000a080808040403050201090c0c0c;
    encBuf[874] = 256'h0b0b00010405050304020101000809090a0a0801040504030202090a0c0d0a09;
    encBuf[875] = 256'h0801040304020201080000000103020201090d0c0b0c0908030403030208090c;
    encBuf[876] = 256'h0c0a0a010205040303030201010a0b0b0e0c0a0800020304040108080a0a0004;
    encBuf[877] = 256'h04060402010109090b0c09010305040302000a0c0d0c09090001020304030000;
    encBuf[878] = 256'h000a090b0c0b090a00030306040201080a0b0d0c090a08010303030301090d0b;
    encBuf[879] = 256'h0a080205040101000a0a0a0a01010305030103010908090b0a0c0d0a0a090101;
    encBuf[880] = 256'h0505040202080a0c0d0c0a090800020404010108090b0a0b0c09090901020205;
    encBuf[881] = 256'h0502030100080b0d0c0b0b0a000103040202010a0c0a0c0b090b0b0a0b0c0909;
    encBuf[882] = 256'h080103050108090c0f0c0a0b0b080000030304020100090c0c0c0b0c0b090908;
    encBuf[883] = 256'h0304040201080a0e0d0a0b0908010305020201080a0b0c0a0a09010100010008;
    encBuf[884] = 256'h0d0b0a090a08030306030100080a0c0c0c0a08080102030400090e0d0d0b0b0a;
    encBuf[885] = 256'h08000404030302080a0c0c0a0b08000303050200090c0c0a0c0a080001020203;
    encBuf[886] = 256'h010008090909080801060203040200080c0d0c09090901030404020100090b0c;
    encBuf[887] = 256'h0b080802050502030108080b0d0b0a0b0a080901000002010a090a0a0b0b0908;
    encBuf[888] = 256'h08030403030301090b0c0a090a0803040302000a0b0b0e0b0a00010305040303;
    encBuf[889] = 256'h0101090a0b0d0b0a0001050503030301090b0f0c0a0a09000203050402020009;
    encBuf[890] = 256'h090a0b0a0801030403030109090b0b0b0a0a0000000001080a080b0901030406;
    encBuf[891] = 256'h03040302080a0c0d0c0a0a0900020404020200090c0c0b0b0b08020603050302;
    encBuf[892] = 256'h0101090b0c0c0a0a0900010304030201000a0a0d0b0a09090204030404000008;
    encBuf[893] = 256'h090c0a0b0c0b0a090909080909080100000908080b0b0a0a090a0909080a0a09;
    encBuf[894] = 256'h0c0c0b0b0c0a0b0908090a01000a0a0908080000020002020009090b0c0b0c0a;
    encBuf[895] = 256'h090801030202020a0a090d0b0a0a09000101080100090b0c0a0b0c0a08090b0a;
    encBuf[896] = 256'h09090a090108000102000808080a0d0a090a09010204040101000a0c0b0c0a0a;
    encBuf[897] = 256'h0a08020204030403020908090a0b0a0b0001000305030402020201090a0b0b0b;
    encBuf[898] = 256'h0b09030703030503020009090a0b0c090802050303050100080b0c0b0b090003;
    encBuf[899] = 256'h06040303020008090b0a0808050503030301000a0c0c0b0a0002040603040201;
    encBuf[900] = 256'h00080a0a080801040405040201010009090a0b08000003060303030201030203;
    encBuf[901] = 256'h030504010202080908090b000202040404020009090b0e0a0a08030604050302;
    encBuf[902] = 256'h020108090c0a0b0a08000404040303020009090b0d0a09000205040403040101;
    encBuf[903] = 256'h0009090a0a0b080001030703030402010009080a0b0801020704030403010100;
    encBuf[904] = 256'h0a0a0a0b0a080005030405020001090909090a010203070302020100080a0a09;
    encBuf[905] = 256'h090103020306010001080a08090b01020003030103020902000a010008010008;
    encBuf[906] = 256'h02010902010804010802020a08090d00080a02010105020103000b00090e0909;
    encBuf[907] = 256'h09080000040101030008090c0c0a0c0b090a0a010303040201020a0d0b0f0b0b;
    encBuf[908] = 256'h0a0a00010207020101080c0b0c0c0b0a09010203060201010a0b0c0d0b0b0909;
    encBuf[909] = 256'h020204030208000a0f0b0b0b0a090801010202000b0c0e0b0b0b0b0908000100;
    encBuf[910] = 256'h00000a0c0b0c0b0a0b0a090b0b0c0d0b0b0d0b0a0a0a09090a0b0c0a0b0c0d0a;
    encBuf[911] = 256'h090a090a090c0d0b0b0d0c0a0b0a0808090a0a0a0c0d0a0c0a09000101020202;
    encBuf[912] = 256'h080b0e0c0c0b0a0b0a09000108000a0b0d0c0c0a0b0a0900080103000901090c;
    encBuf[913] = 256'h0c0c0b0b0d0b0b0b0c0b0a09090908000a0a0b0c0b0c0c0b0a08000103010200;
    encBuf[914] = 256'h0a0b0e0d0a0b0b0a0908020202040100000b0b0b0b0a080a0003010103090101;
    encBuf[915] = 256'h090d090b0c090c0a080908020802040100080b0b0b0c0a090002050203030009;
    encBuf[916] = 256'h090c0d0b0a0900080106010801090b0c0a0c0809020401030309090a0d0b0b0b;
    encBuf[917] = 256'h08010002030000080c0b0a0b0b080103050304020101080900000a0002000100;
    encBuf[918] = 256'h0901010908010a08020908000900000802050203040102000b0b0a0e0a080901;
    encBuf[919] = 256'h030205020800090f0a090a0001020504030201080a0a0c0b0900020603030303;
    encBuf[920] = 256'h00080b0d090a0803050504020201080a0a0b0a000003070304030100080a0b0a;
    encBuf[921] = 256'h0a080304070303010209090a0b0b000005040404020101010809090003040405;
    encBuf[922] = 256'h02020200090b0b0b08010204060202030109090a0a090002070403030300080a;
    encBuf[923] = 256'h0d0b0a0b08000306040203010000090a09080307030603020302000809090b09;
    encBuf[924] = 256'h0002020603040202010009080901050304040403010108080a0b0a0a01000303;
    encBuf[925] = 256'h0201000b0c0b0b0b08040504030503010208090a0a0a0002040504040201080a;
    encBuf[926] = 256'h0a0c0a0a000206040403030200080a0a0a0a0003060503030201080a0c0b0a0a;
    encBuf[927] = 256'h08040404040302010009090b09010106050304020201080a090a0a0002040603;
    encBuf[928] = 256'h03030200000a0b09010206050403040102000808090a00010105040203020001;
    encBuf[929] = 256'h0809000108050503050303040302020201030303060201030401020202030302;
    encBuf[930] = 256'h0503000404010404020304020401010200080100000201010701080101080001;
    encBuf[931] = 256'h0806040206030204030101020001020004040204030103020801080803050206;
    encBuf[932] = 256'h040205020002010801000902030105020103010a010a0e000009050301060200;
    encBuf[933] = 256'h020009000009030402060301030109080a0e00080805030305020001090c090a;
    encBuf[934] = 256'h0c08010005020103020d0a0b0e0a0a0a01010004030801090e0a0c0b0a090902;
    encBuf[935] = 256'h030105010a080a0e0a090b00010004020101090d0a0c0d090909000008010a0e;
    encBuf[936] = 256'h0a0c0c0a0a0a00000802080a0a0e0e0a0c0b090908000108000b0d0c0d0b0b0b;
    encBuf[937] = 256'h09080101030300080c0f0b0c0b0a0a0801020201000c0c0d0d0b0b0a09080002;
    encBuf[938] = 256'h0201000a0e0c0c0b0c0a080800000100090b0d0d0b0c0b0a090800000100090a;
    encBuf[939] = 256'h0d0c0c0b0a0a0a08000808080a0c0d0c0c0a0b0b090a09090a0a0c0d0c0b0b0b;
    encBuf[940] = 256'h0b0b0b090b0b0b0e0c0b0d0b0a0a0b090a090a0b0d0b0e0b0b0b0c090a080809;
    encBuf[941] = 256'h09080c0c0b0d0b0b0a0a090908000a0b0c0f0b0c0b0c0a0a0a08090a080b0c0a;
    encBuf[942] = 256'h0e0b0a0b0b090b0a090a0a0a0f0b0a0c0c0a0b0b0a0c0a090c0a090a0b080b0a;
    encBuf[943] = 256'h080c0b090e0a090c0a000b09080b0c0a0f0b0a0d0b090a09000900030a0a080f;
    encBuf[944] = 256'h0b090d0a080908020800010b0e090f0a090b09080801030000030b0b0a0f0b08;
    encBuf[945] = 256'h0b08040002050808000d0b090d0a080a00020102030809000f0b080b09020802;
    encBuf[946] = 256'h060001020b0b090e0a080a08040003050800020a0a010a000501030701010208;
    encBuf[947] = 256'h08000a08030803070302050000010a08010902070102050101020808010a0004;
    encBuf[948] = 256'h0004050203040001020900020902050304050202040001010000030105040303;
    encBuf[949] = 256'h0502020301010300010402040502030402020301020301040402040502030303;
    encBuf[950] = 256'h0304010203020305020404010304020303020403020403030503020403020403;
    encBuf[951] = 256'h0203040203030303040305030304030403030303030304030403050304030303;
    encBuf[952] = 256'h0402020202030205040304030403030302030203030305050204040203020302;
    encBuf[953] = 256'h0201030202050403050402020301020208020102040404040303030301020108;
    encBuf[954] = 256'h0204020604020403020301000000080303030705020302010201080101000503;
    encBuf[955] = 256'h0405030203020001080902010106040204030202020901000903040207030204;
    encBuf[956] = 256'h020101010900000a03030207040103020001000b010809050302070301030209;
    encBuf[957] = 256'h00090c08080a05020205030002080b090c0c000008050301050109010a0d0909;
    encBuf[958] = 256'h0b00010004020002000e080b0d08090901010804010a000a0e090a0c00090902;
    encBuf[959] = 256'h080a010a0e090a0e08090b00090b010a0d080a0d09090c08090b080a0d080a0d;
    encBuf[960] = 256'h09090c08090c08090c080b0b090b0d08090b080a0e080b0c090a0c08090b0809;
    encBuf[961] = 256'h0c090c0d0a0a0d09090a000909000a0c0b0c0d0a0b0c080909000009090b0f0b;
    encBuf[962] = 256'h0c0c0a0a0b0808000108090a0d0d0c0b0b0b0a0900000002090b0e0d0c0b0c0a;
    encBuf[963] = 256'h090908000000000a0c0c0c0d0a0a0a090008010008090c0d0b0c0c0a0a0a0808;
    encBuf[964] = 256'h000000090a0d0c0c0b0c0a090a08000000080a0b0e0c0c0b0b0a0a0900000000;
    encBuf[965] = 256'h090b0e0c0c0c0a0b0a090800000108090c0d0c0b0c0b0a0908000000010a0b0e;
    encBuf[966] = 256'h0d0b0b0c0a090808010000080c0b0d0c0b0a0b0a08080000080a0b0e0d0a0c0a;
    encBuf[967] = 256'h0a0a09080809080a0c0a0d0b0a0c0b080b09080b0b0a0f0b0a0c0a0a0b0b090b;
    encBuf[968] = 256'h0b0a0e0b090d0a090c09080a09080b0b0b0f0b0a0c0b090a0a000b09000d0b0a;
    encBuf[969] = 256'h0e0b0a0c0a000a00020908000d0b0b0f0b090b09010900040908000d0b0a0e0a;
    encBuf[970] = 256'h08090802080102090a080f0a090b0a000900040800020c0a000d09010a08040a;
    encBuf[971] = 256'h08030c0a010d09020901070000030909000d09000902060102050000010b0b08;
    encBuf[972] = 256'h0e09010003070103030000010b0a090b00040206050201030808080c0a080900;
    encBuf[973] = 256'h050204050102020000080a08010802060204030201020908010b080301040702;
    encBuf[974] = 256'h0205010203000203000304010104000204000305020304010302000203000307;
    encBuf[975] = 256'h0305040303040102010808010802040306040202030201010000020205050304;
    encBuf[976] = 256'h0402020201010100010203050402040302020201030204040403050203020101;
    encBuf[977] = 256'h01010103050306030304020100000808010205050404030202010009090a0900;
    encBuf[978] = 256'h030704040402020000090a0a0908010505040402020108090a0b0b0900020605;
    encBuf[979] = 256'h0304020101090a0a0b0a080105050403030200080a0c0a0b0a00030505040202;
    encBuf[980] = 256'h0100080a0b0b09090205040503010200080a0a0c0a080803050305030102000a;
    encBuf[981] = 256'h090a0a09000205050204010101090a090a0900010307030203020000080a0808;
    encBuf[982] = 256'h0804030306020102080908090a02020207040003010900090b01000907020103;
    encBuf[983] = 256'h0208000a0f080a0a020101070201020109080a0d090a0a01010006020002080c;
    encBuf[984] = 256'h080b0e09080901020206020102000b090c0d0a090b00010804010002080d090b;
    encBuf[985] = 256'h0e08090902030106020001080c0a0b0f09090a08000802020801090c0a0c0c09;
    encBuf[986] = 256'h090a02020206020000090e0a0d0b0b0a0b000008030208010a0f0a0b0e090909;
    encBuf[987] = 256'h010101040108080b0f0b0c0c090a0a000100020108000c0d0b0c0b0b09090102;
    encBuf[988] = 256'h0203020a0b0f0f0a0b0c09090901010101010a0a0e0c0b0c0a09090002020102;
    encBuf[989] = 256'h080c0c0d0c0b0b0a090801020101010a0d0d0c0b0b0b09080001030108090c0e;
    encBuf[990] = 256'h0b0d0b0a09090000000100090b0d0d0b0b0c0a090908080008090b0c0c0c0b0b;
    encBuf[991] = 256'h0c0a0a0908090a090c0b0d0b0c0c0a0b0b0b0a0b0b0a0b0c0b0c0c0b0b0c0a0b;
    encBuf[992] = 256'h0c0a0b0b0b0d0b0b0d0b0b0c0b0b0b0c0a0b0b0b0d0b0a0b0c0a0a0b0a0c0b0b;
    encBuf[993] = 256'h0c0c0b0d0b0a0c0b090b0b090b0b0a0d0b0a0d0b0b0c0a090b09080a09090d0c;
    encBuf[994] = 256'h0a0e0b0a0c0b090909000800010b0b0b0f0d0a0a0b080900020000020a0d0a0f;
    encBuf[995] = 256'h0b0b0b0a08080004020103090b0a0f0d090b09000801030102030a0c0a0f0a0a;
    encBuf[996] = 256'h0a0a0100030501020309090a0f0b090b09010802040102030a0a090f0a090a08;
    encBuf[997] = 256'h030003070101020a08080c0a080b080208010608010309000309010600010408;
    encBuf[998] = 256'h01030901050002070002020800020b09000a02070205050202030001010a0901;
    encBuf[999] = 256'h0902060205040203020108000a0a010a01070304060202020100010a09000901;
    encBuf[1000] = 256'h040306040303030001000b09090a010504040503030301000009090809000602;
    encBuf[1001] = 256'h0504020303010000090909080104040504020304000101080800080104030504;
    encBuf[1002] = 256'h0203030201010900000802050305040303030302020001020304050305030203;
    encBuf[1003] = 256'h0302020202030403060203040202020302040305030403040202020101010103;
    encBuf[1004] = 256'h0503060303040202010100000001030604040304020202000008000800030504;
    encBuf[1005] = 256'h0404030302010100090908080205040503040202010000090909080205030603;
    encBuf[1006] = 256'h0304020000080a08090902030406040202020100000908080802050305040203;
    encBuf[1007] = 256'h0200010009080009020303070501030201020108020101030501050301040200;
    encBuf[1008] = 256'h03010003020104030004020005020106030204040003010801080b0102000704;
    encBuf[1009] = 256'h0105020002000a08090b01020107050204020000000a090a0a00010107030204;
    encBuf[1010] = 256'h020001080a080a0a01030107040104010001080908090b010009050201050300;
    encBuf[1011] = 256'h03020a03080d01090b01010a07010004010902080d080a0c08080a0303000703;
    encBuf[1012] = 256'h0002000b080b0f0a090c00000804020003010a080c0f090a0b00000805020104;
    encBuf[1013] = 256'h0109090b0f0a0a0b090800030303050109080c0e090b0b08080803030104000a;
    encBuf[1014] = 256'h0a0e0d0a0b0c09080801010003000b090d0d0a0c0b09090a00000900080c090c;
    encBuf[1015] = 256'h0d0a0b0d090a0a08090a08090b090b0f090c0b0b0c0c0a0a0b09090a08090c09;
    encBuf[1016] = 256'h0b0d0b0d0c0a0b0b090a0a08090b0a0d0d0a0d0b0b0c0a0a0a09080909080a0d;
    encBuf[1017] = 256'h0a0d0c0a0c0b0a0b0a090a09080a0b0c0d0c0c0b0c0a0b0a0908080008080a0c;
    encBuf[1018] = 256'h0e0c0c0b0b0b0b0a0908000808090d0c0c0c0c0a0b0a090800000008090c0b0f;
    encBuf[1019] = 256'h0c0a0b0b0b090908000800090b0c0e0c0b0b0c0a0909080008010a0a0c0e0b0c;
    encBuf[1020] = 256'h0c0a0a0a090008000009090b0e0b0c0c0a0a0a09000908000a0b0b0f0c0a0b0b;
    encBuf[1021] = 256'h090b09080909080b0b0b0f0b0a0d0a090b0a090c0a090c0a090c0a090b0b090d;
    encBuf[1022] = 256'h0b0a0d0a090b0b000b09010c0a090f0b0a0d0a090a09000800020908080f0b09;
    encBuf[1023] = 256'h0d0a090a08020800040908000e0b090d0a090a08020802040900010d0b090e0a;
    encBuf[1024] = 256'h080a09020908040808020b0a010f0a000c09010900040802040800020c0a080e;
    encBuf[1025] = 256'h09000a01040103060101020909000d09000901060103050102010809000c0900;
    encBuf[1026] = 256'h0802060204040102020808000a09010802070203060101020900000a08010804;
    encBuf[1027] = 256'h0502040401020200000009000200040602030501020300010201020403040602;
    encBuf[1028] = 256'h0204010203010103020306020303030404010303020403030404020303020304;
    encBuf[1029] = 256'h0103040303050203030302040102030305040304030402030102020103030306;
    encBuf[1030] = 256'h0403030403030202020302040404030503040203020201020102040305040303;
    encBuf[1031] = 256'h0303030202020303060304040303030302010201020403050403030402010200;
    encBuf[1032] = 256'h0001010306030503030402000200080202010604030403030303010202010404;
    encBuf[1033] = 256'h0306030304040103020102020203040305030205020203030103030203040103;
    encBuf[1034] = 256'h040004030103030103030903010b02010c04020806020802010b000a0f08090b;
    encBuf[1035] = 256'h01020a06020803020a01090e01080a04040105030204020801000a0101090703;
    encBuf[1036] = 256'h0106030003020801000a01010807030105020803000b08090d08080a03020005;
    encBuf[1037] = 256'h010a010a0f080a0c00080a03010803080b080b0f090a0a02020007030003000a;
    encBuf[1038] = 256'h01080c02020207050204020102000900000a04030207040103010000090b090a;
    encBuf[1039] = 256'h0b02020107020001090e0a0d0b0b0b0b090909000a0c0b0e0d0b0b0d0a0a0b08;
    encBuf[1040] = 256'h0a0a080a0c0a0c0c0a0c0b090a0a09090908090b080b0d090b0c080a0a000009;
    encBuf[1041] = 256'h03010804000901090c080a0c010808050201040009080c0e0a0c0c090b0a090a;
    encBuf[1042] = 256'h0b090b0f0a0b0e0a0c0a0b0a0c090a0b0a0a0c0a0c0c0a0b0c0a0b0c090a0a09;
    encBuf[1043] = 256'h0a09090a0a0a0b0d0a0b0c090a08000001020101010a0c0b0e0c0a0a0a090800;
    encBuf[1044] = 256'h0009090a0e0e0c0c0b0d0b0b0b0b0b0c0b0c0b0d0c0b0c0b0d0b0a0b0c0a0a0b;
    encBuf[1045] = 256'h0a0c0b0b0b0e0a0b0c0a0b0a0b0a0a0a0a0b0a0c0b0b0d0b0a0b0a0909080100;
    encBuf[1046] = 256'h01030000000b0b080c0904010506020303020101090b090c0a080a0003090002;
    encBuf[1047] = 256'h0e0c0b0f0c0a0c0b0a0c0b0a0b0c0a0c0b0a0c0c0a0b0c0b0c0b0a0b0c090b0a;
    encBuf[1048] = 256'h080a0a090c0b0a0d0b090b09010802040202030808000d0a000a010702040501;
    encBuf[1049] = 256'h02020008000a0b000c08020801050809000f0b0b0f0b0a0b0b0a0b0b090c0b0b;
    encBuf[1050] = 256'h0f0b0b0d0b0a0b0c090a0a090a0b090d0b0a0c0b0a0b0a000a00020801040001;
    encBuf[1051] = 256'h0300020701020601030501030402020402020402020302030501020402030401;
    encBuf[1052] = 256'h02030000010909000a08020901050808000f0b0a0f0a0a0b0a080a0800090908;
    encBuf[1053] = 256'h0e0a0b0d0b090b09010002050103030100020800050104070303060203030202;
    encBuf[1054] = 256'h0401020303040502040303030303020302020302030602020401020200010109;
    encBuf[1055] = 256'h01010a00020a00000b09000d09000c09000c09080d0800080307030505020403;
    encBuf[1056] = 256'h0203030204040304050304040203030303030303050304040304030304020102;
    encBuf[1057] = 256'h020101020203040304030102010809090b0a090a00000000090b0e0d0c0c0b0c;
    encBuf[1058] = 256'h0a0b0a0a0a090a0a0b0c0b0b0c0a0a0809010202050303050402040502040304;
    encBuf[1059] = 256'h0303040403030404030305020303030402030304030305020304020203010302;
    encBuf[1060] = 256'h0203030205030203040102020001000802010803040104030004020805010005;
    encBuf[1061] = 256'h0301060202040302040201040302050202050302040302030402030302050302;
    encBuf[1062] = 256'h03030203020801000a00080b02080d080c0f0a0d0c0a0c0b0a0b0b0b0b0d0b0d;
    encBuf[1063] = 256'h0b0c0c0b0c0a0b0b0b0b0a0b0c0b0c0c0a0c0a0b0a0a090a0909090a0a0a0d09;
    encBuf[1064] = 256'h0a0a080008040302050302040302050302060302040302040302040303040402;
    encBuf[1065] = 256'h0303020402020303030503020403020302000201000203020603030502010200;
    encBuf[1066] = 256'h0900080a02030107050103020101000900080a04030307050104010101010800;
    encBuf[1067] = 256'h000802020105020003010a000c0e090b0d090a0a0a0a0c0a0c0c0c0c0b0c0c0b;
    encBuf[1068] = 256'h0b0c0b0c0b0b0b0c0c0a0c0b0b0c0b0b0c0b0b0c0a0b0b0c0a0b0c0a0c0a0b0b;
    encBuf[1069] = 256'h0b0b0b0b0b0c0a0a0a0a090a0a0a0a0a09090802040405040304030203030303;
    encBuf[1070] = 256'h0503050503030503030303030303030403040404030304020302010201010203;
    encBuf[1071] = 256'h0405020402030201010000000001020305030403020201000100090101010503;
    encBuf[1072] = 256'h0205020102010001080b080c0d090b0c090a0b090b0c0c0d0c0c0d0b0c0b0c0a;
    encBuf[1073] = 256'h0c0a0a0c0a0c0b0c0b0d0b0c0b0b0b0c0a0b0c0a0b0c0c0a0c0b0b0c0a0c0a0a;
    encBuf[1074] = 256'h0b0b0b0b0c0b0c0b0c0a0b0b0c0a0a0a0a0a0b0a0b0b0b0b0c0a0a0a08080801;
    encBuf[1075] = 256'h0201040303050403040503040304030502030402030402040302030403030303;
    encBuf[1076] = 256'h0403030403030403030303030303020303030502030303010202000800090801;
    encBuf[1077] = 256'h0102040202020b0c0d0d0b0b0b09000003050100000c0c0c0c0c0a0909000008;
    encBuf[1078] = 256'h01090b0d0f0b0c0b0c0a0b0b090b0c0a0d0c0b0d0b0b0c0b0b0c0b0a0c0c0a0c;
    encBuf[1079] = 256'h0b0b0d0b0a0c0a0b0b0c0a0b0c0a0c0b0a0b0b0b0c0b0b0b0c0a0c0a0a0b0b0a;
    encBuf[1080] = 256'h0a0a090a0a000908010801050104060204030403050203040303040304030403;
    encBuf[1081] = 256'h0403030402030402020303040303040302030302020201020201020401010200;
    encBuf[1082] = 256'h09080e0b0a0d0a0a0a0a0a0a0b0b0f0b0b0d0a0b0b0a090908000908080a0a09;
    encBuf[1083] = 256'h0b09020307060303050202030202040203060204030303030202020800020900;
    encBuf[1084] = 256'h030801030b0b0c0f0f0a0c0c0a0b0b0b0c0b0b0c0c0b0c0c0a0c0b0b0b0b0c0a;
    encBuf[1085] = 256'h0b0a0c0a0b0b0b0b0d0a0a0a0a09080801010204020304030404030603040403;
    encBuf[1086] = 256'h0403030403040303030404030303040304030203030303040203030204020201;
    encBuf[1087] = 256'h020001000908090b0b0b0e0b0b0d0b0c0c0b0b0d0b0b0b0c0b0b0c0a0b0b0a0b;
    encBuf[1088] = 256'h0b0b0a0b0a0a0908020305050503030503040304030403040403040303040303;
    encBuf[1089] = 256'h03040303030402040203020303030302030102010008090a0b0c0c0c0b0c0c0b;
    encBuf[1090] = 256'h0d0b0b0d0b0b0d0a0b0b0b0b0c0a0b0b0b0c0b0b0c0b090a0900000102030305;
    encBuf[1091] = 256'h0302050304050304040304030402040203020403030304030402030203020302;
    encBuf[1092] = 256'h020302020201020008090b0c0d0b0d0b0c0c0b0b0d0b0b0d0a0b0c0b0b0b0c0b;
    encBuf[1093] = 256'h0b0b0c0c090b0a0a0b0a090a0a00080801020105040204050204030306030204;
    encBuf[1094] = 256'h0304030304030402040303030403030402030302030303040202030302030201;
    encBuf[1095] = 256'h02000a080b0d0b0c0c0b0c0c0a0b0d0a0c0b0c0b0c0a0c0b0a0b0b0b0b0c0a0b;
    encBuf[1096] = 256'h0c0a0a0c090a0b09090900000802010003010004020207040305040203030202;
    encBuf[1097] = 256'h020101010002030204030201080c0d0d0c0c0b0b0c0a0c0a0a0c0b0d0b0d0b0c;
    encBuf[1098] = 256'h0a0c0a0a0b0a0a0b0b0b0c0b0c0b0c0a0b0b090a0a0808080000000101080303;
    encBuf[1099] = 256'h0307040306030403040304030304020303040204030304030304030202020102;
    encBuf[1100] = 256'h0201020303040403030200000a0d0c0b0d0a0b0a0a0a0a0a0b0e0c0c0c0b0c0c;
    encBuf[1101] = 256'h0a0a0b0a0a0a0a0b0c0b0d0c0b0c0a0b0b0a090a09090a0a0b0e0b0c0b0b0a0a;
    encBuf[1102] = 256'h09080000010008090c0c0b0d0a0a0a080000010100000a0d0c0c0c0b0b0c0a0a;
    encBuf[1103] = 256'h0a0a0b0d0a0d0b0c0c0b0c0b0b0b0b0b0b0c0b0b0b0d0a0c0b0b0c0b0b0b0a0a;
    encBuf[1104] = 256'h0a08080000020001020001030307050404040304040203030202030305030403;
    encBuf[1105] = 256'h05030304020202020201020103030405020203010100090a0a0d0a0a0a090008;
    encBuf[1106] = 256'h08010b0c0b0f0d0b0c0b0b0b0b0a0a0b0b0d0b0c0c0c0a0c0b0a0a0b090a0a0a;
    encBuf[1107] = 256'h0a0b0b0e0b0b0c0c090b0a090a09080a09080a0a080c0b090c09080900030204;
    encBuf[1108] = 256'h070101040000000809000a08030105060102040800010a0a080c080109020400;
    encBuf[1109] = 256'h02010a0c0b0f0b090b0901000504020402010202080103020605030504020402;
    encBuf[1110] = 256'h0303040204030304030404030303040303030303040203040203040203030202;
    encBuf[1111] = 256'h020101000808080908080a09090d0c0b0f0b0c0c0b0b0b0c0a0a0a0a0a0b0a0b;
    encBuf[1112] = 256'h0c0a0c0a0a0a0a09080808000801000001010404030505030404030403020402;
    encBuf[1113] = 256'h0202020101020002020103040102030808090c0c0a0b0b090901010001090e0c;
    encBuf[1114] = 256'h0c0d0b0a0a090801020304040203030403070304050304040303040302040303;
    encBuf[1115] = 256'h0403030503030502040303030502030304020302030402040203040203020302;
    encBuf[1116] = 256'h0201020202030303030202090a0d0e0b0d0b0c0b0b0b0d0b0b0d0b0c0b0c0a0c;
    encBuf[1117] = 256'h0a0a0b0b0a0b0c0a0c0b0a0b0b0a0a0a08080900010803030406030504040304;
    encBuf[1118] = 256'h0303030403030402030402030303030402020301020201020008090a0d0b0d0c;
    encBuf[1119] = 256'h0b0c0c0b0b0d0b0b0c0c0b0b0b0c0b0a0a0a090a0a090a0a09090b0001000405;
    encBuf[1120] = 256'h0206030305030304040204030304040203040303030303040202030202020202;
    encBuf[1121] = 256'h020202000008090c0c0c0c0b0c0b0b0b0d0b0c0c0b0c0c0b0c0b0b0b0b0a0b0c;
    encBuf[1122] = 256'h0a0b0c0b0c0b0b0c0a0a0a0909090a090a0c0b0c0b0b0a090002020703020402;
    encBuf[1123] = 256'h0202020102030206040305030304030204020202030204030304040203030203;
    encBuf[1124] = 256'h010808090b0c0a0c0a090b0a0b0d0c0c0d0b0c0b0a0b0c09090908080a090b0d;
    encBuf[1125] = 256'h0a0b0c0909080103020703020404010402020403040304030304020202020102;
    encBuf[1126] = 256'h000101010101000009090d0d0c0c0c0c0c0b0b0c0c0a0b0b0b0c0b0c0c0b0c0a;
    encBuf[1127] = 256'h0c0a0a0b0a0a0a0a0a0a0a090a0b0a0a0a080000040403060303040303030503;
    encBuf[1128] = 256'h04030305030403030203030302010102010201020203020008090c0e0c0c0c0b;
    encBuf[1129] = 256'h0c0b0b0b0c0b0b0b0d0b0c0b0c0b0b0a0b0a0a0a09090a090b0a0c0a0a090002;
    encBuf[1130] = 256'h0306040402040202010202030403060304040304030203020202020001000100;
    encBuf[1131] = 256'h00000108090a0d0d0b0e0c0a0c0b0c0b0b0c0c0b0b0d0b0c0c0b0b0b0c0b0b0c;
    encBuf[1132] = 256'h0b0b0c0b0b0c0a0c0a0b0a0b0b0a0b0a090b0a090a0909090808010203040503;
    encBuf[1133] = 256'h0405030503040403030403030304020304020303020303020402020203000002;
    encBuf[1134] = 256'h09090a0f0b0c0d0b0b0c0b0b0c0b0b0c0b0b0d0b0b0d0b0a0c0a0a0b0a0a0b0b;
    encBuf[1135] = 256'h090b0a0909000000020401030601030502040402040304030303040402020302;
    encBuf[1136] = 256'h02040101020001010800010800000b0b090f0d0a0d0b0b0d0c0a0b0c0a0c0b0a;
    encBuf[1137] = 256'h0b0c0a0b0b0a0b0b0b0d0b0b0d0a0b0b0a090908000102030203030002030104;
    encBuf[1138] = 256'h0503060403050303040402030402030403030303030401030201020401030501;
    encBuf[1139] = 256'h03040203030201020900000c09080a00010004050102020808080e0a0a0d0a08;
    encBuf[1140] = 256'h0a08000801020801040105040305040303030203020001000103070405040305;
    encBuf[1141] = 256'h0303030401020201010001010302030603030403020202010009090a0c0b0b0c;
    encBuf[1142] = 256'h0b0a0c0b0b0b0b0c0b0b0b0b0a0b0b0c0e0b0b0e0b0c0a0a0908020504040404;
    encBuf[1143] = 256'h0204020102020102020304040404040304030304020303030302030303030302;
    encBuf[1144] = 256'h030203030305030404030304020201090a0c0d0b0d0b0a0a0a08000003030103;
    encBuf[1145] = 256'h000a0a0c0f0a0a0b090808040402050402030303040301030302040201030302;
    encBuf[1146] = 256'h05030307030305030305020202010000080a0a0b0b0a09080204030602020202;
    encBuf[1147] = 256'h09080a0f0a0c0c0a0a0c0a0a0a09080a000008020809000a0f090b0e090a0a08;
    encBuf[1148] = 256'h0000040403060303040302040200030101020302070303060303050302030302;
    encBuf[1149] = 256'h03010101010800010902010003030105020002090e0a0d0e0a0c0c0b0b0d0a0a;
    encBuf[1150] = 256'h0b090a0b09090b0a0a0c0a0b0e0a0b0c0a0b0c09090a00000004030305030103;
    encBuf[1151] = 256'h0200020100030303070503040303040303030201020009080b0d0a0b0c090b0a;
    encBuf[1152] = 256'h080a0a080a0d0b0f0c0b0d0b0c0c0b0b0c0b0b0b0b0b0a0b090a0a090a0b0b0c;
    encBuf[1153] = 256'h0e0a0b0c0a0a0a09000002030405030204030203030204020203020304040306;
    encBuf[1154] = 256'h030305030203020101080b0a0d0c0b0c0b0a0b0a0b0b0b0b0d0c0b0d0c0c0c0b;
    encBuf[1155] = 256'h0c0c0b0b0c0a0b0b0a0a0b0b0b0c0b0b0d0b0b0c0b0b0b0c0a0b0b0a0b0a0909;
    encBuf[1156] = 256'h0800000302030202010109090000010704040504030402040201020101000009;
    encBuf[1157] = 256'h0a090b0b0a0c0a090b0b0a0e0c0c0d0b0d0c0c0a0c0b0b0d0a0b0b0b0a0b0c09;
    encBuf[1158] = 256'h0b0a0a0b0c0b0d0b0c0b0c0a0b0a0a0a08080000010100020801020001050103;
    encBuf[1159] = 256'h070102030203060103040202040102030008010a0a080d0a080c0a080b0a080d;
    encBuf[1160] = 256'h0b0a0f0c0a0d0b0c0b0c0b0b0c0a0a0a0a0a0b090c0b0b0c0c0a0b0c090b0b0a;
    encBuf[1161] = 256'h0b0b0a0b0b080a09020003070101030001030900040003070304060203030303;
    encBuf[1162] = 256'h040202030001040101050102040202050101030000020908000900010a00030a;
    encBuf[1163] = 256'h09010e0b080d0a010a08020b09080f0d0a0d0b0a0b0900080206020204020102;
    encBuf[1164] = 256'h0900000800020105070202050203040203040203030204030204030304030204;
    encBuf[1165] = 256'h040103030303050102040101010000000900020003060205040102020000000a;
    encBuf[1166] = 256'h09090a0801010306020403020403030403040305020303020402020403040403;
    encBuf[1167] = 256'h0404030304030303040203030204030204030404030404030303030302020201;
    encBuf[1168] = 256'h0102030404040305030203040202020202020103020002010002030307050204;
    encBuf[1169] = 256'h0401030201010109000808000101050402050402030402040301030201020108;
    encBuf[1170] = 256'h0303030704030503020403020402020302020303010402000304020504030503;
    encBuf[1171] = 256'h02030302010009080a0c08000903030107040103020104020003010900090d08;
    encBuf[1172] = 256'h090b010300070601040301030301020108020208040301060302050401040202;
    encBuf[1173] = 256'h02020001010a00080b00000904020905010901080d000b0d090b0e0a0c0c0b0b;
    encBuf[1174] = 256'h0e090a0b080909000009000a0d0a0c0c0b0b0c0a0a0a08080901010804010002;
    encBuf[1175] = 256'h010a020a0e080a0c08080a03040107030103020002000b090c0d090b0d090b0c;
    encBuf[1176] = 256'h08090a00080901000c080d0e0a0c0d0a0b0b0a0a0b09080a08090a09090d090b;
    encBuf[1177] = 256'h0d0a0b0c0a0c0b0a0b0b090908030202070301030100010a0c090b0c0a0b0c08;
    encBuf[1178] = 256'h000804030306030201000b0c0e0d0b0c0b0a0b0b0a0a0a080a0c0b0d0c0c0b0d;
    encBuf[1179] = 256'h0b0b0d0a0b0b0b0c0b0a0b0b0a0b0b0b0b0c0b0c0c0b0c0c0a0b0b0a0b0b090a;
    encBuf[1180] = 256'h080000010302030402010108090a0b0a0801030705050303030302020000090b;
    encBuf[1181] = 256'h0c0b0c0d0a0c0b0b0c0b0b0d0b090b0c0a0d0b0c0c0c0b0c0b0b0c0b0a0a0a09;
    encBuf[1182] = 256'h09080908090a0a0d0b0c0c0b0a0b090900010304050402030203020101010001;
    encBuf[1183] = 256'h030101060102040101040002030000020a0c0a0f0e0a0c0c0a0c0a0a0b0a0a0b;
    encBuf[1184] = 256'h0b0a0d0b0b0e0b0b0d0b0b0c0b0a0b0a0a0b0a090a0a0a0b0b0b0d0a0b0c0b0a;
    encBuf[1185] = 256'h0b0a080900030206050304040304030202030001030801030204060204050202;
    encBuf[1186] = 256'h040102010000000a0a080b0b090b0a000b0a090f0b0a0f0a0b0c0c0a0b0b0a0d;
    encBuf[1187] = 256'h0b090c0a0a0a0b090a0a080a09000b0a080c0a090b0802010705030604020304;
    encBuf[1188] = 256'h0303030203040202030303060203040303050202030101020800000a0a090c0b;
    encBuf[1189] = 256'h090d0a090d0a090d0a0a0c0c0a0b0d0a0c0b0a0c0a0a0a0a090a09080a09090b;
    encBuf[1190] = 256'h0b0a0e0a09090801000505020405020304020304020203020304030305030305;
    encBuf[1191] = 256'h0303040303040203030202040101010001000800010802030204040002020b0c;
    encBuf[1192] = 256'h0b0f0c0a0c0b0a0b0a080909080908080b0a0b0f0a0b0c0b090b0a0000030504;
    encBuf[1193] = 256'h0504020403020304010303020304030404030404030403040304020303020202;
    encBuf[1194] = 256'h0101010100020202050203040203020008080b0d0b0d0b0c0b0b0b0c0b0a0b0b;
    encBuf[1195] = 256'h0a0c0b0a0c0b0c0c0b0b0c0a0b0a090a08010005040305030403040203030202;
    encBuf[1196] = 256'h0203040503060304040304030303030202020102010203030503030503030303;
    encBuf[1197] = 256'h03030202010009090b0d0c0b0c0b0b0a090b000100010208000b0f0c0d0b0c0a;
    encBuf[1198] = 256'h0c09090901010306030304030203020002000802030307050304040304040203;
    encBuf[1199] = 256'h030303030303020102020102040205040306020304020202020000080b090b0c;
    encBuf[1200] = 256'h0a090a010000050202030208010b0f090c0d0a0a0b0a090a0000000302000503;
    encBuf[1201] = 256'h0801010801090d01000a04020107050205030304040103030003010001010003;
    encBuf[1202] = 256'h040207030304030304030103010801080a00090a00080a050201060201040108;
    encBuf[1203] = 256'h01080c090b0e090b0b09090b02010805030004020804000b01090c000a0d0101;
    encBuf[1204] = 256'h0904040106020204010003000901080a00080a05020107040105020103020102;
    encBuf[1205] = 256'h010901090a00000b05030106040104030104020003000902080c080a0c090a0d;
    encBuf[1206] = 256'h00080902000904000b000c0f0a0b0f090a0c09090b08090a08090c080a0d090a;
    encBuf[1207] = 256'h0d0a0a0b0a0a0c09090a00080902000804000902000a03080c01000a02010007;
    encBuf[1208] = 256'h030207040104020102010800090c090b0d09090a00000902090c080c0f0a0b0d;
    encBuf[1209] = 256'h0a0c0c0a0b0b0b0c0b0a0c0c090b0b0a0c0a0b0b0c0a0c0b0b0c0b0b0b0c090a;
    encBuf[1210] = 256'h0a09090900080900090c090a0b0a090901030506040304020203020002090800;
    encBuf[1211] = 256'h090a00090c090b0d090c0c0a0c0b0d0b0c0b0e0b0c0c0c0b0c0b0b0c0b0b0c0b;
    encBuf[1212] = 256'h0a0b0c0a0c0a0c0a0c0a0b0b0c0b0b0a0b0b0b0b0a0b0b0b0b0b0c0a0b0b0b0b;
    encBuf[1213] = 256'h0a0909000000030405040303070201030202030101020009010a080209080408;
    encBuf[1214] = 256'h09020f0b0a0f0d0a0d0b0b0d0b0a0c0b0a0c0b0a0b0c0a0c0b0a0c0b0b0c0c0a;
    encBuf[1215] = 256'h0b0b0a0c0a0a0b0a090a0a080a09000909020a08030900070001060103050303;
    encBuf[1216] = 256'h050202040102020102030002030103060002030801030a0a010f0c0a0c0c0a0d;
    encBuf[1217] = 256'h0b090c0b0a0c0a0a0b0c0a0b0c0a0c0b0b0c0b0b0c0b0b0b0c090b0a080a0900;
    encBuf[1218] = 256'h0909010800020801040004060103060203060202040202040202030203040103;
    encBuf[1219] = 256'h050102040102040101040001020000020808000a08080c09000c09000a0a000c;
    encBuf[1220] = 256'h09080e0b090d0a090c0a090b0801090205000305020304020305020305020403;
    encBuf[1221] = 256'h0305030305030304030305030203040203030303050202040202030303030303;
    encBuf[1222] = 256'h040101020000010801010800010801030908080c0a0c0d0a0b0e090a0b0a0909;
    encBuf[1223] = 256'h0001010406020503020503030304030403040304030503030503030403030403;
    encBuf[1224] = 256'h0303030403030304030305020303040203030303020303020303020304020203;
    encBuf[1225] = 256'h0203050203040302030202030901030a08030103060206040203040204020203;
    encBuf[1226] = 256'h0301050202040401030502030402040303040302040302030302030302040301;
    encBuf[1227] = 256'h05020204020203030103020803000a03010b04010b02080e00090e090a0c090b;
    encBuf[1228] = 256'h0b090b0c090a0c000a0b010a0c04000a05020004020904010802020905020006;
    encBuf[1229] = 256'h020205030104020103020104030004020004020802010b02090d00090d08090c;
    encBuf[1230] = 256'h08090c090a0e09090c0a0a0c09090c080a0b0a0a0d090b0b0a0b0d080a0a0009;
    encBuf[1231] = 256'h0b01090c01090d02080a04010805020805010003000803080b04000902080b02;
    encBuf[1232] = 256'h0a0f080a0c090b0d080b0c080a0c090c0c090a0d0b0b0c0b0b0e0a0a0c0a0b0c;
    encBuf[1233] = 256'h0a0b0b0b0b0d0a0a0b090b0b0a0b0b0b0c0c0a0a0c090b0b0a0a0c080a0a0809;
    encBuf[1234] = 256'h0a01090903010004020206020102010104010002090b080b0e0b0c0c0c0b0d0a;
    encBuf[1235] = 256'h0c0b0a0b0c0a0c0b0b0c0b0c0b0c0b0d0b0b0c0b0b0c0b0b0c0b0b0b0c0b0b0b;
    encBuf[1236] = 256'h0b0c0a0b0b0b0a0c0a0a0a09090a000008010302030303040401010202040305;
    encBuf[1237] = 256'h040203050202040202040100020008000a0b0b0f0d0a0d0b0b0c0c0a0c0b0a0c;
    encBuf[1238] = 256'h0c0a0b0b0c0b0c0b0b0c0a0b0c090b0a0a0b0a0b0d0a0b0c0a0a0b0a0a0b0908;
    encBuf[1239] = 256'h0808020203050205040304040203040203040103030103030303050103040002;
    encBuf[1240] = 256'h030001010908010b0a010e0b000d0c0a0d0c0a0d0c0a0b0c0b0b0d0a0b0b0b0c;
    encBuf[1241] = 256'h0b0a0c0a0a0b0b090b0a0a0b0b0a0c0b0a0c0a090a0900000204030604020305;
    encBuf[1242] = 256'h0203050203050303050204030203040202030302030303030203030202030001;
    encBuf[1243] = 256'h020900020c0a000d0a0a0f0b0b0e0b0b0d0b0b0c0b0b0c0b0a0c0a0a0b0b0a0b;
    encBuf[1244] = 256'h0a080a0801010306030603040304030403040304020304030304030403030404;
    encBuf[1245] = 256'h0203040303040203030204020201030101010100000808090c0a0b0d0b0b0d0b;
    encBuf[1246] = 256'h0b0b0b0c0b0a0b0c0b0a0c0b0c0b0a0d0b0a0b0c0a0a0a0a0a0a000801030405;
    encBuf[1247] = 256'h0503050304030403040303040304020402020402030303030502030402030304;
    encBuf[1248] = 256'h02030304030304030303030303020201020808000a0a0a0b0b0b0a080909080a;
    encBuf[1249] = 256'h0901000802010804020104020004020005030803050103040206030205030305;
    encBuf[1250] = 256'h040204030304030304030303030203030202010202000000010808000908090a;
    encBuf[1251] = 256'h080a09080b0c0a0c0c0b0d0c0b0d0c0a0b0c0a0c0a0b0b0d0a0a0b0a0b0b0a0a;
    encBuf[1252] = 256'h0a08080801000903000b000b0d090b0d090a0b00090a01000902010005020004;
    encBuf[1253] = 256'h040105020204020203030004020001020803000903000a020200040302070402;
    encBuf[1254] = 256'h0503030403020502010302010202010202000201000502010305020403020502;
    encBuf[1255] = 256'h0103020103010003000901080b080c0e0a0c0c0b0d0b0a0c0b0b0b0b0a0b0b0a;
    encBuf[1256] = 256'h0b0c090c0b0b0c0c0b0d0b0b0c0c0b0c0b0b0c0b0a0c0b0a0a0b0b0a0b0b0c0a;
    encBuf[1257] = 256'h0a0c0a0a0b0b0b0c0c0a0c0b0c0c0b0b0c0c0b0b0c0b0b0b0b0c0a0b0b0b0b0b;
    encBuf[1258] = 256'h0b0b0c0b0b0d0b0b0e0b0b0d0b0c0b0c0a0b0b0b0a0b0a0b0b090b0a0a0b0a09;
    encBuf[1259] = 256'h0809020303060303040203030302040304030504040304040403030404030304;
    encBuf[1260] = 256'h0304030304030303020303020203020202040202030203030102010808080a0b;
    encBuf[1261] = 256'h090b0b0c0b0e0b0c0c0c0b0d0b0b0c0c0b0b0b0c0b0b0c0b0b0b0b0a0b0a0b09;
    encBuf[1262] = 256'h0a090b0b0b0e0b0d0b0c0b0c0a0b0b0b0b0b0b0b0b0d0b0b0c0b0c0b0a0b0c09;
    encBuf[1263] = 256'h0b0d090b0d0b0c0c0b0c0c0a0c0b0a0c0b0b0c0b0c0b0b0b0c0b0b0b0c0a0a0b;
    encBuf[1264] = 256'h0a0b0c0a0c0b0b0c0b0b0c0b0b0b0a0a0b090809000100030503060403040403;
    encBuf[1265] = 256'h0403040304030403030502030403030403030502030304030403030403030403;
    encBuf[1266] = 256'h0303030304030203030304020203020302030203020303030204020302020101;
    encBuf[1267] = 256'h0908090d0a0b0d0a0b0c0b0b0c0b0c0d0a0b0b0b0c0b0a0a0a0a0909090a0b0c;
    encBuf[1268] = 256'h0c0c0c0d0b0c0c0b0c0b0c0b0c0b0c0b0b0d0b0b0b0d0b0b0c0b0c0b0b0c0b0c;
    encBuf[1269] = 256'h0b0c0a0c0b0a0c0b0b0b0c0b0c0a0b0b0c0a0b0b0b0b0b0b0c0a0a0a0a090a09;
    encBuf[1270] = 256'h0809080008020301060402050403040403040403040303050303040304030304;
    encBuf[1271] = 256'h0304020402030304030304020402030303040303040303030502030302040203;
    encBuf[1272] = 256'h020402020202030202030302030302040201020201020200020109000a0e090d;
    encBuf[1273] = 256'h0c0a0d0b0b0d0b0b0d0b0b0c0b0c0b0c0c0b0b0c0b0c0b0c0b0b0c0b0c0b0b0c;
    encBuf[1274] = 256'h0c0b0b0c0b0b0c0c0a0b0b0c0b0b0c0b0b0b0c0b0b0c0b0b0c0a0b0c0a0b0b0b;
    encBuf[1275] = 256'h0b0c0b0b0b0b0c0a0a0b0a0a0a0a090909080801020206030306040204030403;
    encBuf[1276] = 256'h0403050203040402030403030403050203040303040303040304030303040303;
    encBuf[1277] = 256'h0502030303040304020402030302040203030304020402020302030302030401;
    encBuf[1278] = 256'h020201010100010809090a0d0a0d0b0c0c0b0b0d0c0a0b0d0a0c0b0b0c0b0c0b;
    encBuf[1279] = 256'h0c0b0b0c0b0c0b0b0c0b0b0c0b0b0c0b0b0c0b0b0c0b0b0c0b0a0c0b0a0c0a0b;
    encBuf[1280] = 256'h0b0b0c0b0b0b0c0a0b0c0a0b0a0b0b0b0a0c0a0a0a0b0a0a0b0a0a0b090a0a00;
    encBuf[1281] = 256'h0900040104050304050204030404030305030305030304030404020304030403;
    encBuf[1282] = 256'h0304030304040203040303030404020304030303040303040203040203030303;
    encBuf[1283] = 256'h0403030402030302040202020201020100010008000a0a0b0d0c0b0d0c0b0c0b;
    encBuf[1284] = 256'h0c0c0b0c0b0c0b0c0b0b0c0b0b0d0b0a0c0b0a0c0b0b0b0c0b0c0b0b0c0a0b0c;
    encBuf[1285] = 256'h0a0b0b0b0c0b0b0b0b0c0b0b0b0c0b0b0b0c0b0a0c0a0a0b0a0b0b0a0c0a0a0b;
    encBuf[1286] = 256'h0b0b0b0c0a0a0b0a0a0a08090001010205020306020304030404030404030404;
    encBuf[1287] = 256'h0303050304030304040204030303040403030403030404020304020402030304;
    encBuf[1288] = 256'h0203040203040203030304030304030203040203020302030203020302020102;
    encBuf[1289] = 256'h010001080a090b0f0a0d0b0c0c0c0a0c0b0b0d0a0b0c0c0a0b0c0a0c0b0a0c0b;
    encBuf[1290] = 256'h0b0d0a0b0b0b0c0b0c0a0b0b0c0b0b0b0c0b0c0b0b0b0c0a0c0a0b0b0b0b0c0b;
    encBuf[1291] = 256'h0b0b0c0b0b0b0b0c0c0a0a0b0b0b0c0a0a0b0b0b0b0a0b0b090b0b0a0b0a090b;
    encBuf[1292] = 256'h0a00090005010506020306020305020403030403030503030403030503040303;
    encBuf[1293] = 256'h0403040303040304020304030204030303040304030303040303030403030304;
    encBuf[1294] = 256'h0303030403030303040303040203030203030203030201020001010808080a0a;
    encBuf[1295] = 256'h0c0c0b0e0b0c0d0b0c0c0b0b0d0b0c0b0b0c0c0a0b0c0b0c0b0b0c0c0a0b0c0b;
    encBuf[1296] = 256'h0b0d0a0b0b0b0c0b0c0b0b0b0c0b0b0c0b0c0a0c0a0b0b0a0c0b0a0b0c0a0b0b;
    encBuf[1297] = 256'h0a0c0a0a0b0b0b0b0b0b0c0a0a0b0a0909090808000201030602030602030403;
    encBuf[1298] = 256'h0404020403040304030403030404020402030304020402030402030403030403;
    encBuf[1299] = 256'h0304030303040304030204030303040304030304030304020402030303030403;
    encBuf[1300] = 256'h03040302040203030402030303030303040202020202010100010808090b0c0b;
    encBuf[1301] = 256'h0e0b0c0d0c0a0d0a0c0b0b0c0c0b0b0c0b0b0d0a0b0c0b0b0c0c0a0b0c0a0c0a;
    encBuf[1302] = 256'h0b0b0b0c0b0b0c0b0b0b0c0a0b0c0a0b0b0b0c0a0b0b0b0b0b0b0b0b0b0b0a0b;
    encBuf[1303] = 256'h090a0a0809000101020502060304040304040402040303040303050203040302;
    encBuf[1304] = 256'h0403030304030403040303040304030303040303040303040303040402030303;
    encBuf[1305] = 256'h0403030403030305020303030305020303040303030403020402020303020303;
    encBuf[1306] = 256'h0203020203020202020002080a090d0d0a0d0c0b0d0b0c0c0b0b0d0b0b0d0b0a;
    encBuf[1307] = 256'h0d0a0b0c0b0b0c0b0c0b0c0a0c0a0b0b0b0c0b0b0b0d0a0b0b0c0a0b0c0a0b0b;
    encBuf[1308] = 256'h0c0a0b0b0a0b0b0b0c0a0a0a090a0a0909090808080101020306030404040205;
    encBuf[1309] = 256'h0203040303050204020304030304040203040203040303040203030304030303;
    encBuf[1310] = 256'h0402030402030402030402030402020303030303030402040202030303030402;
    encBuf[1311] = 256'h03030203030104020003020102020003010a00090d080c0d0b0c0d0a0d0b0b0d;
    encBuf[1312] = 256'h0b0b0c0c0a0c0b0b0b0d0a0c0b0b0c0b0c0b0c0b0c0b0b0c0b0c0b0b0c0b0b0c;
    encBuf[1313] = 256'h0b0b0c0b0c0a0b0c0a0b0b0b0c0a0b0b0b0b0c0a0b0b0a0b0b0b0c0a0a0a0909;
    encBuf[1314] = 256'h0a08000103040404050303050304030403040304030305020304030304030304;
    encBuf[1315] = 256'h0303040303040303030403040203030304030303030304030202040102020101;
    encBuf[1316] = 256'h020201020101020002010009090a0c0c0c0b0d0d0a0c0b0b0c0b0b0d0b0b0c0b;
    encBuf[1317] = 256'h0b0b0d0b0b0c0b0b0c0b0c0b0b0c0b0b0c0b0c0b0b0c0c0b0b0b0d0a0c0a0b0c;
    encBuf[1318] = 256'h0b0b0b0c0b0b0c0b0b0b0c0c0a0b0c0a0c0a0b0b0c0a0b0c0a0b0b0b0c0a0b0b;
    encBuf[1319] = 256'h0b0a0b0b0b0b0b0a0c0909090800080204020405020404030404030403040304;
    encBuf[1320] = 256'h0403030404030303050303040204030204020303040204020203030402030304;
    encBuf[1321] = 256'h020303030304030203020302030202020101010008080b0c0b0d0c0b0c0c0b0c;
    encBuf[1322] = 256'h0b0c0b0c0b0b0c0c0a0c0a0b0b0c0b0b0d0a0b0b0c0b0b0b0c0b0b0c0b0b0b0b;
    encBuf[1323] = 256'h0c0b0a0c0b0a0b0b0b0c0b0b0c0b0b0b0c0a0b0c0a0c0a0a0b0b0b0c0b0a0c0b;
    encBuf[1324] = 256'h0a0b0c0a0a0c090a0c090a0b0a0a0c0a0b0b0a0c0b090a0a0909000100030602;
    encBuf[1325] = 256'h0307020304030404020403040304030305030305030303040403030403030502;
    encBuf[1326] = 256'h0304030204030204030204020303040203030303040203030303040302030302;
    encBuf[1327] = 256'h0303020201020100090a090d0c0a0b0e0b0b0c0c0b0c0a0c0b0b0c0b0b0d0b0a;
    encBuf[1328] = 256'h0c0b0a0c0a0b0b0b0c0a0c090b0b0a0b0c0a0a0b0b0a0b0b0b0b0a0a0a090908;
    encBuf[1329] = 256'h0101000201030502020202040502020303040403040303040203040302030302;
    encBuf[1330] = 256'h0203040201020301010100000101080a090a090a0b0c0a0c0b0a0c0b0a0a0c0b;
    encBuf[1331] = 256'h0a0c090a0a090b0b08090a090809000200080204030303050402040402030304;
    encBuf[1332] = 256'h0403030403030602020403030403020403040202030402020304020203030304;
    encBuf[1333] = 256'h0204020203020104020003010002020801010802080a01000a02080c08090a00;
    encBuf[1334] = 256'h0a0c01080b02000a030400030301070300040400030202040301050301040302;
    encBuf[1335] = 256'h040302040203040101030300020109010809080d0d0a0b0e0a0b0e0a0c0b0b0d;
    encBuf[1336] = 256'h0b0b0d0b0b0c0c0a0b0c0b0c0a0c0a0b0c0b0b0b0d0a0b0c0a0b0c0a0b0b0b0b;
    encBuf[1337] = 256'h0c0b0b0b0b0c0a0b0b0b0a0b0b0a090b0a090800000203040504030404040303;
    encBuf[1338] = 256'h0503030503030503030305030304030304030303040304020303040203030403;
    encBuf[1339] = 256'h0203040302040202030202030402010302020202020302020103010801080900;
    encBuf[1340] = 256'h080b080b0b090a0b080d0b080b0d0a0d0b0a0f0a0a0c0b0b0d0b0b0c0c0a0c0b;
    encBuf[1341] = 256'h0a0d0a0b0c0b0b0c0b0c0c0b0b0c0b0c0b0c0b0c0a0b0c0b0c0b0a0c0b0b0b0d;
    encBuf[1342] = 256'h0a0b0b0c0a0c0a0a0b0b0b0b0c0a0c0a0a0a0b0b0a0a0b0b090b090908000102;
    encBuf[1343] = 256'h0307030404030404030404030305020403030305030304030304030403020403;
    encBuf[1344] = 256'h0304020304020303040203030304030203030204020202020202020102010000;
    encBuf[1345] = 256'h0008090a0b0c0c0c0d0a0c0b0c0b0c0c0a0c0b0a0c0b0c0b0b0b0c0c0a0b0c0a;
    encBuf[1346] = 256'h0c0a0b0b0b0c0b0c0a0c0a0a0c0a0b0b0b0c0b0c0b0b0b0c0b0b0c0b0b0c0b0b;
    encBuf[1347] = 256'h0b0d0a0b0a0b0d0a0a0c0a0a0b0b0b0c0b0a0b0c0a0b0b0a0b0b0a0b0b090b09;
    encBuf[1348] = 256'h000a010202060303070402040304030503040303050303040402040303040303;
    encBuf[1349] = 256'h0502030403020403030304030304030303040303030403020304020303020303;
    encBuf[1350] = 256'h020303010202020000080a0a0c0c0c0c0c0b0c0c0b0c0b0c0b0c0b0c0b0c0b0b;
    encBuf[1351] = 256'h0c0b0b0c0b0c0b0b0c0b0b0c0b0b0c0a0b0c0a0b0b0c0a0b0b0b0b0c0b0b0a0b;
    encBuf[1352] = 256'h0c0a0b0b0b0b0b0b0c0a0a0a0b090b0a090b09000a0802090106000206020204;
    encBuf[1353] = 256'h0304030306030204030205030204040203040204030305020304030304030305;
    encBuf[1354] = 256'h0203040303040204030303040303050203030402030402040202030304020303;
    encBuf[1355] = 256'h04020303020402020203020302020202020100000008090a0d0b0c0d0b0c0c0b;
    encBuf[1356] = 256'h0c0c0b0b0d0b0b0b0d0b0b0c0b0c0b0a0c0b0b0c0b0b0b0c0b0c0a0b0b0c0a0b;
    encBuf[1357] = 256'h0b0b0b0c0a0b0b0a0b0c090b0a090a0a08080901000004040204040204040303;
    encBuf[1358] = 256'h0502040303040402040302030502030402030402030304020402030302040302;
    encBuf[1359] = 256'h03030304030204020203030203030203030203040101010001010901000c0809;    

    decBuf[0] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[1] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[2] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[3] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[4] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[5] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[6] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[7] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[8] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[9] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[10] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[11] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[12] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[13] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[14] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[15] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[16] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[17] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[18] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[19] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[20] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[21] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[22] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[23] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[24] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[25] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[26] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[27] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[28] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[29] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[30] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[31] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[32] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[33] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[34] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[35] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[36] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[37] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[38] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[39] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[40] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[41] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[42] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[43] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[44] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[45] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[46] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[47] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[48] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[49] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[50] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[51] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[52] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[53] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[54] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[55] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[56] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[57] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[58] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[59] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[60] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[61] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[62] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[63] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[64] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[65] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[66] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[67] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[68] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[69] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[70] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[71] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[72] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[73] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[74] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[75] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[76] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[77] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[78] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[79] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[80] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[81] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[82] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[83] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[84] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[85] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[86] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[87] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[88] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[89] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[90] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[91] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[92] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[93] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[94] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[95] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[96] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[97] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[98] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[99] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[100] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[101] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[102] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[103] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[104] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[105] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[106] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[107] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[108] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[109] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[110] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[111] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[112] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[113] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[114] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[115] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[116] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[117] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[118] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[119] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[120] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[121] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[122] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[123] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[124] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[125] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[126] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[127] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[128] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[129] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[130] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[131] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[132] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[133] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[134] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[135] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[136] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[137] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[138] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[139] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[140] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[141] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[142] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[143] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[144] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[145] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[146] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[147] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[148] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[149] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[150] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[151] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[152] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[153] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[154] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[155] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[156] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[157] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[158] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[159] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[160] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[161] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[162] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[163] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[164] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[165] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[166] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[167] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[168] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[169] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[170] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[171] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[172] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[173] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[174] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[175] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[176] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[177] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[178] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[179] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[180] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[181] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[182] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[183] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[184] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[185] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[186] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[187] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[188] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[189] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[190] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[191] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[192] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[193] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[194] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[195] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[196] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[197] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[198] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[199] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[200] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[201] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[202] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[203] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[204] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[205] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[206] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[207] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[208] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[209] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[210] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[211] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[212] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[213] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[214] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[215] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[216] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[217] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[218] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[219] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[220] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[221] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[222] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[223] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[224] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[225] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[226] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[227] = 256'h010000000100feff010000000100000001000000010000000100000001000000;
    decBuf[228] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[229] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[230] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[231] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[232] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[233] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[234] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[235] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[236] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[237] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[238] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[239] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[240] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[241] = 256'h0100000001000000ffff00000100000001000000010000000100000001000000;
    decBuf[242] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[243] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[244] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[245] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[246] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[247] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[248] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[249] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[250] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[251] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[252] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[253] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[254] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[255] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[256] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[257] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[258] = 256'h0100000001000000010000000100020001000000010000000100feff01000000;
    decBuf[259] = 256'h0100000001000000ffff00000100000001000000fffffeff0100000001000000;
    decBuf[260] = 256'h01000000010000000100feff010000000100000001000000010000000100feff;
    decBuf[261] = 256'h0100000001000000010000000100feff01000000fffffeff0100000001000000;
    decBuf[262] = 256'h0100feff01000000010000000100000001000000010000000100000001000000;
    decBuf[263] = 256'h01000000010002000100000001000200ffff0000010000000100000001000000;
    decBuf[264] = 256'h0100000001000000010000000100000001000000fffffeff01000200ffff0000;
    decBuf[265] = 256'h01000000ffff000001000200ffff000001000000ffff00000100000001000000;
    decBuf[266] = 256'h01000000010000000100000001000000ffff0000010000000100000001000000;
    decBuf[267] = 256'h01000000ffff00000100000001000200ffff0000010000000100000001000000;
    decBuf[268] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[269] = 256'h010000000100000001000000fffffeff010002000100feffffff000001000000;
    decBuf[270] = 256'h010000000100feff0100000001000000010000000100feff0100020001000000;
    decBuf[271] = 256'h0100000001000000010000000100000001000000010000000100000001000200;
    decBuf[272] = 256'hfffffeff01000000ffff00000100000001000000010000000100000001000000;
    decBuf[273] = 256'h0100feff0100020001000000010000000100feff0100020001000000ffff0200;
    decBuf[274] = 256'h01000000010000000100000001000200ffff0000010000000100000001000000;
    decBuf[275] = 256'h01000000010000000100000001000000010000000100000001000200ffff0000;
    decBuf[276] = 256'h01000000010000000100000001000000010000000100000001000000ffff0000;
    decBuf[277] = 256'h01000000010000000100feffffff000001000000010000000100000001000000;
    decBuf[278] = 256'h0100000001000000ffff000001000000010000000100000001000200ffff0000;
    decBuf[279] = 256'h01000000010000000100000001000200fffffeff01000000fffffeff01000000;
    decBuf[280] = 256'h01000000010000000100feff01000200ffff0000010000000100000001000000;
    decBuf[281] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[282] = 256'h01000000010000000100feff0100000001000000010000000100000001000000;
    decBuf[283] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[284] = 256'h01000000010000000100000001000000ffff0000010000000100000001000000;
    decBuf[285] = 256'h0100000001000000010000000100000001000000010002000100000001000000;
    decBuf[286] = 256'h010000000100000001000200ffff000001000200fffffeff0100000001000000;
    decBuf[287] = 256'h010000000100000001000000fffffeff01000000010000000100000001000000;
    decBuf[288] = 256'h0100000001000200010000000100000001000000010000000100000001000000;
    decBuf[289] = 256'h01000000010000000100feff010000000100feff010000000100feff01000000;
    decBuf[290] = 256'h0100000001000000010000000100feff0100020001000000ffff000001000000;
    decBuf[291] = 256'h0100000001000200ffff000001000000ffff000001000200ffff0200fffffeff;
    decBuf[292] = 256'h01000000010000000100000001000000ffff0000010000000100000001000000;
    decBuf[293] = 256'h0100feffffff00000100000001000000010000000100000001000000fffffeff;
    decBuf[294] = 256'h01000200ffff00000100000001000000fffffeff01000200ffff00000100feff;
    decBuf[295] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[296] = 256'h010000000100feff010000000100000001000000010000000100000001000200;
    decBuf[297] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[298] = 256'hffff000001000000010002000100000001000000010000000100000001000200;
    decBuf[299] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[300] = 256'h010000000100000001000000fffffeff01000200fffffefffffffeff01000000;
    decBuf[301] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[302] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[303] = 256'h010000000100feffffff000001000000ffff0000010000000100000001000000;
    decBuf[304] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[305] = 256'h0100feff01000200010000000100000001000000010000000100000001000200;
    decBuf[306] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[307] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[308] = 256'h010000000100020001000000ffff000001000000010000000100000001000000;
    decBuf[309] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[310] = 256'h0100000001000000010000000100000001000200ffff00000100000001000000;
    decBuf[311] = 256'h01000000010000000100000001000000010000000100feffffff00000100feff;
    decBuf[312] = 256'hffff00000100000001000000010000000100feff010000000100000001000200;
    decBuf[313] = 256'h010000000100000001000000010000000100000001000200ffff00000100feff;
    decBuf[314] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[315] = 256'h0100000001000000010000000100feff01000000fffffeff01000200fffffeff;
    decBuf[316] = 256'h01000000010000000100000001000000010000000100000001000200fffffeff;
    decBuf[317] = 256'hffff000001000000010000000100feffffff00000100000001000200ffff0000;
    decBuf[318] = 256'h010000000100000001000000010000000100000001000000010000000100feff;
    decBuf[319] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[320] = 256'h01000200ffff0000010000000100000001000000010000000100000001000000;
    decBuf[321] = 256'h0100000001000200ffff0000010000000100000001000200ffff00000100feff;
    decBuf[322] = 256'h01000000010000000100000001000000fffffeff0100feff01000200ffff0000;
    decBuf[323] = 256'h01000000fffffefffffffeffffff00000100000001000200fffffeff01000200;
    decBuf[324] = 256'hfffffeff01000000010000000100000001000200fffffeff0100000001000000;
    decBuf[325] = 256'h01000000010000000100feffffff00000100000001000200010000000100feff;
    decBuf[326] = 256'h01000000ffff000001000000010000000100feff01000200ffff000001000200;
    decBuf[327] = 256'h01000000ffff000001000200ffff00000100feffffff00000100000001000000;
    decBuf[328] = 256'h010000000100000001000000010000000100feff01000200fffffeff01000000;
    decBuf[329] = 256'h0100000001000000010000000100000001000200ffff00000100000001000000;
    decBuf[330] = 256'h01000000010000000100000001000000010000000100feffffff000001000000;
    decBuf[331] = 256'h01000000fffffeff010000000100feffffff0000010000000100000001000000;
    decBuf[332] = 256'h0100000001000200fffffefffffffefffcfffbff01000c0018001300ffffeaff;
    decBuf[333] = 256'hf8ffffffecffdeffeffffeff0400100018000b00f4fff1fffaff01000d000f00;
    decBuf[334] = 256'h0d0008000a000b000f001b0028002d0029001500fdff0d002d002800eeffd6ff;
    decBuf[335] = 256'hddfff2ffdffffbff29002f001f00240032002d0012000800050007000f000800;
    decBuf[336] = 256'hf9fff3fff9fffdfff9ffe7ffcdffc2ffd2ffd5ffbdffcdfff8ff24001e002e00;
    decBuf[337] = 256'h45001600c5ffbaffecff0700deffb8ffa4ffb6ffc7ffe1ffe6ffeaffeeffe3ff;
    decBuf[338] = 256'hdaffe2fffaff160031002700f8ffacffcafff8ff1100450083005a0007002800;
    decBuf[339] = 256'h6e002e00b3ff59ffabfff4ff1c0029001e0000000900110009000300f0ffc8ff;    
    decBuf[340] = 256'h9aff94ff8eff94ffd9ff5b00250015005f00370099ffafff5f00e9ff51ff7800;
    decBuf[341] = 256'hef023d08830ad309730ae1095d09e4085209b5095b09ad09f809b40976093e09;
    decBuf[342] = 256'ha5081a089b0775070c07ed0643075d0716072b073f07e6065306f10598054705;
    decBuf[343] = 256'h5505e905720684067406470604062906600692068906a106c706ce0606077707;
    decBuf[344] = 256'h4a081309ca09410a2b0af009de09ef09e0093d0ac30a400bd20b340c460c360c;
    decBuf[345] = 256'h620c700c330ce60bc80b880b3e0b480b9a0bbb0bb10bba0ba10b4f0b020bbc0a;
    decBuf[346] = 256'h6a0af109c009940951092c0937092d09ee08b4087f08180876073507fa06e806;
    decBuf[347] = 256'hf906250732073e0749076707700779078f078807690763077d079407cb073c08;
    decBuf[348] = 256'hae08f7085509c209ee09fc09200a150a0b0a140a3e0a810ad30a360b790b9d0b;
    decBuf[349] = 256'h920b880b490bfe0ae00ad70acf0ad60add0acb0aa30a750a3d0a080ad809b909;
    decBuf[350] = 256'h9209630938091009e208b6088f0861081008c30769072c0721073f075a077307;
    decBuf[351] = 256'h6c0757072b07ed06d506cd06e206010728075707760787079607a407b907d407;
    decBuf[352] = 256'hed07fc0711081e082e08410854086008620864086208640871088b089f089b08;
    decBuf[353] = 256'h85085a08fd0784071207c906bb06af06a4069a066d062206c8055b05f4049604;
    decBuf[354] = 256'h5a0439042f0426040d040504f103de03cd03b3039c0376034803290318032703;
    decBuf[355] = 256'h51038303a603b903be03a5039703a303c60302043c048004c004d804e004e704;
    decBuf[356] = 256'h060539057605b005d605ea05f105e005d005c205ad058a0557050c05b2045d04;
    decBuf[357] = 256'h2604f403d903af036c0307038f021d0299013f010e01e200ba00960049001700;
    decBuf[358] = 256'hc5ff78ff46ff06ffdcfe99fe6bfe42fe1dfe08fe02fefcfde2fdb9fd86fd56fd;
    decBuf[359] = 256'h37fd3cfd56fd92fddcfd22fe75feacfedefe0bff34ff69ffb5fffbff4d009a00;
    decBuf[360] = 256'he000fb000301fc00e700d400c400be00b1009b00780046001500ddffa9ff86ff;
    decBuf[361] = 256'h67ff4bff27ff07ffe9fecefeaefe88fe50fefdfd9afd3dfdcffca3fc60fc54fc;
    decBuf[362] = 256'h33fc01fcaffb62fb1cfbdcfab3fa8dfa6bfa3ffa0dfaddf9caf9c4f9def907fa;
    decBuf[363] = 256'h3afa6afa89fa9afa9ffa9bfa97fa9afabafae9fa21fb73fbc0fbf2fb20fc39fc;
    decBuf[364] = 256'h31fc0ffcd7fba2fb80fb6dfb7efb98fbaffbaafb97fb63fb2efbfefac6faaffa;
    decBuf[365] = 256'ha8faa2fa91fa82fa61fa33faeef9aef974f94ff948f94ef95ff95af943f903f9;
    decBuf[366] = 256'hb1f84ef8f0f7b4f793f7b1f7def739f88ef8c5f8bbf88df843f8e9f7acf78bf7;
    decBuf[367] = 256'hbdf722f89af80cf973f99bf98ff96ef928f9fbf8f2f809f939f97ef9bef9f7f9;
    decBuf[368] = 256'h2cfa40fa3afa1efae6f9b1f981f955f939f93ef930f924f9f9f8b0f856f819f8;
    decBuf[369] = 256'hccf7aef7b7f7aff7a8f778f733f7cef671f634f6fdf5f3f5fcf515f62cf640f6;
    decBuf[370] = 256'h53f64df61ff6daf5adf573f55df57ff5abf5f4f53af67af692f6a9f6a2f6a8f6;
    decBuf[371] = 256'hb9f6c9f6e9f618f750f793f7e6f71df84ff88ef897f8adf8c2f8e1f814f952f9;
    decBuf[372] = 256'h7bf991f998f985f95ef93af91af90df909f9f8f8e8f8daf8b8f897f879f847f8;
    decBuf[373] = 256'h09f8cff77df730f712f709f701f717f710f7f1f6bef680f647f621f60df6faf5;
    decBuf[374] = 256'hfff5e6f5cff5c2f5a7f5a3f5b3f5bcf5d8f5fbf512f630f65bf682f6b0f6e9f6;
    decBuf[375] = 256'hfff62ff75bf782f7bbf70df844f88af8caf8e3f8eaf8f1f8ebf8daf8dff8dbf8;
    decBuf[376] = 256'hdff8faf819f948f974f990f99ff99bf97df96af966f95df965f978f971f959f9;
    decBuf[377] = 256'h37f9fbf8c1f89cf879f84df831f8f9f7c4f794f775f764f769f765f769f76df7;
    decBuf[378] = 256'h5bf758f772f792f7c9f7fdf72df84df874f898f8c2f8f4f824f944f96bf97af9;
    decBuf[379] = 256'h91f9b8f9e6f912fa4ffa79fa8ffa96fa90fa95faa5fab3fab7fac3fab8faaffa;
    decBuf[380] = 256'hb7fabffae3fa11fb30fb41fb46fb26fb08fbf5fae3fad4facbfaa4fa7cfa4efa;
    decBuf[381] = 256'h16fafff9ebf9d8f9c7f9adf984f95cf943f935f939f94df965f987f9b1f9d8f9;
    decBuf[382] = 256'h07fa3ffa73fab1fadafa00fb30fb68fb9dfbe8fb2efc5cfc75fc7cfc83fc96fc;
    decBuf[383] = 256'hbdfcf6fc39fd79fdb3fdd8fdedfde7fde1fddcfdcefdcafdbefdb4fdaafda7fd;
    decBuf[384] = 256'haafdb1fdb8fdb2fd97fd74fd38fdeefcbcfca1fc88fc8ffc89fc82fc7dfc59fc;
    decBuf[385] = 256'h2ffc08fceefbd7fbd3fbcffbcbfbd5fbd2fbd5fbd7fbddfbeffb0efc34fc6dfc;
    decBuf[386] = 256'hb0fcf0fc3afd80fdc0fdfafd2ffe5ffea3fed1fefafe2fff51ff70ff8dffbbff;
    decBuf[387] = 256'hf3ff270065009f00c500cb00d200b600a6008f007a006600550045003d003500;
    decBuf[388] = 256'h320039003b00390027000400cbff88ff48ff0effdafed3fed9fe00ff2eff5aff;
    decBuf[389] = 256'h76ff71ff5aff34fff1feb1fe88fe63fe5cfe6efea1feedfe47ff9cffe9ff1b00;
    decBuf[390] = 256'h36003e0046004d005f009200d0002b017f01e201250231023c02320229022102;
    decBuf[391] = 256'h29023d025c02790288028d028002740271027a028802a502c002d202db02d802;
    decBuf[392] = 256'hc602b10297027e027502780285029602a0029a028002550223020002ee01f301;
    decBuf[393] = 256'h170253028d02b202d502db02e102d102ba02b602c202d30202034e03a8031504;
    decBuf[394] = 256'h5e04870493045c041604c4038d0383039e03d8030c044a0473047b0474045504;
    decBuf[395] = 256'h2d04ff03e003b903a903a503a903c403e303f9031404330440044c0448043204;
    decBuf[396] = 256'h18040004de03d003dc03e80308042e043d04540461046504760486049a04b704;
    decBuf[397] = 256'hd204eb040d0537056905b505fb053b0675068b06920698069306a206cc06f306;
    decBuf[398] = 256'h1707400751074c073e072107f606cf06a00681067c0681068f06a406af069e06;
    decBuf[399] = 256'h7c063f06f505af058205690552053e052b0531052b051e0522051605fe04e804;
    decBuf[400] = 256'hbd049104750465046104650469045e045b04580456047504a304cf0402051605;
    decBuf[401] = 256'h10050b05f104da04e70409054605a005f50542069c06d906e406ee06c0069706;
    decBuf[402] = 256'h80066c067f06b106e1060d0734073a072c0727071c07110714070c07ef06dc06;
    decBuf[403] = 256'hbc06a706ab06ae06b106b406a2067e0665063b061406fa05da05bc05a1057a05;
    decBuf[404] = 256'h6105530557055b056c05630549052a05fb04c304ac048a0477047d0477046004;
    decBuf[405] = 256'h5c0450043f043604270410040604f203e003e703f103fb030b040d0403040204;
    decBuf[406] = 256'hf903f503ff03fb03ec03da03c003a1039c03a803c703ff033304560468045704;
    decBuf[407] = 256'h34041304ed03de03eb0301041c04490469046e047e04700463045f0455045104;
    decBuf[408] = 256'h5a0462046e04810489048b049a04a004a504b704c304c504cb04bf04a7048004;
    decBuf[409] = 256'h52040d04e003b603a003a703ad03be03cd03bf0388034503ce025c021202ea01;
    decBuf[410] = 256'hc601e70105022002390232020102c90186013401fd00df00c300dc00f200f900;
    decBuf[411] = 256'h0c01fb00d700ae007b004b0045003f0044005b00680074007e008e009c00b900;
    decBuf[412] = 256'hd400f4001a0134014b016001730185019b01af01c101d701eb01fd0112022102;
    decBuf[413] = 256'h290222020e02f701e101cd01c001bd01bb01b901bb01b601a9019c018a017501;
    decBuf[414] = 256'h6101490133011f010801f200d200ac00920072005d0051004e003e002400feff;
    decBuf[415] = 256'hc5ff82ff54ff2bff14ff1bff21ff32ff37ff2aff0cffe1febafea0fe89fe7cfe;
    decBuf[416] = 256'h78fe83fe93fea7feb4febbfeb5fea3fe88fe70fe67fe6ffe82fe9cfeb4febefe;
    decBuf[417] = 256'haffe98fe7bfe68fe5efe61fe69fe7cfe91fe9afe9cfe95fe86fe74fe64fe5dfe;
    decBuf[418] = 256'h5ffe76fe98fecbfefbfe1bff37ff3cff25ff10fffcfef2fe08ff33ff5eff86ff;
    decBuf[419] = 256'h9fffa4ff8fff6cff4cff3fff43ff54ff77ff8effa3ff9fff95ff85ff77ff6fff;
    decBuf[420] = 256'h68ff65ff5bff4cff3dff27ff07ffe9fecefea1fe75fe4efe2afe13fe0efe12fe;
    decBuf[421] = 256'h16fe0cfee1fd9dfd4afdfdfccbfcb0fcb8fcedfc0ffd22fd28fd18fdf8fcd2fc;
    decBuf[422] = 256'haefc97fc8afc95fca7fcd0fc02fd32fd5efd7afd7ffd7bfd6efd62fd6dfd8ffd;
    decBuf[423] = 256'hb9fdebfd29fe53fe78fe9afeadfed5feeefe0fff35ff4eff5cff61ff64ff68ff;
    decBuf[424] = 256'h71ff7aff82ff89ff8bff85ff7cff71ff5aff38ff0effdcfeb9fea7fea1fea6fe;
    decBuf[425] = 256'hc7fed3fedffed4feacfe79fe49fe11fefafde6fdecfd08fe22fe30fe2bfe18fe;
    decBuf[426] = 256'he3fdaffd71fd48fd31fd2afd3dfd65fd88fda0fdacfdb0fd9ffd8ffd81fd74fd;
    decBuf[427] = 256'h7bfd8afda0fdbffdddfdf0fdfbfd04fefcfdf9fdf2fdebfdedfdeffdeefdeffd;
    decBuf[428] = 256'heefde0fdd0fdc1fdabfda3fda0fd9efda4fdaafda1fd96fd88fd72fd68fd6bfd;
    decBuf[429] = 256'h7efda1fddafdfffd21fe34fe2ffe1ffe11fefcfd08fe19fe3cfe65fe8dfea6fe;
    decBuf[430] = 256'hb4feb8fea5fe8cfe7dfe7afe8cfeb0fee8fe1dff4dff6cff72ff6dff56ff49ff;
    decBuf[431] = 256'h35ff2bff28ff2bff28ff2aff24ff12fffdfed7fea9fe7dfe56fe47fe42fe4ffe;
    decBuf[432] = 256'h53fe56fe40fe15feddfd99fd6cfd53fd4cfd52fd65fd60fd46fd26fdfffcd1fc;
    decBuf[433] = 256'hbefcaefca8fcb6fcc3fcdefcfefc24fd48fd68fd7dfd81fd7efd81fd95fdbcfd;
    decBuf[434] = 256'hfafd45fe77feb6fecffed7fedefee4fee9fef9fefdfe0aff16ff20ff36ff56ff;
    decBuf[435] = 256'h74ff8fffa7ffa4ff9bff8eff79ff6bff72ff7eff96ffacffc0ffcdffcfffcdff;
    decBuf[436] = 256'hc3ffb0ff8eff64ff31fff4fecafeb4fe9ffea5feabfea6fea1fe8cfe71fe58fe;
    decBuf[437] = 256'h43fe2efe1cfe15fe17fe25fe3cfe5efe7ffea5febefeccfed1fecdfec2feb3fe;
    decBuf[438] = 256'ha4fe9cfe95fe97fea1feb8fecefee8fe07ff14ff10ff06ffeafecefebdfeb4fe;
    decBuf[439] = 256'hc2fedffe02ff2bff47ff57ff52ff3dff22fffbfed7feb7feaafeaefec7fee9fe;
    decBuf[440] = 256'h13ff24ff33ff38ff22ff07fff6fee0feddfeeafe04ff32ff6aff9effc1ffe0ff;
    decBuf[441] = 256'he6ffe1ffd3ffbdffbaffc4ffd4fff3ff11002c003e004d005600590064006f00;
    decBuf[442] = 256'h81008d0098009e009800900083007a007200730077007b007c0071005b002c00;
    decBuf[443] = 256'he0ff9aff48ff11fff3fed8fee0fef7fe19ff2cff26ff0cffe3feb0fe80fe54fe;
    decBuf[444] = 256'h43fe53fe73fea2fedafe00ff07ff0dfffcfee2fed4fed0fee4fe03ff32ff6aff;
    decBuf[445] = 256'h90ffb2ffd1ffccffd1ffd5ffebff0d004a009400da0007012001280121011b01;
    decBuf[446] = 256'h2b0145016f01a101c401e301dd01b90199016a014b012f0120011b011f011b01;
    decBuf[447] = 256'h11010101e700c1009d0073004c003d0038004d00700090009d008a0063002b00;
    decBuf[448] = 256'hf6ffc6ffc0ffc6ffeaff0a001f00230019000300e3ffd6ffd2ffebff1a005800;
    decBuf[449] = 256'h9100c600f600fc000201f300ee00f2000d0134016c01a101d101e401de01c401;
    decBuf[450] = 256'h9b0173015a0143013e01520163017f018b018e0185016b01530137012b012001;
    decBuf[451] = 256'h240126012401260120011e01200128013801470155015a015f015b0154014901;
    decBuf[452] = 256'h38012901230125013d016b01a301e70114021c0224020202e201d101e1010102;
    decBuf[453] = 256'h30027502a202cc02e202db02c802b8029e0287027a0267025c025f025c026402;
    decBuf[454] = 256'h6b0261024f022b02fd01c5019f017d016a0165015f015b015701430132012201;
    decBuf[455] = 256'h0e010101f500ef00ed00eb00f000fa0009011f013901590176019201aa01ba01;
    decBuf[456] = 256'hc801d501dc01e301ed01f201fa0105021102230242025f027b0293029c029f02;
    decBuf[457] = 256'h97028c0285029302aa02cc02f6021d0337034e034a033e031f03e702b3027502;
    decBuf[458] = 256'h3b021602010214021a021f020802d90188012501e200a50084008e0097009f00;
    decBuf[459] = 256'ha700bc00c200de00f8000f0113010f010501f500f200fa000b0126013a013d01;
    decBuf[460] = 256'h3a012c012e013a0151016e0189018c018901860184019401b401f0012a025e02;
    decBuf[461] = 256'h810287028d02730265025802550258025b02640266025f0248022602f301b501;
    decBuf[462] = 256'h7b0138010a01e100d900d200d900c800ae00840052002f001000fffffaff0800;
    decBuf[463] = 256'h1500200032003b003e0046004d0054006200710084009700ac00bb00cd00d900;
    decBuf[464] = 256'he300e900f6000801260144016f019601b001c701d401d001c501bc01b301b101;
    decBuf[465] = 256'hb801c201c801c301ab018401600137011b010b01fd00f100dd00c500a2008200;
    decBuf[466] = 256'h5c0042002b000d00faffe8ffd9ffc5ffbdffb6ffafffadffa8ffa3ffa2ffa3ff;
    decBuf[467] = 256'hacffbdffd2ffecff0b0021003c00540064007e008f00a500b900d100da00e900;
    decBuf[468] = 256'hfb0002011101230134014701590160016701610154013f012b010e01fb00e900;
    decBuf[469] = 256'hda00cb00c400b800a50088005d003600fdffc9ffa6ff87ff76ff5dff4fff3aff;
    decBuf[470] = 256'h26ff1cff0cff09ff07ff04fffefef8feecfee3fee8fef7fe11ff31ff4eff69ff;
    decBuf[471] = 256'h7bff84ff98ffabffbbffd3ffe9fff7ff040010001b003100500077009a00bb00;
    decBuf[472] = 256'hd000dc00df00e200e500ed00f900ff0005010401fb00f100df00ce00b7009b00;
    decBuf[473] = 256'h780045001500ddffa8ff78ff59ff32ff18fff8fedafeb7fe97fe81fe66fe55fe;
    decBuf[474] = 256'h4bfe43fe45fe51fe64fe86fea7fecdfef1fefffe0cff0fff05ff02fff9fefcfe;
    decBuf[475] = 256'hfefe09ff17ff27ff3aff51ff61ff75ff82ff85ff87ff85ff7fff81ff89ff95ff;
    decBuf[476] = 256'hadffd4fff8ff210032004200460039001e000600e3ffbaff92ff6fff45ff29ff;
    decBuf[477] = 256'h19ff0cff07ff03fff9fef0fedbfecefec7fecefee0fefefe1cff30ff3aff3dff;
    decBuf[478] = 256'h3aff2dff26ff1bff15ff14ff0cff0dff09ff05ff02fffbfeeefed4feb4fe8efe;
    decBuf[479] = 256'h60fe41fe24fe15fe1afe2ffe4afe6afe7ffe92fe9dfea6fea9fea6fea4fe9efe;
    decBuf[480] = 256'h94fe8bfe86fe84fe8bfe9cfeb7fed2fef9fe1dff34ff52ff5dff68ff6bff6eff;
    decBuf[481] = 256'h70ff81ff90ffa6ffbaffd2ffdbffe9ffe7ffe4ffdeffd0ffb6ff9bff74ff50ff;
    decBuf[482] = 256'h27fff4fec4fe98fe65fe35fe0afeedfdcafdb2fda6fd9afd90fd80fd77fd7afd;
    decBuf[483] = 256'h7cfd87fd99fdaafdb4fdb6fdb1fda9fd9efd95fd93fd99fda8fdbffde2fd0bfe;
    decBuf[484] = 256'h3efe6efe9afec1fed1fed5fed1febefeb3feaafeb2fec5fedffefefe1cff28ff;
    decBuf[485] = 256'h32ff2fff21ff09ffe7feb4fe84fe3ffefffdc5fd82fd54fd2bfd06fdf1fcdefc;
    decBuf[486] = 256'hc2fcbdfca6fc99fc7efc6cfc50fc35fc16fc00fcedfbeafbf9fb19fc50fc94fc;
    decBuf[487] = 256'he6fc49fda6fdfbfd48fe8efecefef7fe0eff15ff0efffefeeefee0fee5fe00ff;
    decBuf[488] = 256'h26ff5fff84ffa6ffadff9cff6eff35fff2fea0fe69fe23fee3fdbafd94fd80fd;
    decBuf[489] = 256'h6dfd67fd58fd37fd09fdd0fc8dfc5ffc26fc00fcebfbd9fbbdfb99fb6ffb3cfb;
    decBuf[490] = 256'h0cfbe1fad0fadffaf6fa2dfb71fbb1fbfbfb2dfc5bfc84fca9fcbefcddfc10fd;
    decBuf[491] = 256'h4efd98fd06fe6dfecbfe08ff3fff5dff53ff2aff05ffc7fe8dfe4afe1cfef3fd;
    decBuf[492] = 256'hcdfdabfd98fd87fd78fd6afd4cfd31fd0bfde7fcc6fcbafcbdfccffcf8fc1ffd;
    decBuf[493] = 256'h39fd50fd43fd28fd01fdc9fc94fc64fc45fc29fc1afc1efc33fc4ffc6efc8cfc;
    decBuf[494] = 256'h97fc94fc78fc4dfc26fc0cfc08fc2efc70fcc3fc26fd83fdc0fdf7fd15fe30fe;
    decBuf[495] = 256'h38fe40fe39fe33fe2dfe1efe19fe15fe19fe23fe39fe53fe6cfe81fe96feadfe;
    decBuf[496] = 256'hc9fee4fef6fefffefcfeeafed5fec1febefec5fee1fe04ff24ff31ff35ff31ff;
    decBuf[497] = 256'h2eff37ff59ff95ffdfff39008e00c500e300fe0017013d018801ce0133027502;
    decBuf[498] = 256'h9a02a50287026b0253022d02190212020d02fd01ef01e301e701f1010d022802;
    decBuf[499] = 256'h410244024102390237024a027102c6021b037e03db031804390443041504cb03;
    decBuf[500] = 256'h71030403ba0277023b021a02fc01e001b7018201520127011601fc00e500bf00;
    decBuf[501] = 256'h7200f9ff67ffddfe84fe53fe62fe8afeaefecffed9fed0fea7fe72fe5efe58fe;
    decBuf[502] = 256'h52fe57fe49fe34fe19fe0efe24fe4ffeadfe76ff3f00c2003801a40107023c02;
    decBuf[503] = 256'h6d02b702df0203030e03dc029c0252020c02f10109023e02a5020c034f038c03;
    decBuf[504] = 256'h810363032303e902b502920273026d025e0250025d028002c5023303b8035904;
    decBuf[505] = 256'hc5040005ee04bd043804bb034a03e202850260023f02490265028e02e0022d03;
    decBuf[506] = 256'h8703f5033e044c0458044d042f0426041d044304580477049e04ae04bb04d104;
    decBuf[507] = 256'hdc04d904e804d404b70495044f04cd0350039d02c801380181003a0024005f00;
    decBuf[508] = 256'h0001ee01cb020704da044d05b605d505b9056a0552051205fe04ec04dc040805;
    decBuf[509] = 256'h30058505fe0590061a07bb075208b408ea08d908cb08a3087e083108ff07ad07;
    decBuf[510] = 256'h60070607c90692069c06ef0668071a08c10801093c09e3085108790776063c05;
    decBuf[511] = 256'h150409035a02bc019f01ba0160022203d90350043a04d803cc0226012dff51fd;
    decBuf[512] = 256'haafae5f84af73ff573f4b9f3a1f2a2f117f1f0ef16f07ff09bf1dbf3bff678f9;
    decBuf[513] = 256'ha6fceffd52feadfefffe4aff2601cd036608c70c0b13e018aa1c7d21df25b728;
    decBuf[514] = 256'h4e2bb72c492c1f2b5a29bf2774274028e82a802f6336ce3ca4427649364c0b4d;
    decBuf[515] = 256'h494cd8483543633c4d32e8285d206116ab0f2007940189fcc9f9f3f321ede0e4;
    decBuf[516] = 256'he4dad0ce71c327b637add8a16a9d63992b9847994e9cb9a28ea8e4b0a8b8bdc1;
    decBuf[517] = 256'h47cad3cfe3d64edd79e1c7e69aeb7df2e8f813029e0ad216f11e4729ac32373b;
    decBuf[518] = 256'hc340ca43b444df439941c63c2437523011284d203e19d212fd0c33096004feff;
    decBuf[519] = 256'hdffa4bf33bec25e210d6b1ca5bc0f5b6faab98a4339b8a9736943393f4951e9a;
    decBuf[520] = 256'he89dbba21da719aba7ac10aea2ad06ae60aefbaf9cb280b631bc03c36ec99ad2;
    decBuf[521] = 256'h24dbe8e2f8e963f039f687fb98fd79ff2e01b2013a018302ad037205b107bd09;
    decBuf[522] = 256'h990bcd0c050d060c650a8b07450325fef2f771f05de7d3ded7d471cbe7c2ebb8;
    decBuf[523] = 256'he4b4caaeaeada7aa92abbcaa7eabceaa2eaa79a8eba673a6e0a60ba839ab13af;
    decBuf[524] = 256'hcdb538bc64c55fd0b5da1ae416ef78f62efd48039c06a209630c380d7e0f8f11;
    decBuf[525] = 256'h2f12c1124613ec10c80e100ce108080568012dfd0df8daf159ea45e1bbd8bfce;
    decBuf[526] = 256'h59c5cfbc43b733b09dab1da9d7a627a607a8bda94aaba4ad11ae75aecfaed9ad;
    decBuf[527] = 256'hf8acb4ace9ade2af56b382b855bdb7c1b3c541c7b9c726c835c625c5d3c41ec5;
    decBuf[528] = 256'h72c610cab0cddcd270da80e1c0e984f190f6d0fe9406a90fa41aee2771340f43;
    decBuf[529] = 256'hd250e860b76b8b75e87ac87f4e7e477a0e7982737c70bb6d3b6bf5682364405d;
    decBuf[530] = 256'h2a53154736359024c80c9ef679e229d0c1ba5dac84a4619de596dc981297b298;
    decBuf[531] = 256'h209d789e21a275a585acc6b4c2be85cd48db5eeb80fa4308eb1b0029a639c948;
    decBuf[532] = 256'h8c560e632d6b8f724679ef7c0b7e0d7f4d7c22785874246e4f6801636d5b5d54;
    decBuf[533] = 256'h1c4c5844443b4930f325de197f0e290414f8f5ef93e8dde1c3dba7daa5d98fda;
    decBuf[534] = 256'h65db2fdf40e1a2e57ae811eb5bee7ff070f2eaf42af735f911fbc1fcbafe9600;
    decBuf[535] = 256'hc202380414064907f107be073307b8058703e6006cfe88fbd0f80bf770f5bbf5;
    decBuf[536] = 256'h87f6b2f8e9fbc2ff6b048c07880b280f8211a513d014df15d6164c18a019cb1b;
    decBuf[537] = 256'h6c1ee62025233125fd253a26922561232b20761bd415020fc106fdfee9f55eed;
    decBuf[538] = 256'h9ae58fe024daf9d52fd21ed0fdcc47cbb1c838c8cbc72ec83ec97ecb1ece02d2;
    decBuf[539] = 256'haad64ddc1fe38ae90af11ffaa9026d0a7d11be194a1f5524eb28162d5c2f6d31;
    decBuf[540] = 256'h4d33df335b33e2329a31a82fe42d002b472819253f21a01d64194414720f100b;
    decBuf[541] = 256'hcd04a20054fbe2f701f629f3a4f23bf1cdf031f1d6f0cdf118f25cf215f3ddf2;
    decBuf[542] = 256'h10f33ef369f328f4a8f5d9f77afaa8fda7005f038e06b1086a0be30d23102e12;
    decBuf[543] = 256'h1a15d3174c1a8c1c971eeb1f2021c821c722af232e243a25a32502261f266825;
    decBuf[544] = 256'h33240f226f1f401c6718be135c0f3d0a6a0508010cfd63f842f569f2d3ef88ec;
    decBuf[545] = 256'h8ae90ae6c0e2e6de47dbedd8a4d741d79bd792d808dae4db10deb0e02ae30ee6;
    decBuf[546] = 256'hc7e8aaec4af0a3f27df613f96dfb91fd82ff470187039205e60696083e09d709;
    decBuf[547] = 256'h060adc091c0928080b071805b402d0ff17fde9f9eaf66bf311f1c9ef9eeedaec;
    decBuf[548] = 256'he3eb03eb27e9f2e7f9e51de46ce273e01fdf6fdd56dcf1da0ada8bd965d988d9;
    decBuf[549] = 256'h26dab6daa1db00dc8fdca9dcc1dcacdce6dc1cddcfddd4de0ee089e154e304e5;
    decBuf[550] = 256'h8de6bee8c9ea2ded6def0ef287f4c7f63df891f9c6fa6efba1fbcffba5fb32fb;
    decBuf[551] = 256'hcafa2bfa62f977f85af74ef6cef403f3d7f0a1eda3ea5ce660e2c0de76db9cd7;
    decBuf[552] = 256'h06d5acd23ed214d1b9d00cd1ecd1b8d2edd376d5dbd6d9d82dda58dc64de40e0;
    decBuf[553] = 256'h6be20ce53be814ecb4efeff3ebf782faccfdcb00bc02cc03c3040d05c9049503;
    decBuf[554] = 256'h0c0275fffbfc17fa5ff730f40df28dee33ec5ae8c3e588e18cddecd9a1d6c8d2;
    decBuf[555] = 256'h28cfcfcc86cb5cca01ca53ca34cb88ccb3ce29d005d2b5d33ed5a3d68bd706d9;
    decBuf[556] = 256'h6bdab0db7fddabdf21e1ede121e3e9e2b6e22be204e1abdf20dfa1de15df4ee0;
    decBuf[557] = 256'h1ee24ae480e77eea70ece9ee29f19ff203f5e7f72efc9403a90ca417ee240335;
    decBuf[558] = 256'h2644e9516b5eca69386e906fc870746d6968d363a85f5a5ae956c753a84ed549;
    decBuf[559] = 256'hb241b637a12bc2191c09a7f557e3b0d28ec3bab9cab02aafa4b0fcb116b86abb;
    decBuf[560] = 256'h7ac2e5c8bace08d49ddbb1e43bed6ff9cf04250fe81dab2b9b343a43fc50ec59;
    decBuf[561] = 256'h4b65a16f5776717c8d7d8f7ea47d7a792c74f86d7866685f2757634f5448e841;
    decBuf[562] = 256'h133c4135d52e00292e22ed192912190bae04d8fe8af919f638f4a6f334f59df6;
    decBuf[563] = 256'hc0f840fc9afe980151041506b0079108d508a007f7062c0501038b01affffffd;
    decBuf[564] = 256'h56fdbdfc32fc5cfc83fc60fc7ffc9cfc4efca8fb10fb60fae9f9fef9affa13fc;
    decBuf[565] = 256'h10ffc5036709b50ee8141319611e34231525ca265728d0286228382728263225;
    decBuf[566] = 256'h51248523cc22b321b420b61e521cca189d13cb0ee807a7ff1bfa07f1edea61e5;
    decBuf[567] = 256'h56e096dd6bd9a9d8f8d799d82ad9c1db1bde19e160e539e8e1ec43f13ff5dff8;
    decBuf[568] = 256'h0bfedd023f075f0c92126818321c042166256229f92b622df52c912c182a3327;
    decBuf[569] = 256'hb423781f7c1bdd1792146f12b60ff20d560ce10a8d095808cf066a05c9034002;
    decBuf[570] = 256'ha7011c019a01a70226045706f808710b560e0e1188132315031647168e15e614;
    decBuf[571] = 256'he7134512bc10f10e410db80b530ab20899070007d206a8061b07c9072808f108;
    decBuf[572] = 256'h74091a0add0afc0b560df70ef010cc12f81403176719a71b481e0c200321e321;
    decBuf[573] = 256'h9f216a20011e1d1bd616da12310e100b140774032a002bfdacf961f663f3aaf0;
    decBuf[574] = 256'h7ced7deafee6a4e45be331e2d6e1cde243e4a7e68be90bed64ef63f21bf5e0f6;
    decBuf[575] = 256'h20f92bfb8ffd2aff35018902be0367040005d10453049303e502c8016f002aff;
    decBuf[576] = 256'h5bfdaafb41f901f760f432f10eef56ecdce941e836e65ae425e30de274e145e1;
    decBuf[577] = 256'h6fe1e2e191e2f0e27fe39ae3e1e322e484e401e5b4e52ae6c2e6fde60fe7fee6;
    decBuf[578] = 256'hd2e674e638e617e695e518e544e408e38de18ee049dfcbdef1de5adf77e0d0e1;
    decBuf[579] = 256'h15e33ce495e57de6f8e7c3e973eb6cedd0ef6cf177f3cbf400f618f7b1f73cf8;
    decBuf[580] = 256'hbbf82ef9c5f866f89df77ef624f583f3faf1c9efbeede2eb3be9c1e681e476e2;
    decBuf[581] = 256'h9ae0eaded1dd38dd50dcd2dbf8db1bdc7adcb6dd31dffce028e3c9e542e827eb;
    decBuf[582] = 256'h18ed92ef2df1a3f2f7f32bf5b4f619f817fa6bfb1cfd34fecdfe58ffdafe1afe;
    decBuf[583] = 256'he0fc11fbe5f844f6cbf342f0e8edeaeaf8e8e9e7f2e612e646e58de474e375e2;
    decBuf[584] = 256'heae16be1f8e0d5e034e151e19fe116e282e233e368e48fe535e7bee8bde948ea;
    decBuf[585] = 256'h1eea5ee9dee713e663e4f9e1badfaeddd2db22da0ad90bd87fd7fed7bed8f8d9;
    decBuf[586] = 256'h73db3edd72defbdf60e148e2c3e3f4e595e8e3edb5f4f5fc29098814c624e933;
    decBuf[587] = 256'hac41c151915c7662d3677369f967f263d85d4c583c51a74c7c48b244df3f3d3a;
    decBuf[588] = 256'he731eb272719640bbcf76be5c5d4a3c5cfbbdfb2ffad85acddadf7b383b993c0;
    decBuf[589] = 256'hd3c85fce6fd5dadbb0e182e8c3f087f8a003f60d0a1a6925bf2fd43b33478951;
    decBuf[590] = 256'hee5a08619466a06b8a6c0a6a40660d60375ae1511d4a0941ef3a6335532ebe29;
    decBuf[591] = 256'h9325c921571ef519d5140310600a9606c401a3fecafb3cfac4f90cfbfefc77ff;
    decBuf[592] = 256'hb7015804d1066d08b708fb08c7075d051e0352ffa9fa48f64bf2a3ed82ea85e6;
    decBuf[593] = 256'hf8e48fe321e34ce410e6abe7b7e993eb43edccee31f0d2f1cbf32ff6b8f9f3fd;
    decBuf[594] = 256'h13034709c710d7176c1c42229027022ba22b342ca62a5c278223da1e781a7c16;
    decBuf[595] = 256'hdc12920fb80b1908ce04f50055fd29f856f3b4ed66e833e25ddc0fd73cd21bcf;
    decBuf[596] = 256'h42ccbecb36cc5ace12d1f6d495d8c1dd94e236e800ecd3f0f4f3f0f787fad2fd;
    decBuf[597] = 256'hf5ffae022705b008fa0baf101115541b7f1fcd243f281f2ab12a2429ca26f022;
    decBuf[598] = 256'h511f151b19177a132011fc0ed20dc20ccc0b810bb50a05097c07e504b601ddfd;
    decBuf[599] = 256'h3dfae3f7c0f55cf5b7f5f7f72dfb2bfeab01050428061a087408c6087c08b007;
    decBuf[600] = 256'h7b06f204270377015e002b00130137036d06460ae60d31112f14e816ac18ec1a;
    decBuf[601] = 256'h621cb61dea1e73207221fd21d022dd23d124ed25fa267a281329e4286927d224;
    decBuf[602] = 256'hef203d1bef15bc0fe6099804c5ff64fb67f7c8f36ef14bef59ed4aec53eb73ea;
    decBuf[603] = 256'ha7e972e8e9e684e53fe415e4d5e4e0e616eaf0ed98f2faf6f6fa96fed102aa05;
    decBuf[604] = 256'h41089a0abe0ce80df80e010e210dcd0b980a0f0910088507b3063f0606053603;
    decBuf[605] = 256'h8f0015fe8dfa42f744f48bf15dee39ec81e9bce77ce59ce4d0e389e432e5fde6;
    decBuf[606] = 256'h31e8bae953ea82ea03eaf7e803e8e6e673e6c4e526e5d0e44de4a7e366e353e3;
    decBuf[607] = 256'h88e33be4e1e4a4e5f2e57ce562e409e368e14fe01ce004e1d3e2ffe435e834eb;
    decBuf[608] = 256'h25ed9fef3af145f399f4cef576f60ff7e1f663f6a3f53af5dbf4bff40df584f5;
    decBuf[609] = 256'hc5f58af5e9f4a4f3a6f1caef9fed93eb2fe994e71ee642e40ee385e186e0fbdf;
    decBuf[610] = 256'h25e0e5e064e22fe45be666e8caea0aed80ee5cf00cf225f38af4cef5f5f602f8;
    decBuf[611] = 256'hf6f8d3f9d6fa10fce2fca2fd51fe31fedbfdf0fc55fbccf901f8d5f55ff493f3;
    decBuf[612] = 256'hdaf232f2fff173f1f5f082f08eef2fefd9ee56ee3eee29eeeeed71edffec7aec;
    decBuf[613] = 256'hd9eb6deb0bebd5ea06eb6debe6eb78ec50ede0ed2eee46eeaeedafec30eb65e9;
    decBuf[614] = 256'hbde6f9e4b9e218e054de5ddd7ddcb1db73dbcbdafeda2cdb02db75dbafdcd6dd;
    decBuf[615] = 256'hc9dfb5e234e67fe958edf8f033f577fb4c01260b3b179a22d832fa41ac53905f;
    decBuf[616] = 256'h606a3474fd755d74e3722d6ca363175e07579c50c64afc462942473bdb34062a;
    decBuf[617] = 256'hbc1ca60c84fdd2eb2cdb0acc47be57b5b8b332b5e8bb02c2c6c9dad264db28e3;
    decBuf[618] = 256'h38eaa3f079f64bfd8c05500d6416ef1eeb28ff341f3d694a5853785bce65846c;
    decBuf[619] = 256'h2d7049714b728b6fb5696764d35cbf53344b7043603ccb37f5312b2e1a2c392a;
    decBuf[620] = 256'h8428ed259423ba1f1b1cdf17e3134310da0e920dbc0ecc0f67117213c6148015;
    decBuf[621] = 256'hb8151f15da135f122e10620cc3089703c4fe22f950f2baed8fe9c5e515e574e4;
    decBuf[622] = 256'h2ae6c0e80becbff021f541fa13ff75037107110b5c0e5a111314f6179f1c4122;
    decBuf[623] = 256'h8f27c22d98336237d43a743be23a43370733e82d152932229c1dc7177912a60d;
    decBuf[624] = 256'h04083a0467ff46fc4af8aaf460f186ede7e99ce6c3e22ce0e1dc99db6eda14da;
    decBuf[625] = 256'h0bdb80dce4de6de2a9e6c8ebfcf127f675fb47002802dd036b05f2048504e804;
    decBuf[626] = 256'h43053a06af078b093c0ba50de50f5a11261264124c11810fd90cab09ac06bb04;
    decBuf[627] = 256'h4102ef01a4017002a5032e059306d807a709570be00cab0ed7104d121913d213;
    decBuf[628] = 256'h0a143d14c8144615a016e41760195f1a8d1aba19611863167713f70fad0cd308;
    decBuf[629] = 256'h2b04c9ffa9fad7f5b5f200f17cf0e5f12df31ff5e3f67ef88afadefb09fe1500;
    decBuf[630] = 256'h01038006cb09c90c4910a312a1159317c11ae51c6420be22e2240c26fd246123;
    decBuf[631] = 256'h2b20521cb21877149e11fe0da50b8109900716057b030502b100f8ff4fffeafd;
    decBuf[632] = 256'hecfb88f9a4f6ecf327f230f111f265f390f59cf778f931faf9f960f91bf8a0f6;
    decBuf[633] = 256'h3bf5f6f3cff229f130efccec8ceaece727e68ce4ace3f0e32de466e499e46ae4;
    decBuf[634] = 256'h94e407e5fce557e756e9baeb55ed60efb4f0e9f101f366f465f6c9f8adfb9efd;
    decBuf[635] = 256'h18006a001f0043fe9cfb6ef894f4f5f0aaedabeaf3e7c4e4c6e146defcdafdd7;
    decBuf[636] = 256'h45d580d38ad2a9d1ddd024d00bcf72ce44ce17cf0ad1f6d375d7b0dbaddf43e2;
    decBuf[637] = 256'h8ee58ce87eeaf7ec37ef42f196f2cbf393f3faf259f1d0ef6bee83edb0ec8aec;
    decBuf[638] = 256'h67ecc9ebc6ea46e97be750e544e368e1afe007e06edf3fdf15dfefdeccde2bdf;
    decBuf[639] = 256'hf4df14e1bae2b3e48fe63fe858e9f1e91fea49ea70ea92eab2eacfeab5ea3eea;
    decBuf[640] = 256'h7be9c4e8bfe711e7b2e622e608e6c1e5fee413e436e3c0e1c1e036e060e020e1;
    decBuf[641] = 256'h9fe26ae41be6a4e709e94deac8eb2ded72eeedef52f1ddf107f247f1c8effded;
    decBuf[642] = 256'h4dec53eaffe846e82ee795e6ade586e493e22fe04bddcbd990d5b7d20fceedca;
    decBuf[643] = 256'h15c87ec524c3dcc178c11ec170c150c2a4c3d9c462c6c7c7c5c929ccb2cfedd3;
    decBuf[644] = 256'h0dd940df16e56cedf8f20cfc9704930ea71a462909371e47415615600569e46d;
    decBuf[645] = 256'h5e6f576bae67ea5fd6564b4e8746783f0c398c317c2a3c2240182b0c8cfdc9ef;
    decBuf[646] = 256'hb4df91d0cfc24cb62daebfa967a810acd4b3e8bc73c56fcfd4d85fe123e937f2;
    decBuf[647] = 256'h51f84d02b30b3d14011c1525a02d6435743cdf425f4a6f510556305afa5daa5e;
    decBuf[648] = 256'hc95cf1593f546d4d0247823f6d365330c72abc25fc22272265211522f6236423;
    decBuf[649] = 256'hd6217d1fa31b0418c813cc0f3e0ed50c430da60d4c0dfa0c840b20093c06bc02;
    decBuf[650] = 256'h81fe84fadcf57af15aec88e7e6e198dc26d9c4d4ebd167d1dfd103d482d7aedc;
    decBuf[651] = 256'he2e262ea72f1b2f976018608f10e1c13e616581a791d762115255129702ee231;
    decBuf[652] = 256'h033595351135c631122d6f279d20321ab212a20b370561ff13faa1f63ff243ee;
    decBuf[653] = 256'ha4ea4ae826e635e470e2d5e05fdf0bde52ddaadcdddcc5ddebde92e08be2efe4;
    decBuf[654] = 256'hd3e752eb9dee52f3b3f7b0fb4fffa901f1025503fa025f017f00b3ff75ff8e00;
    decBuf[655] = 256'hf3014e043207ea09640ca40eaf10031238137013a313d113a713cd137c14d815;
    decBuf[656] = 256'h3318171b961ed222aa253827c0267725bf22db1e331a111715137f10340d100b;
    decBuf[657] = 256'h1f095a0764068305b7047a04d103d2023101a8ff77fd01fcadfaebfa74fc0bff;
    decBuf[658] = 256'hee028e06c90ac60e6512b0158919201c6a1f4423da2543278c28ef28e027e926;
    decBuf[659] = 256'h09263d2584244c24b323cb2250211f1f7e1c4f195116d112870f880c0909be05;
    decBuf[660] = 256'hc00207008efd97fce2fc36fee6ff4f02ea0360052c06ee05b6051d0535040b04;
    decBuf[661] = 256'he503c203e203c50377035f0349038403010473046404b6035202bbff8dfc8ef9;
    decBuf[662] = 256'hd6f611f51af4d0f314f451f46af569f651f7ccf831fa19fb94fc93fdc1fd97fd;
    decBuf[663] = 256'hd7fc58fb59fa14f941f81bf8f8f718f835f8b2f77df6aef4fef294f054eedfec;
    decBuf[664] = 256'h8beb56eacde868e7c7e5cee37ae2c0e188e121e266e3e1e446e62ee755e815e9;
    decBuf[665] = 256'hc3e9e0eaeceb6cedd1eeb9efe0f0ecf1e0f23cf4def5d7f73bfa7afcf0fd44ff;
    decBuf[666] = 256'h06ffeefd23fc7cf902f7c2f44df381f243f20bf2d8f1a9f1d7f064f0fbef9cef;
    decBuf[667] = 256'hb9ef07f04ef039f0feef5deff1eeb6eeeceedfef19f1e9f299f4b2f5b1f63cf7;
    decBuf[668] = 256'hbaf72df8dcf8b9f9bcfab0fb0ffcf2fba4fbfdfa91fa2ffa88fa3bfb40fc35fd;
    decBuf[669] = 256'h12fe68fe4efea8fd8ffccffbdbfafdf96ef9ebf845f8d9f74ff71af76bf7d2f7;
    decBuf[670] = 256'h80f856f9acf9c6f9aef9c0f8e3f7e0f632f6d3f5b6f5d0f5e8f5d3f549f585f4;
    decBuf[671] = 256'h65f30cf2c7f0a0efe0ee78ee19eefced7aed74ec3aeb14eabae8d2e754e747e6;
    decBuf[672] = 256'hdfe541e504e4dde21ee2e4e065e03fe0d6dff6df4ce032e04ae0b6e067e16ce2;
    decBuf[673] = 256'h31e4d8e652e9dbec16f112f5bbf99e00de08da12ef1e8e2d513bd34772564660;
    decBuf[674] = 256'h3669d66a506c4968a064145f04589951c34b75464240c138b1317129751f6013;
    decBuf[675] = 256'hc104fef6e9e619dc57ce67c588c00ebf65c07fc60bcc1fd5aadd6ee57eecbef4;
    decBuf[676] = 256'h4afa5a019b09270f3b18551e1926292d9433bf37913e2743fc484a4ebc511e56;
    decBuf[677] = 256'hd3575858ef56cb548550654b9246af3f44391935cb2f592c3829a6282b29a329;
    decBuf[678] = 256'h112a742a652925278424a1200a1ec01ac117d0150b1470126510010e780a2d07;
    decBuf[679] = 256'h790217fe1bfa72f511f114ed6ce80ae40ee06edc24d900d79dd6f7d6dbd95bdd;
    decBuf[680] = 256'h87e2bae83bf04bf78bff87093d10c818541e5f232026a028e62af72cd82eb031;
    decBuf[681] = 256'h3e33a73439340f339530c42b9025101e00179510150909049efdc8f7fef38df0;
    decBuf[682] = 256'h6bed93ea0eeaa5e812e976e9d0e923ea6deab1ea6beb13ec12ed57eed2efd1f0;
    decBuf[683] = 256'h5cf1daf101f224f2c2f28bf3aaf450f6d9f73ef926fa50fa2afa36f9d7f881f8;
    decBuf[684] = 256'h9bf8d0f99ffbcbfd6b009a03bd053d09880c860f0613501674189e19f919a619;
    decBuf[685] = 256'h5c19181955198e198d1ad11ba41cca1c1c1c411add1755140a11310d91095605;
    decBuf[686] = 256'h5901bafd7ff9a6f606f3acf089ee5eed04ed56eda1ed6deea2efbaf01ff21df4;
    decBuf[687] = 256'h81f60afa55fd2e01d705f808f40c9d11be14ba18511b9b1ebf20e92144224d21;
    decBuf[688] = 256'hac1e331caa186f147310dc0d910a9307da041603d600cbfeeffc3ffbb6f951f8;
    decBuf[689] = 256'h0cf791f52cf4e7f215f255f178f116f252f3cdf498f6cdf775f8a8f87af850f8;
    decBuf[690] = 256'hddf774f7d6f60df622f505f45ff2d6f00bef5bedd2ebd3ea48eac9e9f0e913ea;
    decBuf[691] = 256'hf3e910eac1e9aae9bfe9d3e950ea44eb7eeca5edfeee43f069f1c3f2abf37df4;
    decBuf[692] = 256'hf0f413f575f439f315f175eefbeb17e95ee69ae45ae24fe073de47dca6d9e2d7;
    decBuf[693] = 256'ha2d597d343d28ad1e1d048d0bdcf3fcf65cf42cfa1cfa4d0ded1add3d9d5e4d7;
    decBuf[694] = 256'hc0d970dbf9dcf8dd9adfb2e0b1e1f6e274e3e7e3c4e366e30fe3f5e20de379e3;
    decBuf[695] = 256'h78e427e5c5e58ee6dce6f4e635e721e733e764e755e748e723e77ee679e585e4;
    decBuf[696] = 256'h29e3e5e112e105e011dfb2de23dea0dd59dd18dd04dd5eddcfdd8fdeaedfbbe0;
    decBuf[697] = 256'hafe18de21ce3d3e3d8e4cde568e761e93deb69ed74efc8f078f291f32af458f4;
    decBuf[698] = 256'h2ef421f32df2d1f08def12ee13ed2becaceb86eb1debfeeae1ea93ea4beadfe9;
    decBuf[699] = 256'h07e93ee887e7b1e622e6d3e5ebe582e682e7bbe88beab7ecc2ee9ef04ef267f3;
    decBuf[700] = 256'h9af3c8f3f5f2e9f1aff034efcfed2deca5ea40e9fbe7d4e67be536e40fe369e1;
    decBuf[701] = 256'h70df0cddccda2bd8b2d572d3fcd130d16ed117d27cd3d6d516d8b7da30dd15e0;
    decBuf[702] = 256'h06e235e533e825ea53ed52f098f494f84fffba059010e61afb269a355c434c4c;
    decBuf[703] = 256'h6b54d958e05ca85b1c561051a54ad044fe3d9237bd316f2c3b26662094195311;
    decBuf[704] = 256'h570742fbe3ef99e217d6f7cd95c68ec256c1aac4b1c7f2cfb6d7c5de31e5b1ec;
    decBuf[705] = 256'hbcf127f8fdfd4b037e09540fa2147519171f65243829992db9328c37ed3b0d41;
    decBuf[706] = 256'he0450149b64a444ccb4b834a0347c842cc3e1a395035de31bd2e082d832cfc2c;
    decBuf[707] = 256'h442ea82e022f0c2e2b2dc72a3f27f4233f1fde1ae1163912d70ddb093205d100;
    decBuf[708] = 256'hd4fc2cf8caf3f1f05bee01ecdee925e7ace410e305e1b1dff8de30df2fe0e7e2;
    decBuf[709] = 256'hf4e7c7eceaf4aefcc2054d0e4918ff1e19256d28742b5e2c342df62d452da52c;
    decBuf[710] = 256'h132c8f2b162bce29dc2763257f22ff1ec41ac8162813dd0fdf0c260aad071206;
    decBuf[711] = 256'h9c04d0039203ca0363044b0572067f07730811092e09430826073305cf028f00;
    decBuf[712] = 256'h59fd5bfadbf681f483f191ef82ee8bedd6eda2eedfee88efbbef8cef62efd5ef;
    decBuf[713] = 256'h84f01ff2f9f478f8a4fd3805480c5e16c41f4e2812302237b83be33fa540f43f;
    decBuf[714] = 256'h143e3b3ba4385a355b32a32f292de92a74299827f0240d21641c0318e312100e;
    decBuf[715] = 256'hef0a1608890610067e06a807b808530ac90ba50d5e0e770faa0f7b0fa90ee90d;
    decBuf[716] = 256'h690c040bc0094508e0069b05740401046a044705f606190a170d9710e213e016;
    decBuf[717] = 256'h99195d1baf1bfa1b3e1c001ca91c421d861e56200622ff23db251027b827eb27;
    decBuf[718] = 256'h03278825bd239121f11ec21bc4184415fa11200e8a0b3f086504cf0184fe61fc;
    decBuf[719] = 256'h6ffaabf810f79af5cef490f4e8f3b5f3cdf2a6f1e6f038f097f099f1a4f345f6;
    decBuf[720] = 256'hbff8a3fb94fd59ff50009a00ceff15fffdfdfefc16fc43fb1dfb40fbdefb6dfc;
    decBuf[721] = 256'hf0fc67fd51fd3efd08fdd7fc70fc48fcf3fb90fb4dfbf8fa95fa38fab2f9a6f8;
    decBuf[722] = 256'h00f707f5a3f263f0c2ed49ebaee90de748e509e368e0eedd0adb19d909d8b7d7;
    decBuf[723] = 256'h02d8ced87eda77dcdbde1be1bbe380e5c0e7cbe91feb4bedc0ee24f164f305f6;
    decBuf[724] = 256'h7ef863fb54fd19ffb400ff00bb00010079fe14fd72fbe9f984f840f719f6bff4;
    decBuf[725] = 256'h1ef395f130f0ecee70ed0bec24eba8e9a9e865e792e6d2e56ae54ae567e51ee6;
    decBuf[726] = 256'hf3e6f6e730e9abeaaaebefec16ee22ef5cf083f143f2acf2cbf2aef2f8f122f1;
    decBuf[727] = 256'h59f0d6ef5fef75efb0efc2eff2ef3cf064f0d1f091f17cf2d8f379f592f6f7f7;
    decBuf[728] = 256'hdff809f97cf99ff9bff915faccfaa2fba4fc53fdb2fd22fdcefbd0f9e4f62cf4;
    decBuf[729] = 256'hfdf0ffed46eb82e9e6e7dbe5ffe34fe2c6e061df1cdef5dc36dc41dba6d91dd8;
    decBuf[730] = 256'h52d627d4b1d2e5d12cd164d163d204d46ed652d90adceedf8de3b9e88cedeef1;
    decBuf[731] = 256'h31f807fe55038809081118182e22432ea239ec466f53ce5e3066376a6f6b1b68;
    decBuf[732] = 256'h0b61cb58cf4eba429b3a45308e290421781b6814270c63044bf9f5ee8fe594da;
    decBuf[733] = 256'h3ed088c96ec31ac01cc1b2c587cb61d5c7dec2e924f18afa1403a008ab0d4112;
    decBuf[734] = 256'h6c16ba1b8d20ae23aa274a2ba42dec2ea53169330435a5376a39a93b1f3deb3d;
    decBuf[735] = 256'h293e803d813ce03a5739f237ae36db35b535a936c537b839943bc93ce23daf3d;
    decBuf[736] = 256'h0d3c3439b4358830552a7f24ad1d4217c10fb208710075f6bfef34e770df65da;
    decBuf[737] = 256'hcfd5a4d1e2d0d1ce71cf03d088d0e1d205d584d8c0dce0e113e893efa3f6e4fe;
    decBuf[738] = 256'he0084512d01a94229f27352cb52e772fc72ee62c0d2a6e263222591fb11a9017;
    decBuf[739] = 256'h70129d0d3c091c04aa0048fc6ff9e2f779f60bf66ff6c9f6c0f7a0f87cfab1fb;
    decBuf[740] = 256'haafd86ff3601300384043d0505056c04ca0261007dfd36f93af588ef3aea68e5;
    decBuf[741] = 256'h06e1e6db74d894d6ded45ad4c3d50cd7c4d9f3dcf1df71e3ace7ccec9ef141f7;
    decBuf[742] = 256'h8ffcc2029808e60d191444180e1c1f1e0020b5213021b8204b20e71fd81ee11d;
    decBuf[743] = 256'h6b1c8f1adf187516ed12a20fc90b2007be02c2fe23fbd8f7b4f5c3f368f3bbf3;
    decBuf[744] = 256'h30f584f6b9f742f9a7faecfb67fd66feaaffd10077020004cb05f7076d09490b;
    decBuf[745] = 256'h7e0c960d2f0e5e0e880eae0e8b0e2c0ed60d1f0dea0b6f0a0a09c6074b064c05;
    decBuf[746] = 256'h1d05f3041905c805a506a8075608f40884099e0987091a091b08e1061205e602;
    decBuf[747] = 256'hdb00fffe4ffd36fcd1fae9f9c2f81cf704f69ff4fdf2e5f1e6f0feef7fefc0ee;
    decBuf[748] = 256'h57ee77ee93ee4aef7ff0a6f14cf3d5f43af67ef7faf8f9f9e0fab3fb26fc49fc;
    decBuf[749] = 256'ha8fc8bfc71fc59fc18fcdefb84fbf2fa41fa6cf969f875f758f64bf5ccf367f2;
    decBuf[750] = 256'hc5f03def72edc1eb38ead3e8d5e6f9e4c5e3cbe177e0bedfa6de0dde81dd03dd;
    decBuf[751] = 256'h90dc27dcc8db39db1fdb07dbf1da05db17db06db33db40db64dbc7dbf0db14dc;
    decBuf[752] = 256'h35dc03dce8db00dc44dccddcf3ddc2df73e1dce377e583e7e7e982ebf8ecd4ee;
    decBuf[753] = 256'h08f021f1baf1e8f167f28df2b0f2d0f2b3f2fcf1f7f077efe0ec67ea27e8f1e4;
    decBuf[754] = 256'hcde215e050de10dc9bda47d912d8dad7a7d78fd80adad5db00de37e135e4b5e7;
    decBuf[755] = 256'hffea23eddbef55f2f0f3d0f414f5d7f42ef495f3adf2dbf1cef094ef6dee14ed;
    decBuf[756] = 256'hcfebfdeaf0e9fce81fe88fe70ce7c5e65ce70de842e9bdea88ec38ee31f00df2;
    decBuf[757] = 256'hbdf346f545f62df7acf7d2f769f7cbf6c8f58ff468f3c2f1a9f0aaefc2ee44ee;
    decBuf[758] = 256'hd1edaeed10ed46ec5bebffe9bbe894e787e61fe6c0e5a3e589e571e505e5a3e4;
    decBuf[759] = 256'h49e4f8e3aee3bce397e31ee36ce296e15ae033df26de78dd58ddaedd65de6bdf;
    decBuf[760] = 256'ha4e020e285e326e51fe773e81aeb49ee22f2d4f72a00260a3a16d9249c32b242;
    decBuf[761] = 256'hd451975ff364d3694d6b46672c6168595450c9470540f6388a32b52ce325a21d;
    decBuf[762] = 256'ha613910732fcf4eb25e162d372ca93c525c17cc226c6b2cbc6d450dd4ce7b2f0;
    decBuf[763] = 256'h3cf900010c06770ca210f015c21a241f2023c0261a29622a8d2b9c2c932d092f;
    decBuf[764] = 256'h6d31ad33e336e1399a3ca93da03ec03df43c3b3c923bc53bad3c7c3ea8404943;
    decBuf[765] = 256'h0d45a946f346af46ff440643923f473c9337f131a32c6f269a204c1b1815980d;
    decBuf[766] = 256'h880647fe83f674ef33e7a7e1a0deb5dde0dca2ddb3dfd4e2ade53be795e993ec;
    decBuf[767] = 256'h4cefe4f386f9d4fe0805dd0aaf1145161b1ce51f57233725ed266826ff24b623;
    decBuf[768] = 256'hfe20cf1dd11a511707140811890d2f0b0b091a070a065d06d207360a640e6012;
    decBuf[769] = 256'h11185f1dd120f323a8252c26c324a022ae20801da6190716bc12080ea6098604;
    decBuf[770] = 256'hb3ff11fac3f490eebae86ce39ade38da83d8f5d66dd791d910dd4ce16ce63eeb;
    decBuf[771] = 256'he0f02ef662fce203f60c81157d1f3326be2e4a345539403a153b533ae136c033;
    decBuf[772] = 256'hc42f1b2bba269a21c71c65184613730ed108830311006ffaa5f633f352f1c0f0;
    decBuf[773] = 256'h4ef289f6ccfc4d04610dec15b01dbf245529d52b972c482de82d332cae2b5429;
    decBuf[774] = 256'h5626d6229b1e7b19a91447106e0dcf097507510527041703c502100364041406;
    decBuf[775] = 256'h5e09990d95113e16a01a9c1e3b2295249427be28ce29202ad529f927d724fd20;
    decBuf[776] = 256'h551cb2166411920c70099806f8029e007bfec2fb49f9aef7a2f5d6f414f5bcf5;
    decBuf[777] = 256'h87f7b3f954fccdfe5602a1059f08580bd10d1110f11035117c10630f640ec30c;
    decBuf[778] = 256'h3a0b6f09bf07c60562037e00c5fd97fabdf627f4bdf29af036f091f0e3f0c3f1;
    decBuf[779] = 256'h8ff2c4f3ddf442f6e3f76cf937fbe7fc70fe3b00700118024b02c001ee0047ff;
    decBuf[780] = 256'hdefcfaf97af63ff243eea3ea68e68fe302e2a8df84dd93dbced933d853d70fd7;
    decBuf[781] = 256'h4cd746d9aadb32df7de231e753ea4feeeef12af626fabdfc07002b0255036504;
    decBuf[782] = 256'h1204c803740248003dfe51fbd1f787f4adf00eedc3e9c4e6d3e40ee3bce271e2;
    decBuf[783] = 256'hb5e2eae373e5d8e679e8e3ea23edc3ef3df27df41df7e2f8d9f923fadff9a2f9;
    decBuf[784] = 256'hf9f860f8d5f7abf738f789f62ef52ff3cbf0e7edf6eb7ce9e1e76be69fe5e6e4;
    decBuf[785] = 256'haee415e443e4c2e4cee54ee719e945eb50ed3cf0f4f26ef5aef7b9f995fbcafc;
    decBuf[786] = 256'h72fd3ffd57fcdcfa11f961f7d8f5d9f4f1f3caf2bdf184f0b4ee88ec7deaa1e8;
    decBuf[787] = 256'hf1e6d8e53fe56ee5ece5ace615e773e790e7aae7c2e703e865e806e99de927ea;
    decBuf[788] = 256'h5cea8dea43eab0e9d8e8d6e756e68be45fe2bedf90dc6cdab4d7efd554d409d4;
    decBuf[789] = 256'h4dd407d5afd514d759d828dad8dbd1dd35e075e216e544e843eb50f084f6afff;
    decBuf[790] = 256'haa0af4170a282c37de48c254915f66699c67fc658e6129582e4dd842213c9733;
    decBuf[791] = 256'h0b2e00293f266a201c1b27129c0968fd09f2bfe4d0dbb0d34eccf7ca2fccbbd1;
    decBuf[792] = 256'hcbd8e1e246ecd1f495fca0010b088c0a560e671088136116f718511b9a1cc41d;
    decBuf[793] = 256'h891f24212f231b26d428022cdc2f7b33d535d338fe39583aab3aca3976384237;
    decBuf[794] = 256'h99366636f1366d38d239733b8c3c253d3d3c6d3ac637e3333a2fd82adc263422;
    decBuf[795] = 256'hd21dd61936160a11370c9506c3ff58f9d7f1c8ea32e607e23dde2cdc8cdbfada;
    decBuf[796] = 256'h75daeeda36dc61dd25df0ae289e5c4e9c1ed60f19cf598f937fd820080037205;
    decBuf[797] = 256'h8106d4068906bd050405cc04330461043704c4031503b90118001ffe43fc0efb;
    decBuf[798] = 256'h66fafffafdfce9ff6803a4077d0a1c0e850fce106a105b0f1b0de509e606a002;
    decBuf[799] = 256'ha3fefbf999f579f008eda6e8aae40ae1cfdcf6d956d6fdd3d9d13dd24cd330d6;
    decBuf[800] = 256'hb0d9ebdde7e190e6f2eaeeee96f3f8f718fdeb018d07db0cad110f16e818751a;
    decBuf[801] = 256'hee1aa5197b1801161d139e0f440d450a5408da053f043402e000abff92fe2dfd;
    decBuf[802] = 256'he9fb16fb56fa33fad1fa0efc31fed2004c0330062108e609380a830a3f0a010a;
    decBuf[803] = 256'h5909c00891081308a00737075a061e05f703ea02b001de006a004800a6007001;
    decBuf[804] = 256'hc3026504ce060e09af0b280e6810de113213eb132314f013c213ef122f123b11;
    decBuf[805] = 256'ha00f170e800b06092206a30258ff35fd7cfa4ef72af572f2adf06deef8eca4eb;
    decBuf[806] = 256'heaeab2eae5ea70ebefeb62eccaec69edf8ed4cef91f060f210f499f5fef689f7;
    decBuf[807] = 256'h08f8e1f7bef720f757f6a0f5caf4c8f3d3f2f6f1f3f0ffefe3ee23eebaed1ced;
    decBuf[808] = 256'hffec19ed31ed47ed82ed70ed5fed6eed61ed6deda4edaeeda5ed7ced0bed79ec;
    decBuf[809] = 256'ha1eb9eeaaae98de834e793e50ae4d9e1cedff2ddc6dbbbd9dfd7aad691d55ed5;
    decBuf[810] = 256'h30d55ad51ad6c8d6e5d73ed926daa1db06dda8de30e0fbe1ace3a5e581e731e9;
    decBuf[811] = 256'h2aeb7eecb3ed5beef4ee7fef55ef7cef59effaeeddee8fee48ee07eecceddeed;
    decBuf[812] = 256'h0eee1dee45ee6aee49ee17eec5ed4cedb9ec7eec25ecf4eb03ec2bec50ec9dec;
    decBuf[813] = 256'hbbecd6ecefecf6ec19ed5ded9dedf8ed4dee84ee7aee5eee04eeafed78ed5aed;
    decBuf[814] = 256'h51ed7aed81ed5fed1aed91ecbaebf0ea39eac3e904eadbea18ec93ed5eef93f0;
    decBuf[815] = 256'h1bf21af302f4d5f448f5f6f5d4f62af744f72cf76af6b3f5ddf4a1f3cef2c2f1;
    decBuf[816] = 256'hcef0b1efa4ee6aed98ecd8eb6feb50eba6ebf4eb6becd7ec12ed24ed14ed22ed;
    decBuf[817] = 256'h15ed6aedf9edaaeeafefa3f041f15ef10ff13af08aee56ed3dec3eebb3ea89ea;
    decBuf[818] = 256'h16ea67e90be80de6a9e36ae1f4df18de5fdd97ddcaddb2de84df44e038e1d6e1;
    decBuf[819] = 256'hd9e213e437e66de921ee45f64100550cf41aa52c4b3d6e4c315a206300687a69;
    decBuf[820] = 256'h7365595f5d55f84b6d43a93b9e363330082c3e286b23881c48144c0a37fed8f2;
    decBuf[821] = 256'h76eb10e267de4bdd4edee3e264ea78f303fcff05640f7e150a1b111ed120a621;
    decBuf[822] = 256'he4209521f4206320de1f661fd31f701fca1f1c2092216e239a253b28b42af42c;
    decBuf[823] = 256'h6a2ebe2f77309031f53296348f367b39fb3c45404443c3461d49414ba44b4a4b;
    decBuf[824] = 256'h0a49d445fa41523df038d033fd2e5b290d243b1f98194a14170e41086f01dafc;
    decBuf[825] = 256'h04f73af3c8efa7ec15ec88ea00eb92eaf6ea05eca1edacef20f36bf644faedfe;
    decBuf[826] = 256'h0e02e7047d07f5073e09da083509e3080208be078107b907ec0777084a09090a;
    decBuf[827] = 256'h430b160c890c7d0ddc0df90db00eb50f3511661306168018641b1d1ee11fd820;
    decBuf[828] = 256'h8d20c11f951d5f1a8616e612ab0eae0a0606a401cbfe2cfbe1f7e3f42af266f0;
    decBuf[829] = 256'hcbee55ed89ec42ed5bee26f0cdf2fbf5d5f974fdb00189042808820a800d3910;
    decBuf[830] = 256'h671366161e19981b331da91eed1eaf1e261d5b1bb4183b16fb13851231117810;
    decBuf[831] = 256'hb010af11f4121a14c115d916d8176318e2185519491a231c0f1f56237628482d;
    decBuf[832] = 256'hea32b436c6386639b1371134e52eb228dc228e1d5b173013ea10780d970bbe08;
    decBuf[833] = 256'h3107c8057f045503fa024c032d048105ac074d0a310ed9127b18c91d3b219d25;
    decBuf[834] = 256'h5227e02867281f276624ed21091fc21ac6162613fa0d2809c604ca002afdc1fb;
    decBuf[835] = 256'h79fadcfaa1fce0fe8101fb033a06db08a00a3b0c1b0d6f0ead0ee50eb20e270e;
    decBuf[836] = 256'h540d480c820a56084b06d7028dffd8fa76f67af2d2edb0ead8e74ae6e1e473e4;
    decBuf[837] = 256'hd7e431e528e673e6c7e7fce885ea50ec7bee1cf196f3d5f5e1f7bdf96dfb15fc;
    decBuf[838] = 256'h48fc1afc9bfb8ffa55f92ef888f66ff50af469f250f1ebefa7ee80ed73ecc5eb;
    decBuf[839] = 256'he7eae5e936e959e8c9e77be7c2e72ee8dfe8b5e97eea35ebdbeb1cec2fec65ec;
    decBuf[840] = 256'h75eca2ece4ecf1ece6ecdcec9cec62ec5aec46ec72ecbbecedec1aed44ed1eed;
    decBuf[841] = 256'hfcece9ecb6eccbec10ed50edcbed48ee9aeee3ee41ef65ef86efcceffaef34f0;
    decBuf[842] = 256'h77f093f0abf0d1f0caf0c4f0d5f0c5f0caf0f9f018f156f1b1f1edf124f242f2;
    decBuf[843] = 256'h15f2a9f107f119f0fdeea3ed02ec79ea14e9cfe7a8e6e9e53ae59ce446e42ce4;
    decBuf[844] = 256'h14e455e490e4e9e45be5c2e53ae6cde608e761e7d3e7ffe75de8b1e8d2e8f0e8;
    decBuf[845] = 256'h1ee905e9e0e8bde860e802e8dee77be738e744e74fe7bde77de868e945ea81eb;
    decBuf[846] = 256'ha8ec68ed5ceebbeed8eef2eeabee13ee8aede9ec27ec3beb1feac5e881e7b1e5;
    decBuf[847] = 256'h86e37ae19edf73ddfddba9daf0d947d9aed8ddd807d9e0d803d962d97fd9cdd9;
    decBuf[848] = 256'h44dab0da88db8bdcc5dd40df0be1bbe295e514e940ee74f4f4fb080504104e1d;
    decBuf[849] = 256'hd0296f384342334b5253cc547553cb4f3f4a3043ef3a2b33202e8a29b423ea1f;
    decBuf[850] = 256'h781c1718d311fe0ba803e4fbd0f2b6ec2ae727e612e792e964f0d0f6fbff8508;
    decBuf[851] = 256'h49105917191a991cd71b271b06182d1597124c0f030ed90cc90b770b570c9b0c;
    decBuf[852] = 256'hd00d590f24115013f1156a184e1b071e802009245427522ad22d0d32e6348538;
    decBuf[853] = 256'hd03bf33d1e3fc33ecd3dc13b4d3812341630642a16254420e21bc216f0118e0d;
    decBuf[854] = 256'h6e089b03f9fd2ffa5df5fbf0ffec68ea0ee8c6e662e608e65ae63ae706e83be9;
    decBuf[855] = 256'h54ea53ebdeeb05edc4edb9ee96ef26f074f0bbf04ff0c6efddee00ee37edb4ec;
    decBuf[856] = 256'h6dec57ec92ecc8ec5aede3ed84ee47ef32f04ff1f5f27ef4aff64ff9c9fb52ff;
    decBuf[857] = 256'h9c0276060c09570c7a0ea50f4a0f540ede0cf209720628034effaffb64f841f6;
    decBuf[858] = 256'h88f30ff1cfeec4ece8eab3e99ae867e896e8bde9afeb13eef8f077f4b3f8affc;
    decBuf[859] = 256'h4e00a802a7059807a808fa08af08f3083a08020869073a07bc0649069b053c05;
    decBuf[860] = 256'hac045e041604010414046e040005ff053907b408190aba0b430d420e2a0ffd0f;
    decBuf[861] = 256'hbd106b110912991250139713ad137213ad128e113410930e0a0da50bbd0aeb09;
    decBuf[862] = 256'h780955097409cb09810a570b5a0c940dbb0e1410591180128c13c614ed154617;
    decBuf[863] = 256'h2e185519c819eb190e19d11702165b13e110fd0d7e0a240825056d02f3ff58fe;
    decBuf[864] = 256'h4dfc71fac0f838f739f6f4f421f4aef346f3e7f2caf218f360f3ccf355f4d2f4;
    decBuf[865] = 256'h23f550f578f56cf561f543f53af521f50af5daf4a2f45ef41ff4d4f3b6f39bf3;
    decBuf[866] = 256'h93f3a9f3bef3d1f3edf3fcf3f7f3d1f399f346f3e3f286f249f212f2f4f1ebf1;
    decBuf[867] = 256'h04f20bf212f2fff1e3f1bff196f185f175f17af176f162f13cf104f1c0f06ef0;
    decBuf[868] = 256'h21f0efefafef65ef1fefbaee27ee4fed86ec9bebbeeaf4e972e9fbe8bae87fe8;
    decBuf[869] = 256'h91e8a1e809e981e934ea0aeb0cec00eddeede1eed5efb2f0b5f1a9f205f4a6f5;
    decBuf[870] = 256'hbff624f868f93bfaaefa17fb76fb92fbe1fb28fc69fccbfcddfcedfcdefc81fc;
    decBuf[871] = 256'h2cfcc9fb36fbacfa2ffa7df9d6f83ff8b6f738f7e7f680f63df631f610f62ef6;
    decBuf[872] = 256'h6ef6d9f65ef722f8d9f880f96dfa0cfb9bfb1efc95fc7ffc6bfc12fc5ffb8afa;
    decBuf[873] = 256'hc0f9a1f894f7a0f684f52af4e6f2bff165f021ef4eeedbedb8edd8ed67ee1eef;
    decBuf[874] = 256'hc5efb2f090f120f2d6f21ef35ff372f319f3e8f29ef25bf237f258f28af2eef2;
    decBuf[875] = 256'h82f30bf464f475f42bf462f35ff2e0f07befd9ed31ed98ecc6ec45ed05eef9ee;
    decBuf[876] = 256'h97ef27f0d8ef32ef19ee73eceaea1fe96fe7e6e5e7e4ffe381e35ae337e357e3;
    decBuf[877] = 256'h3ae320e3d9e26de20be2b1e1a1e1cde146e239e3b9e4eae68be96eed17f2f9f8;
    decBuf[878] = 256'h65ff90088b13e11df6295535b73c1c46364c8a4f884ec84bf245203fdf365331;
    decBuf[879] = 256'h442aae252e23641f531d311a5917b0124e0e2f095c04faff21fd94fbfdfcfcff;
    decBuf[880] = 256'h09053c0bbd12cd1938206324a926f82518241b206a1a1c154910e70b0f098107;
    decBuf[881] = 256'h090751080a0b380e1212b115ed19e91d8821d324ad284c2ca62e7f321f366a39;
    decBuf[882] = 256'h683ce83f414265448f45ea454f44ae417f3ea63afd355b300d2b9b273a233d1f;
    decBuf[883] = 256'ha71c4d1a2918381628158d1317123b10100e040ca0090508fa05a604ed034403;
    decBuf[884] = 256'hab02da020403dd020003e1025102ce01f90083ff1efe20fc44fa18f80df631f4;
    decBuf[885] = 256'h77f35ff22cf25af22df339f4b9f584f7b9f842faa7fbebfc12fe1fff59008001;
    decBuf[886] = 256'hd9027a0473064f087b0a1c0d950f7a126b147b15cd15ed141113ee0fef0c7009;
    decBuf[887] = 256'h250627036e005fff68feb3fef7feb0ffe8ff810053007d00570034005300e300;
    decBuf[888] = 256'h0202a903a2050608450a510c2d0e610f9a0fcd0f410f1b0e5b0d210c4e0b420a;
    decBuf[889] = 256'h9309b608ed0736078f062306e805fa056c062c0717087309b70a330c980ddc0e;
    decBuf[890] = 256'haf0f6f10d710b810d41086109e10b310ee106b11dd1144126d124812cf11fc10;
    decBuf[891] = 256'hf90fbf0e980dd90c700c900c1f0d0a0e660f08119112f613dd1404167716e016;
    decBuf[892] = 256'h001756177017b717cd17b9178417121752163315d91338123f10630e370c9609;
    decBuf[893] = 256'h1d07dd04d202f600cafe54fd88fc54fbabfa78fa4afa20fa93fab6fad5faf2fa;
    decBuf[894] = 256'hd8fa91fa25fa9bf9d7f820f84af781f6caf524f58cf403f462f39ff2e9f142f1;
    decBuf[895] = 256'h54f0b6efedee6aee53ee68eea3ee20efd3ef79f067f145f20ef3c5f33bf4a8f4;
    decBuf[896] = 256'he2f4adf47cf432f4d5f398f38df383f38cf3a5f39df389f36af32cf3f2f2bdf2;
    decBuf[897] = 256'h64f20ff296f1e3f00ef044ef59ee7cedb3ecfceb26eb5dea72e9d4e80ae888e7;
    decBuf[898] = 256'h40e72be73ee774e7e6e712e855e8aae80de985e938eaafea46ebcfeb05ec36ec;
    decBuf[899] = 256'h62ec55ec49ec6aec4cec42ec5bec63ec77ecc9ec16ed84ed26ee92eef4ee71ef;
    decBuf[900] = 256'he3ef68f0e5f016f142f185f160f16bf19df1b9f103f285f202f394f31ef4bff4;
    decBuf[901] = 256'h2bf5b4f50df63ef64df625f6d0f56df5f5f4a3f495f487f4acf4e3f401f5f7f4;
    decBuf[902] = 256'hdff48cf413f460f35bf267f14af0f1ee09ee8bed18ed3bed99edf0ed3eee26ee;
    decBuf[903] = 256'h8feddeec09ec06eb57ea38ea1bea9eeaa3eb97ecf3ed94efadf012f2faf278f3;
    decBuf[904] = 256'hebf30ef4aff359f3d6f260f2c8f18df110f1bff075f0fdef8bef06ef66eeceed;
    decBuf[905] = 256'h1eeda7ec0fecd5eb7beb4aeb1eebf6eaeaeac9ea97ea69ea1feac5e970e9f7e8;
    decBuf[906] = 256'h85e81ee8a6e755e728e71be73fe78ce7d2e724e887e8e5e83ae9c9e952eaf3ea;
    decBuf[907] = 256'h0cec19ed99ee64f00bf339f613fabbfe5e04300b9b111b192b209626c12a8b2e;
    decBuf[908] = 256'h9c303c31872ff12ca629cd252421031e2a1b94182a17e215b714f312b310120e;
    decBuf[909] = 256'he40ae5072d05b302180163013f03e605ca09720ed412ad154c19c51957192d18;
    decBuf[910] = 256'hb31586118a0dea099f067c045103f70292049d06110a4d0e4912e9153319571b;
    decBuf[911] = 256'h0f1e1f1fba209a2166221f23382437257c264e275b28c428a428db275326e923;
    decBuf[912] = 256'haa21731e9a1a0318b91495126b11a60f540f090f4d0f100f480f150f8a0e630d;
    decBuf[913] = 256'h090cc50af50845072c06c704e003b902ac01b800dbffd8fe29fe8bfd35fde7fc;
    decBuf[914] = 256'h9ffcb5fc7afc21fcd0fb2dfb96fa0dfa8ff93ef96af9c8f94dfa12fb95fbdcfb;
    decBuf[915] = 256'hf2fbb7fb81fb30fb04fbf6fa02fb39fb93fb31fcf4fc13fe6cff0e0107035b04;
    decBuf[916] = 256'h0b06b3064c07c106ef059504f4026b01a0ff6bfe53fdbafce8fc12fdd2fd80fe;
    decBuf[917] = 256'h1fffaeffc8ffb1ff9bff87ff99ff0b00e80005025e03000518067d07c2089509;
    decBuf[918] = 256'hbb099809fa08f707bd064205dd039902c6015301ea00cb00e700cd00b5007500;
    decBuf[919] = 256'h610073008300af000d017a01e101240279029a02900287025e02290215022702;
    decBuf[920] = 256'h4f029c0215038603ee0330043d0432040004ad0360031a03ed02d402eb022803;
    decBuf[921] = 256'ha40345040805f305d00699071c08c2085a09e309840a1b0bcc0b430caf0cea0c;
    decBuf[922] = 256'hb40c630cde0bf60a180aa3083e079c05a303c70117001efecafc19fb01fa02f9;
    decBuf[923] = 256'h1af847f7d4f6b1f692f675f65bf614f6a7f51ef5a1f4eef348f3b1f24ef2f5f1;
    decBuf[924] = 256'ha4f178f14ff143f122f1dcf09cf031f0caef87ef63ef6eefa0ef16f0c9f06ff1;
    decBuf[925] = 256'h32f21df3faf3fdf4f1f5cff65ef715f88cf8cdf8e1f8f2f803f92ff957f994f9;
    decBuf[926] = 256'hf7f91ffa43fa38fab6f915f927f80bf7b1f56df446f339f28bf1aef01ef0cfef;
    decBuf[927] = 256'h29efbdee5bee02ee90ed46ed03eddfecbeecb4ecbdecd6ecfbec47edb5ed1cee;
    decBuf[928] = 256'hafee39ef6eef9fefaeefa0efacefe3ef29f0b2f063f139f23bf330f40df5d6f5;
    decBuf[929] = 256'h8df604f770f7f9f72ff8a1f808f99bf924fac5fa31fb94fbc9fbd9fbe8fbf6fb;
    decBuf[930] = 256'he9fbf4fb12fcf7fbbdfb7afbf1fa68fac7f9d9f83bf871f7eff678f637f64bf6;
    decBuf[931] = 256'h80f6f2f63cf7b4f747f8a9f802f953f9bbf9fdf96bfa97faa4fa98fa77fa45fa;
    decBuf[932] = 256'h05fabbf975f923f9c0f862f80df8c0f78ef773f75af735f705f7b3f650f60df6;
    decBuf[933] = 256'hd1f5c6f50cf670f603f7b4f72bf897f8aaf8bcf88cf842f8fff7c2f78bf759f7;
    decBuf[934] = 256'h2cf702f7b0f663f61df6b9f576f551f530f526f52ff5f6f4b2f43cf489f384f2;
    decBuf[935] = 256'h8ff134f0efee1cee10ededeccdec23ed0feeeceeefefe3f081f111f25ff277f2;
    decBuf[936] = 256'h61f226f214f245f2acf225f3f8f3fbf4eff5ccf6cff77df89af9a7fae1fbb0fd;
    decBuf[937] = 256'h60ffca01ae0466074a0be90e34123215b2180c1b541cb81c5d1c0b1c951ab918;
    decBuf[938] = 256'h09178015b51389111410c00e0f0df70b920aaa092c0905092809c6098f0ae30b;
    decBuf[939] = 256'h840dee0f2e12ce1448178819281ced1d881f68203421f7204e204f1f0b1ee41c;
    decBuf[940] = 256'h241c751b561bac1bfa1b711c091d431d551d251ddb1c981c741c691cc31c301d;
    decBuf[941] = 256'hd21d951e4b1f2120ea20a12148220a23592341235623f4225322bc21e4201b20;
    decBuf[942] = 256'h641f8e1e8c1d971cba1b441a7918c916601420127f0f060d6a0bf50929096f08;
    decBuf[943] = 256'ha808db08c209950aa20b960cb20dbf0eb30f91102011d7117d12be12f912e712;
    decBuf[944] = 256'h7612d311ba10140f8b0dc00b94098907ad05fd03e402e501fd00d300fa001d01;
    decBuf[945] = 256'hbb0184026f03cb0410063607dd08f509f40adc0b060c2d0c0a0c2c0b2a0a3509;
    decBuf[946] = 256'hda0738062005bb037602a301e3007b005b007800c6003d01d401ac0276039504;
    decBuf[947] = 256'hee0590071909e40a940c1d0e1c0f04108210a810cb10ac101c10990fc30ec10d;
    decBuf[948] = 256'hcd0cef0bec0af8095a09ca084808d1073a07ff06c90698068a067c0670067b06;
    decBuf[949] = 256'h8506a106eb0631077107cb07f00711080708d9078f074907d2064006b7053a05;
    decBuf[950] = 256'ha7041e04c5039403a303cb0307048004f2047705f4056606ea068b074e083909;
    decBuf[951] = 256'h560a620b9c0c6f0d2f0edd0efd0ea60e240e4e0dd80b730a750899066d04f802;
    decBuf[952] = 256'h1c01e7ffcefe35feaafd2cfd6cfcbefb1ffb1dfa29f98af8c1f773f72cf716f7;
    decBuf[953] = 256'h02f7cdf67bf6f7f57af5c7f421f489f300f383f211f26ff103f1a0f023f0f3ef;
    decBuf[954] = 256'hc6efd4ef10f073f006f1def1e1f21bf496f595f6daf701f9c0f929fac7fa57fb;
    decBuf[955] = 256'hdafb50fc91fca5fc6ffc1efc5efba7faa2f9aef891f738f650f529f4d0f2e8f1;
    decBuf[956] = 256'h15f109f0a0ef02ef72eef0ed79ed0ded83ec2aecd9ebcaebf2eb5fec01edefed;
    decBuf[957] = 256'h0cefccefc0f05ef1b4f103f2bbf14ff1edf04cf0e0efa5ef93efe5ef69f00af1;
    decBuf[958] = 256'hcdf184f22af396f3d1f3e3f3d3f3e1f30af446f4d5f45ff523f6daf6b0f779f8;
    decBuf[959] = 256'h30f9a7f9e8f9fbf97ef9ecf814f811f763f685f52ff5adf465f424f49bf31ef3;
    decBuf[960] = 256'h6bf2c5f102f180f0d9ef99ef36ef25ef35ef61efbfef5cf01ff10af227f333f4;
    decBuf[961] = 256'he2f4fef5bef66df70bf89af81df994f900fa14fa02fad1f987f92af9bcf838f8;
    decBuf[962] = 256'hdef74cf7c3f669f6d7f54ef5f4f483f41bf4f3f3b7f396f38cf35ef314f3cef2;
    decBuf[963] = 256'h45f2bbf11bf158f0a1effbee63eeb3ed3cedd0ec47ecedeb5bebd2ea78eae6e9;
    decBuf[964] = 256'h35e9bfe852e8f0e7bbe7aae77ee7a6e79ae7bbe7ede752e8cae89de966ea1deb;
    decBuf[965] = 256'hc4eb5bec96ecefecffec0eed36ed42ed63ed95edc3edeced12ee0beef8edd1ed;
    decBuf[966] = 256'h84ed21eda9ec37ecd0eb8deb81ebb8eb3aecfeece9ed45ef8af005f26af3aff4;
    decBuf[967] = 256'h81f58ef6f6f655f772f758f740f72bf717f770f7c2f70bf869f88df898f8a2f8;
    decBuf[968] = 256'h99f8b2f813f9a7f97efa81fbbbfce2fd3bff8000a70100034504c0058b07c008;
    decBuf[969] = 256'h490aae0b950cbc0d7c0ee50e830f13106110d81019117b11b011e111f011fd11;
    decBuf[970] = 256'hd911a2115c111c11c110b510c01006118f116712301350145c1550162e173018;
    decBuf[971] = 256'hdf187d19d319561a9d1a091b1d1b521b631b541b2c1bbf1aff191419f7179e16;
    decBuf[972] = 256'h5915321426137712d9114911fb10b4109e10d9103211a41164121b13c1135814;
    decBuf[973] = 256'hbb14f0142115f514971412144d132e12d410330faa0d790b6e0992075d064405;
    decBuf[974] = 256'h45041704ed03c703e903ca03ad03c703af03c50300045904ab04f4040205f604;
    decBuf[975] = 256'hbf0465041004ad033403e3027c021e02c9017c013601e4008100090077ffedfe;
    decBuf[976] = 256'h70fefefdd2fdfafd4ffec8fe5affe4ff3d008e00bb00c800bc009b007d002b00;
    decBuf[977] = 256'hdeff70ff08ffabfe56fe1ffe15fe0cfef3fdddfdacfd68fd16fdc9fc97fca0fc;
    decBuf[978] = 256'heafc58fdfafd92fe42ffe8ff55008f00a100910065003d00180023005500a700;
    decBuf[979] = 256'h0a018301b401e001d201ae0177016d018801e30181021803c9039f04f5047705;
    decBuf[980] = 256'h8f057a051705be046d040604dd03b903c403e203100439047c04aa04b204ab04;
    decBuf[981] = 256'h5104cc0307031c020001f3ff45ffa7fe17fec8fd52fde6fc35fc8ffbf7fa6efa;
    decBuf[982] = 256'h15fac3f9b5f9ddf919fa66fad4fa3cfb99fb06fc6efc96fcd2fcf3fcfdfcd0fc;
    decBuf[983] = 256'ha6fc45fccdfb5bfbb9fa4cfac3f98df97df98cf9cff924fab3fa15fbb6fb22fc;
    decBuf[984] = 256'habfc05fd76fda3fde5fd22fe2dfe37fe2efe15fef0fddbfdaffdaafda5fda9fd;
    decBuf[985] = 256'hb6fdc2fdbefdb5fd95fd55fd03fda0fc28fcb6fb4ffbf1fab5fa94fa8afaa5fa;
    decBuf[986] = 256'hcefa12fb52fb8bfb93fb8cfb6dfb2ffbe5fab3fa60fa29faf7f9b8f96df927f9;
    decBuf[987] = 256'hc3f865f841f820f83ef86cf8b6f8fcf83cf975f9c8f915fa6ffadcfa43fb86fb;
    decBuf[988] = 256'hc3fbcefbb0fb94fb6bfb46fb08fbcefa6dfa0ffaa2f93bf9ddf888f867f849f8;
    decBuf[989] = 256'h2ef815f80df8f9f7e6f7ecf7f1f7fff703f816f828f83ef869f8baf81df995f9;
    decBuf[990] = 256'h07fa8cfa2dfb99fbd4fb2dfc3dfc2ffc21fce5fb82fb3ffbd2fa6afaf2f980f9;
    decBuf[991] = 256'hdef847f86ff76cf6bef5e0f417f460f319f3d8f213f349f3baf33ff498f40af5;
    decBuf[992] = 256'h54f561f586f591f5aff5dcf537f68cf6d9f61ff74df755f72ff7e4f68af61df6;
    decBuf[993] = 256'hb5f558f51bf5e4f49ef44cf4fff3a5f338f3d1f28ef239f218f20ef217f261f2;
    decBuf[994] = 256'he3f284f347f432f50ff6d8f65bf7d2f713f875f8cef81ff9a4f945fadcfa66fb;
    decBuf[995] = 256'h2afcadfc53fdebfd74fecdfe1fff68ff91ff9dffbeff04006800fb00ac018202;
    decBuf[996] = 256'h840378045605e605d1063007f907b0085609190a040be10baa0cca0d8a0ec30f;
    decBuf[997] = 256'hea10aa11e412b713771425158415da15f415dc159c1561154f15fe140c153415;
    decBuf[998] = 256'ha21561164c172a182d19211afe1ac71b7e1c241de71dd21e701f73202121ff21;
    decBuf[999] = 256'h8f2245238d23f9233424fe23cd238423f0228e223522c321b4218c2168218921;
    decBuf[1000] = 256'ha721b021ea210022f9210022d8218b2112218020f71f9d1f6d1f401f691fa51f;
    decBuf[1001] = 256'hb01fe21fb51f491fc51e001e151d371c351b411aa219d918ee17111747162815;
    decBuf[1002] = 256'h6814ba13dc12c01271122a121412da118011ee103d10970fd40e1e0e480d7f0c;
    decBuf[1003] = 256'hc80b210b8a0ad9093309c7083e08e40793072c0799063706b90548051b05f304;
    decBuf[1004] = 256'hcf04f004fa04f1040a05110518052b051a05ec04b3044304b1034f03d1026002;
    decBuf[1005] = 256'h5102440250028702a502ae02a6028f0251021702b6013e01cc004700caff58ff;
    decBuf[1006] = 256'h0effe6fef2fe13ff6dfff3ff700002016401be01ce01dd01cf0193015c012a01;
    decBuf[1007] = 256'hfc00d300ad009900860080007b0077006a005e003f001800e0ff9dff4afffdfe;
    decBuf[1008] = 256'h8ffe28fee5fdc1fdccfd12fe76fe09ffbaff31009d00ff003501450154017c01;
    decBuf[1009] = 256'hb80105027302f8027503e70331047404980477045904f5037c03ca02f4012b01;
    decBuf[1010] = 256'h3f0062ff5ffeb1fdd4fc44fcc1fb4afb0afba7fa72fa41fa15fad2f97df904f9;
    decBuf[1011] = 256'h72f8c1f71bf758f6d6f52ff5eff4b4f4a2f4d3f41cf5aff512f68ff600f70ff7;
    decBuf[1012] = 256'h02f7c5f64cf6daf556f5d9f487f45bf44ef442f44df443f427f41ff4eaf3c8f3;
    decBuf[1013] = 256'hc2f3c7f300f461f4daf44bf5b3f5f6f5e9f5c8f546f5c9f417f470f3d9f250f2;
    decBuf[1014] = 256'hf6f1c5f1b7f1c4f1d0f1f1f1d3f181f11ef18bf002f0ccefbcef05f099f070f1;
    decBuf[1015] = 256'h3af259f3ccf37bf49af47df4fbf384f3c1f2d6f138f1a8f05af072f087f0eaf0;
    decBuf[1016] = 256'h43f194f185f178f10bf186f0e5ef4eefc5ee6bee1aee0bee19ee3dee74eef6ee;
    decBuf[1017] = 256'h73ef05f08ff030f19cf14cf294f200f362f3bbf3ecf318f4f0f3b3f37cf30ef3;
    decBuf[1018] = 256'hc5f2b7f2abf2ccf226f37bf3b2f3f8f3eff3d6f3a2f33bf3d3f290f254f233f2;
    decBuf[1019] = 256'h65f292f2fef2a0f30cf495f413f523f514f5ecf47ff4faf3a1f34ff323f34bf3;
    decBuf[1020] = 256'ha0f32ff4e0f486f5c7f502f685f5f2f41bf4def20cf2fff051f031f04ef068f0;
    decBuf[1021] = 256'hdff076f1fff159f2aaf2d6f2c9f2bdf2b2f294f29df284f27df284f24bf208f2;
    decBuf[1022] = 256'hb6f127f176f0d0ef0def56eee0ed48edbfec42ecf0eb89eb61eb0cebebeae1ea;
    decBuf[1023] = 256'hd8ea01eb27eb65ebbfeb45ece6eca8ed93ee71ef3af0f1f068f1a9f1bcf1aaf1;
    decBuf[1024] = 256'h9af1a9f1b6f10bf284f2f6f298f32ff492f4ebf41cf50df500f5f3f4fef444f5;
    decBuf[1025] = 256'hcdf5ccf606f82df987facbfb46fd45fe2dff00000c01bb0198029b038f042d05;
    decBuf[1026] = 256'h3006240701080409f809d60a9f0b560ccd0c0d0d210d0f0dff0cd30cc50cd10c;
    decBuf[1027] = 256'h080d3a0d8d0df00d4d0ed30e730f361021117d12c2133d15a2164318cc19cb1a;
    decBuf[1028] = 256'h561bd51bfb1bd81bb81b9c1b4d1b651b7b1b671b791b481bc31a231a6019a918;
    decBuf[1029] = 256'hd3177d172f174617de17b618b819f21a191cd91ccd1d2c1e821e681e211eb51d;
    decBuf[1030] = 256'h041d5e1cc71b161b701a041a7a192119af180d181f1742163f150514de121e12;
    decBuf[1031] = 256'h2a11cb103b10b90f420fd60e250eaf0dec0c350cbe0b520bf00aba0a8a0a5d0a;
    decBuf[1032] = 256'h350af909960938099a08d80755077f06f0056d05c7042f04cd035003be025c02;
    decBuf[1033] = 256'hbb014f01ed0070003f00130005002a0061009300c000c8008500fcff24ff21fe;
    decBuf[1034] = 256'he8fc15fc55fbecfacdfa23fba6fb4cfce3fc1efd0cfdbbfc19fc56fb9ffa29fa;
    decBuf[1035] = 256'he8f9fbf955fae7fa98fb3efcd5fc37fd25fdd4fc14fcf5fa9cf957f830f724f6;
    decBuf[1036] = 256'h75f516f5faf4dff427f568f5a2f5d8f54af6b1f60ff77cf7c6f7eef7c9f766f7;
    decBuf[1037] = 256'heef65cf6faf5e8f518f6bbf67df79df85df90bfaebf922f99af7a1f5b5f2fdef;
    decBuf[1038] = 256'hceecabeab9e85fe855e9f6eb25efd9f33bf837fcd7ff30029e027301fafe16fc;
    decBuf[1039] = 256'h96f84cf503f4d9f233f32af435f699f8d9fa4ffc1bfdddfc54fb23f982f609f4;
    decBuf[1040] = 256'h6df2f8f0b4f0e8f152f436f7b6fa00feff00f0024b0354024900d5fc8af9b1f5;
    decBuf[1041] = 256'h1af3c0f053f0b6f0c6f1aaf49bf6caf9edfb18fd27fed5fdf5fc29fc79faf0f8;
    decBuf[1042] = 256'h8bf746f6c8f5a1f5c4f523f6b3f66af7b1f7f2f706f8f4f7e3f7f2f750f806f9;
    decBuf[1043] = 256'hf1f90dfb67fcabfd7efe8bfff3ff1300bdff3aff64fe62fd28fc01fbf4f900f9;
    decBuf[1044] = 256'h62f80cf8f2f7daf7eff703f8f1f7e1f7d2f7c5f7d1f7f2f738f878f8d3f80ff9;
    decBuf[1045] = 256'h1af924f9e4f879f812f864f78ef6c5f50ef538f4a9f3f2f2aaf26af256f244f2;
    decBuf[1046] = 256'h54f263f270f295f2b6f2fcf260f3d9f38bf432f5f4f5abf651f714f897f80df9;
    decBuf[1047] = 256'h4ef989f9bff9aef982f975f950f945f963f991f9ecf959fac0fa39fbaafb12fc;
    decBuf[1048] = 256'h6ffcacfce3fc29fd44fd5dfd64fd5efd57fd52fd57fd6efdaefd00fe4dfebbfe;
    decBuf[1049] = 256'h05ff47ff54ff5fff2dff11ffe8fee0fef5fe21ff6affc4ff31007b00be00e200;
    decBuf[1050] = 256'hed00e300b5009d0095009c00c80011017f010402a5026703ea039004fc045e05;
    decBuf[1051] = 256'h9405a40595056d051805cb045d04d9035c03c902190272010601a4006f007f00;
    decBuf[1052] = 256'hab0009018e01e7015902a302cb02ef0210031a0336034f0356037803b103e503;
    decBuf[1053] = 256'h31049f042405c4055c060c078307ef072a086008500841084e087308aa081809;
    decBuf[1054] = 256'hba09510a020bd80b670c520df10dba0e3c0f1210a2102511cb116212ec126913;
    decBuf[1055] = 256'hda1342148514a914e014ea14e114fa1410151715361552155715651561154615;
    decBuf[1056] = 256'h5015601574159c15f015a61691176e18fe18e919871a171b651bad1b971b831b;
    decBuf[1057] = 256'h721b611b531b7b1b871bea1b621cd41c761d0e1e701ec91efa1ece1ea51e511e;
    decBuf[1058] = 256'hd81da71d7b1d6d1dda1d5f1e241f0f20ec207c21ff21462230221d229f21ed20;
    decBuf[1059] = 256'h7620b31ffc1e861eee1d3e1df61c8a1c281cf31bc21b781b351be01a511aef19;
    decBuf[1060] = 256'h4e198c1809189217fb1699163f16ee15c2157f155b15661548152c152415f014;
    decBuf[1061] = 256'h96144114b21302135b12c41113119d100510a30f6e0f3d0ff30ecb0e5e0ed90d;
    decBuf[1062] = 256'h5c0da90cd30b440b8d0ae709a60944093209420951099409d009db09d109a409;
    decBuf[1063] = 256'h2809630878075b064f051504ee02e101ed00100047ff90fe19fed8fd9dfd8bfd;
    decBuf[1064] = 256'h7bfd4ffd0cfdb7fc28fc9ffbdafa58fa82f9f2f8a4f82df8c1f786f72df7fcf6;
    decBuf[1065] = 256'hd0f6a7f69bf690f69af6c8f6f1f626f764f77cf784f78bf778f75cf757f740f7;
    decBuf[1066] = 256'h33f71ff7ebf689f611f67ff5f5f478f407f4bdf395f370f339f31bf3dbf281f2;
    decBuf[1067] = 256'h44f2e1f183f147f1e4f086f019f0b2ef39efe8ee81ee74ee80eeb7ee25efc7ef;
    decBuf[1068] = 256'h8af075f152f21bf306f4a5f434f5b7f5fef514f627f616f6a4f55af5fcf4a8f4;
    decBuf[1069] = 256'h71f467f482f4ccf426f57bf5c8f50ef617f630f637f631f643f66bf6a3f6f6f6;
    decBuf[1070] = 256'h6ff7e0f765f8e2f854f980f98ef951f9d8f846f86ef7def627f6b0f570f55cf5;
    decBuf[1071] = 256'h4af55af569f541f51df5e6f478f4f3f376f304f39df28ff283f2baf228f38ff3;
    decBuf[1072] = 256'h23f4acf405f577f5def521f676f6eff640f7c5f742f873f8bdf8e5f8c0f889f8;
    decBuf[1073] = 256'h2ff8aaf72df7bbf636f6b9f568f501f5a3f44ef4d5f384f33af312f306f33df3;
    decBuf[1074] = 256'h83f3d5f338f460f43cf4d9f310f30ef2d4f0adef53ee6ced99ecd9eb70eb51eb;
    decBuf[1075] = 256'h34eb82eb6beb80eb94eb5eebedea68eaa3e9ece876e835e821e89ee830e908ea;
    decBuf[1076] = 256'h0bebffebddec6cedefed36ee77ee8bee9deeadeebceec9ee06ef27ef59efbdef;
    decBuf[1077] = 256'he5ef09f040f04af066f07ff095f0aaf0e2f0daf0e1f0e8f0b5f093f080f064f0;
    decBuf[1078] = 256'h69f089f096f0a9f0bbf0a5f091f07ef05bf022f0fdefbfef85ef60ef14eff6ee;
    decBuf[1079] = 256'hedeec4eecbeed2eecceeddee01ef21ef61efd7ef49f0cef06ff106f2b7f25df3;
    decBuf[1080] = 256'hf4f3a5f41cf5b3f53df6baf62bf793f70bf85cf8a6f804f940f98df9d3f913fa;
    decBuf[1081] = 256'h5dfaa3fabffae8fafffa05fb18fb29fb4dfb92fbecfb59fcfcfc93fd1cfebdfe;
    decBuf[1082] = 256'h55ffdeff7f00eb007401ce0140028902e7023c037303a503d203fc033f047f04;
    decBuf[1083] = 256'hea046f051006d30689075f08ef08a6091d0ab40a3d0b970b290cb20c530deb0d;
    decBuf[1084] = 256'hc20e8c0f431048113c125913b2149a156c16e016021722179216db1535154714;
    decBuf[1085] = 256'ha9131913cb1284129912ad12bf1210131f132c1351135c137a13a71302146f14;
    decBuf[1086] = 256'hf414951501168a169c168c166016e7153515be1426149d134413f212a9126612;
    decBuf[1087] = 256'h2912c61183114711fa10b41074103a10421056108e10ff1091111b12bb122813;
    decBuf[1088] = 256'h3b134d13fc1295121c12aa112611a9105710f00fad0f580f0b0fb10e2c0e8b0d;
    decBuf[1089] = 256'hc80cdd0b000bfd094f09b1085a080c08c507af074d07d0063e06b4055b052a05;
    decBuf[1090] = 256'hfe040b0530053b051d05ef0484041d04a4031203b00256022602170224023002;
    decBuf[1091] = 256'h51026f0266023d02fa018301f1006700eaff78ff11ffb4fe8ffe6efe64fe6dfe;
    decBuf[1092] = 256'h97febcfedefe17ff2dff34ff2eff06ffcefe9afe40fed3fd6cfdf3fc61fcd8fb;
    decBuf[1093] = 256'h37fb74fabdf9e8f8e5f737f759f6c9f57bf563f579f58df5c2f5f3f51ff62df6;
    decBuf[1094] = 256'h39f65af68cf6ccf616f75cf777f76ff749f7fef6a4f64ff602f6d0f5b5f5bdf5;
    decBuf[1095] = 256'hd3f503f648f688f6c2f6e7f6fcf6f6f6daf6a1f66df63df604f6dff5caf5b7f5;
    decBuf[1096] = 256'ha7f5a1f59df599f5a4f59af58af57cf554f52df513f505f512f535f55ff586f5;
    decBuf[1097] = 256'haaf5a5f5a1f59df5a1f5c3f508f64ef68ef6c8f6b2f681f630f6cdf58af566f5;
    decBuf[1098] = 256'h87f5f5f597f65af745f822f9ecf9a2fa49fb8afbecfbfefbedfbdffbd1fbc5fb;
    decBuf[1099] = 256'he6fb18fc6afccdfc2bfd80fd8bfd81fd1cfda4fcf1fb1bfb8cfad5f92ff997f8;
    decBuf[1100] = 256'h35f8fff7eff7fef726f87bf8c8f822f977f9c4f9f6f911fa2afa31fa38fa32fa;
    decBuf[1101] = 256'h2cfa3cfa65faaffa1dfbbffbadfc8afd53fe0affb0fff1ffdeffa8ff57fff0fe;
    decBuf[1102] = 256'h92fe55fe1efe14fe0bfe24fe49fe7afeb2fed7fefafe19ff35ff44ff5cff68ff;
    decBuf[1103] = 256'h83ffaaffd8ff10006300b0001e016801aa01b701ac015201e400420080ffc9fe;
    decBuf[1104] = 256'h22fe60fd11fd9bfc5afc46fc58fc48fc57fc64fc40fc09fcd7fb84fb37fbf1fa;
    decBuf[1105] = 256'hc4faabfab3fab9fad9fa00fb2efb66fbaafbeafb34fc7afca8fcf2fc24fd64fd;
    decBuf[1106] = 256'haefd08fe5dfeaafef0fe0bff03ffedfebcfe9dfe81fe86fea7fed5fe0eff42ff;
    decBuf[1107] = 256'h72ff78ff68ff2fffddfe64fed1fd48fdcbfc39fcd7fba1fb70fb44fb1cfbdffa;
    decBuf[1108] = 256'h92fa4cfafaf9c3f991f976f97ef985f9b6f907fa54fad6fa53fbe5fb47fca1fc;
    decBuf[1109] = 256'hd1fce0fcd3fc96fc75fc6bfc62fc8bfcc0fcd4fcf4fc05fd14fd34fd74fdfdfd;
    decBuf[1110] = 256'haefeb3ffa70084014e0204037b03e70322045804a904f3045005be0507068006;
    decBuf[1111] = 256'hf10676071708da089109960a440be20b720cf50c3c0d520d650d770d870db40d;
    decBuf[1112] = 256'hc10dfe0d4b0e7d0ecf0e320f750fe20f4910c1103311b8111112831208136113;
    decBuf[1113] = 256'hf3137d141e150b16e916b217d118de198c1a2b1bba1bd41bbd1ba71b451bec1a;
    decBuf[1114] = 256'h7a1af519bf196e195f196d19a919ca19241a611a6c1a621a471afc19b6196419;
    decBuf[1115] = 256'h0119be1882184b18551870188918bd18e018da18bd187118e21731175b165815;
    decBuf[1116] = 256'haa14cd13031381123a12f9110c121e122e125b124d1229121e12d811aa119211;
    decBuf[1117] = 256'h9911a011cc11fe11211259127e129312a612951267122f12cd115511e3105e10;
    decBuf[1118] = 256'he10f6f0f080f750ec40def0cec0bf80a1a0a1809af081108bb076c07f5065e06;
    decBuf[1119] = 256'hd50510055904b3034703bd0264021302ac0169011401c70081002f00ccff6eff;
    decBuf[1120] = 256'h01ff9afe21feb0fd48fdebfc96fc49fc03fcd5fbbcfba6fb9ffb8cfb65fb37fb;
    decBuf[1121] = 256'hfffacafaa8faaefae1fa3afb8ffbdcfbfafbdefb73fbd1fa3afa62f9d2f84ff8;
    decBuf[1122] = 256'hd9f7c3f788f752f701f79af622f68ff5dff438f4a1f33ff3c2f271f244f237f2;
    decBuf[1123] = 256'h5bf292f2d8f22af3a3f3f5f33ef49cf4a8f4c9f4bff4b6f4aef4b5f4a1f49af4;
    decBuf[1124] = 256'h8af447f4f5f392f319f3a8f27bf253f247f27ef2b0f2def2f7f2eff2cdf294f2;
    decBuf[1125] = 256'h51f211f209f2f2f122f274f2d7f26af3f3f394f400f58af5bff5cff5a3f560f5;
    decBuf[1126] = 256'h0bf5bef464f428f407f4e9f3e0f3e8f3c2f3a0f374f32bf3e5f2b8f27ef267f2;
    decBuf[1127] = 256'h6ef274f27af294f28ff29cf2bff2dff21ff395f307f4a9f46cf523f6c9f635f7;
    decBuf[1128] = 256'h97f786f775f72cf7cef691f62ef6ebf5dff5bef5c8f5f6f50ff616f61df6e5f5;
    decBuf[1129] = 256'h92f52ff59cf4ecf345f3aef2fdf1b6f175f13af105f1d4f0a8f080f05bf03af0;
    decBuf[1130] = 256'h58f061f08bf0bff0c6f0b3f097f04af0fdefb7ef77ef3eef36ef14eff4eefaee;
    decBuf[1131] = 256'he0eed3eee8eee4eee0eef0eed0eea2ee76ee2deefbed16ee3feeb0ee83ef4cf0;
    decBuf[1132] = 256'h38f115f2def22df374f389f34ff3f5f2a4f278f26af246f23bf245f22af2f0f1;
    decBuf[1133] = 256'hbbf154f1edf0aaf055f0f2efafef2aefadee3beed4ed76ed52ed47ed79edefed;
    decBuf[1134] = 256'h61ee03efc6ef49f0bff02cf166f19cf1acf19ef190f16cf14bf141f15cf1a6f1;
    decBuf[1135] = 256'h14f2b7f24ef3fff3a5f43cf59ef5d4f5c4f5d3f5c5f5d1f5f2f54cf6b9f63ef7;
    decBuf[1136] = 256'hbbf74ef8d7f854f9a5f90dfa6afaa7fa0afb4dfba2fb05fc62fce8fc88fd20fe;
    decBuf[1137] = 256'hf8fe87ff3e008600c60001011301230132017501e2014902c20213033f034d03;
    decBuf[1138] = 256'h2803f102bf0292029a02ce023603ba035b041e05a0051706af06e9061f075007;
    decBuf[1139] = 256'h7c07bf07fc074908a308100977090a0abb0a610b240c0f0dad0d760ef90e6f0f;
    decBuf[1140] = 256'hb00feb0ffd0f2e105a108210bf100c115211b6112f1280120513821314149d14;
    decBuf[1141] = 256'h1a156c15b515de15b915981552150015c914ab147d1475148c14ae14f3145715;
    decBuf[1142] = 256'hb5152216a716dc164e177a176d1761174017fa16ba165f160a16a7154a15f514;
    decBuf[1143] = 256'ha814621422140914f313c313a313711333130a13e412c212e11214135113bd13;
    decBuf[1144] = 256'h24144c14701465141f14cd136a13f212c1129512a212c712e812de12c2127812;
    decBuf[1145] = 256'he2114b119a10f40f5c0fd30e320ec60d3d0d9c0c300c7f0b080b710a0f0a9209;
    decBuf[1146] = 256'h40091409ec08f8082f097509fe09870a280bc00b490c7f0cd00cc10c990c5c0c;
    decBuf[1147] = 256'h0f0cc90b9c0b620b3d0b360bfd0aba0a680ad9092809b108ef076c07f506b506;
    decBuf[1148] = 256'h7a0668067806870679066d064c06060690051e0599044004ef03e00308045d04;
    decBuf[1149] = 256'hc0041d0542054d0507057e04cd03c802d401f700f4ff45ff68fe9ffd1cfda5fc;
    decBuf[1150] = 256'h39fcd7fba2fb71fb62fb55fb49fb28fb0afbcafa90fa4cfa1ffa06fafff9f8f9;
    decBuf[1151] = 256'h0afa05fae1f9b7f963f90ef9c1f87bf84df856f85df880f8abf8bcf8b7f8a9f8;
    decBuf[1152] = 256'h7af84ff833f80ff801f805f8f9f7eff7ecf7c6f7a3f779f746f716f7eaf6adf6;
    decBuf[1153] = 256'h62f608f69bf516f599f428f4a3f36df33cf310f338f344f37bf3adf3c9f3e2f3;
    decBuf[1154] = 256'he9f3d4f3c2f3b1f3a1f3a6f3d5f30df460f4d9f44af594f5d7f5e3f5c2f590f5;
    decBuf[1155] = 256'h2cf5cef491f45af43cf446f46ff4a3f4fdf452f5cbf53cf686f6e4f639f75af7;
    decBuf[1156] = 256'h78f781f768f751f758f75ff786f7d3f720f87af8e7f813f93bf960f955f937f9;
    decBuf[1157] = 256'h2ef925f92df94ff955f945f92bf9e6f850f8b8f708f761f6f5f593f581f591f5;
    decBuf[1158] = 256'hbef5e6f53bf65cf68ef6a9f6b1f6b9f6cdf6e0f6f1f61ff74bf77ef7d7f714f8;
    decBuf[1159] = 256'h61f8a7f8d4f8edf8f4f8e0f8b4f898f86af857f873f897f8d3f82ef96bf9a2f9;
    decBuf[1160] = 256'hc0f992f958f906f98df81bf8d1f774f737f700f7cef68ef654f602f6b5f55bf5;
    decBuf[1161] = 256'heef486f444f4eff3cef3ecf3f5f31ef453f467f461f445f4f8f3abf379f339f3;
    decBuf[1162] = 256'h41f376f3c1f32ff4b4f40ef57ff58ef581f544f5f7f49df448f411f407f435f4;
    decBuf[1163] = 256'ha0f425f5c6f532f6bbf615f766f775f782f78ef76df777f792f79bf7c0f7f0f7;
    decBuf[1164] = 256'h29f86cf8acf8d5f80af92cf932f943f934f926f933f937f956f996f9faf958fa;
    decBuf[1165] = 256'hf5fa62fbebfb68fcb9fc03fd61fd85fdbcfd02fe30fe69febcfef3fe61ffe6ff;
    decBuf[1166] = 256'h6300f500cd019602b603c204b60594065d07e00756089708ab08e00832097b09;
    decBuf[1167] = 256'hf409a70a4d0b0f0cfb0c990d9b0e4a0fe80feb109911761240132b140815d115;
    decBuf[1168] = 256'h8816ff16961720187918eb1835195d199919a4199a199119891964196a197119;
    decBuf[1169] = 256'h7619c319261a841a091baa1b161ca01cf91c4a1d941df21d161e791ef11e431f;
    decBuf[1170] = 256'he51f5120b3203021612170217d2171213a2130211521eb20f320fa20e7200e21;
    decBuf[1171] = 256'h28213621652177217221772156211721c5206220ce1f6c1f131fa11e3a1edc1d;
    decBuf[1172] = 256'h571dfe1c6b1ce21b411baa1ad219091952184c179e168115c214cd132f136612;
    decBuf[1173] = 256'he3116d110111c6106c10fb0fb10f530fce0e510ebe0d350db80c460c1a0c0d0c;
    decBuf[1174] = 256'h190c3a0c800c9b0cb40cac0c7c0c1e0c8b0bdb0a050a3c095108b207e9066706;
    decBuf[1175] = 256'hc0055405f2045104e50334035f02cf01180172000600a4ff4aff19ffedfee0fe;
    decBuf[1176] = 256'hbbfe9afe7cfe4ffef4fd87fd20fd72fcccfb34fb84faddf946f995f81ff887f7;
    decBuf[1177] = 256'h25f7a8f636f6cff571f535f5fef4ccf4c3f4baf4d1f4f3f406f52df551f57bf5;
    decBuf[1178] = 256'hb9f5f2f545f6a8f6ebf640f777f781f753f72af7b9f627f69ef5fdf465f403f4;
    decBuf[1179] = 256'haaf359f32cf31ff3e2f2c1f253f2cff152f19ff0f9ef8cef03efcdeedeeeecee;
    decBuf[1180] = 256'hfaee36ef2bef21ef06efabee56ee09eeafed5bed24ed06edeaece2ecdaece1ec;
    decBuf[1181] = 256'hf4eceeece9eceeecd9eccdeccaecbaecb1ecc9ecd9ecfeec4bed82eddced31ee;
    decBuf[1182] = 256'h7eeeb0ee02ef23ef55efa7efdeef38f0a5f0eff032f156f14bf105f1c5f05af0;
    decBuf[1183] = 256'h10f0e8efc4efcfef01f01cf035f04bf01bf0e3ef9fef29efd8eeabee83ee8fee;
    decBuf[1184] = 256'hdcee22ef87ef1af07cf0d5f027f153f17bf19ff1c0f1def10cf235f25bf2a6f2;
    decBuf[1185] = 256'hd8f218f362f394f3e7f334f466f4a5f4dff405f519f539f533f52ef53cf526f5;
    decBuf[1186] = 256'h1bf525f51cf530f557f58af5d6f544f68df6ebf658f767f78ff783f74cf706f7;
    decBuf[1187] = 256'hc6f67cf64af62ef626f63df66df699f6b5f6cef6aef677f633f6bdf54bf501f5;
    decBuf[1188] = 256'ha3f47ff474f47ef487f4b0f4a9f4a2f476f422f4b5f34ef3d5f263f237f20ff2;
    decBuf[1189] = 256'h1bf252f25cf278f290f27af265f246f21ff205f21cf231f264f2aff2e1f20ff3;
    decBuf[1190] = 256'h38f331f30ef3eff2a6f274f246f20df2f6f1e1f1c2f1b1f1a2f178f146f116f1;
    decBuf[1191] = 256'hd1f091f057f014f0e6efbdef97ef90ef97ef91ef96efa4efa0ef9cef91ef82ef;
    decBuf[1192] = 256'h7fef97efbfef14f099f016f1c9f16ff2dbf23df373f383f392f385f391f3def3;
    decBuf[1193] = 256'h38f4bdf45ef521f6a3f649f7e1f743f89cf8eef81af95df9b2f915fa8dfafffa;
    decBuf[1194] = 256'h83fb24fc90fc1afdbbfd52fe03ffa9ff970074013d02f402ca0393044a05f005;
    decBuf[1195] = 256'hb3066a0740080909c009660afd0a870b280cbf0c480dc60d580eba0e370f880f;
    decBuf[1196] = 256'hd20ffa0f371058109e100211951146121c13e513d014ad1577162e17d4176b18;
    decBuf[1197] = 256'hf518b919701a461b491cf71c141ed31e821f2020e9203821ae211a227d22d622;
    decBuf[1198] = 256'h27235323b123ee23f9233f247f24b8240b256e25962503266a269226cf260627;
    decBuf[1199] = 256'h10272b2734270e270727dc2687264b26fe257c25fe248d24ea235323ca222922;
    decBuf[1200] = 256'h912108214320c11f1b1f581ea11d2a1d681ce51b3f1ba71a1e1a7d19bb186c18;
    decBuf[1201] = 256'hf5175e174a171517e416f316cb1676163f16bd151c158514fb133713b4123d12;
    decBuf[1202] = 256'hd1116f111611a4103d10a90ff90e530e900da50c070c3d0b870ae00949099808;
    decBuf[1203] = 256'h2208b5072c07af063d06b8053b05a90420047f03e70237029101ce004b00a5ff;
    decBuf[1204] = 256'h0effacfe76fe25fef8fd06fee1fdd6fdccfd9ffd76fd5ffd2ffd03fdfefce4fc;
    decBuf[1205] = 256'hdffcecfcf0fc01fd24fd3bfd50fd64fd59fd3dfd12fdbefc69fc06fc8efb1cfb;
    decBuf[1206] = 256'hd2fa75fa38fa17fa0dfa16fa2ffa45fa68fa87fa8dfaa6faabfa9efa9afa97fa;
    decBuf[1207] = 256'h8dfa90fa93fa9afaa9fab7fabcfac7fac6fab7faa1fa7bfa43fa00fac0f975f9;
    decBuf[1208] = 256'h43f904f9ebf8e3f8eaf809f93cf97af9b4f9f7f925fa3efa54fa4dfa3afa2afa;
    decBuf[1209] = 256'h10fa02fa06fa1afa32fa61fa91fab0fae3faf8fafefa04fbf4fad4faaefa7ffa;
    decBuf[1210] = 256'h47fa22fafff9f9f90afa19fa30fa46fa3afa14fad1f95af9e9f864f8e7f795f7;
    decBuf[1211] = 256'h69f741f74df758f762f76bf763f73ef71bf7fcf6d5f6bbf6c0f6bbf6c7f6dff6;
    decBuf[1212] = 256'hfcf626f759f77bf79af7cdf7eff71bf84ef870f883f89ff890f882f875f862f8;
    decBuf[1213] = 256'h50f853f85cf86ef892f8acf8c3f8d8f8dcf8d1f8cef8aff888f864f832f801f8;
    decBuf[1214] = 256'he2f7c6f7b7f7c5f7d1f7ddf7fcf7f8f7edf7dbf7acf77cf750f71ef7fbf6f5f6;
    decBuf[1215] = 256'hfbf6f6f616f71af716f71af710f7fcf609f71af736f770f7cbf707f854f886f8;
    decBuf[1216] = 256'hb4f8cdf8d4f8cdf8ecf809f937f994f9f2f95ffae4fa3dfb8ffbf6fb03fc0ffc;
    decBuf[1217] = 256'h1afce8fbbbfba2fb6dfb4bfb51fb40fb27fb35fb1ffbf5fad9fa96fa44faf7f9;
    decBuf[1218] = 256'h9df930f904f9a6f869f85ef82cf811f8f8f7b5f787f75ef71af7fff6f7f6eff6;
    decBuf[1219] = 256'hf6f615f71bf716f708f7c8f688f63ef6d0f5a4f57cf557f578f5d2f50ff672f6;
    decBuf[1220] = 256'hd0f6f4f615f71ff7dff6b6f672f60ef6e6f5c1f5b6f5c0f500f62af67cf6c9f6;
    decBuf[1221] = 256'h0ff761f782f7a0f797f77ef74af735f716f710f753f7b7f74af822f9ecf9d7fa;
    decBuf[1222] = 256'hb4fb44fcc6fc0efd4ffd89fd9bfdedfd54feccfe7fff55001e01d501da028803;
    decBuf[1223] = 256'h2704f0047205e9058106e3063c07ce075808b10864090a0acd0ab80b950c5e0d;
    decBuf[1224] = 256'h4a0e270fb70f6e10e4102511af1108125912c0123913ab134d140f1592156816;
    decBuf[1225] = 256'h3117b4175a18f1185319ad19fe192a1a6d1a921ac91a231b771bda1b6e1cf71c;
    decBuf[1226] = 256'h501de31d1d1e531e631e721e4a1e561e4b1e411e811e9a1ece1e1a1f381f531f;
    decBuf[1227] = 256'h6c1f551f331f141fcb1e851e571e0d1edb1dad1d631d1d1ddd1c721ced1b941b;
    decBuf[1228] = 256'h011b781a1f1a8c192a19ad183b18b7173a176616d71520151a146c138f12c511;
    decBuf[1229] = 256'hda103c10ac0ff60e7f0ebc0d3a0d930ca50b070b3e0a53097608e6072f078906;
    decBuf[1230] = 256'h1d066c05c6042e047e03d70240028f01e90052007affeafe68fec1fd2afdc8fc;
    decBuf[1231] = 256'h27fcbbfb59fbb8fa4cfac2f921f98af801f860f7c8f666f6e9f598f54ef5d6f4;
    decBuf[1232] = 256'h85f43bf4c2f351f307f3a9f285f264f246f261f26af262f25bf23cf2fef1c4f1;
    decBuf[1233] = 256'h81f12ff10ef1f0f0d4f0ccf0d4f0cdf0d3f0c2f0b3f0aef099f07ef06cf050f0;
    decBuf[1234] = 256'h3df032f01cf019f02cf038f04ff07ef0a0f0ccf0f3f0f9f0f4f0f8f0edf0e9f0;
    decBuf[1235] = 256'h05f120f155f1a7f1def124f276f2adf2b7f2d3f2dbf2e3f2f7f20af331f35ff3;
    decBuf[1236] = 256'h7ff3b1f3d4f3cdf3b1f398f352f30cf3dff2a5f27ff286f28df29df2b7f2bcf2;
    decBuf[1237] = 256'ha6f2a3f26ef23af217f2dff1b9f1b3f193f182f192f17bf165f15af133f105f1;
    decBuf[1238] = 256'hf2f0b5f07bf055f017f0cdef87ef35efe8eea2ee62ee28ee03eed3edb4eda3ed;
    decBuf[1239] = 256'h75ed3ced17edcbec85ec58ec1eecf8ebffebf9ebffeb2dec3fec50ec74ec70ec;
    decBuf[1240] = 256'h74ec78ec6dec64ec67ec5aec57ec6aec6dec8cecccecf9ec43ed9deddaed11ee;
    decBuf[1241] = 256'h43ee4cee54ee5cee47ee4eee6aee83eebfee1aef6fefd2ef30f06cf0b9f0ebf0;
    decBuf[1242] = 256'hf4f01ef143f166f19ef1f0f13df297f2ecf239f37ff3d1f31ef464f4c9f40cf5;
    decBuf[1243] = 256'h60f5adf5b7f5d3f5cbf5a5f590f597f59cf5caf51cf669f6aff613f73bf760f7;
    decBuf[1244] = 256'h81f777f780f777f77ff794f7bff7f2f730f87af8acf8ecf826f94bf96ef999f9;
    decBuf[1245] = 256'hb5f9e4f90ffa37fa65fa91fac3faf3fa38fb66fb8ffbc3fbe6fb12fc2efc29fc;
    decBuf[1246] = 256'h24fc20fc05fcecfbd0fbadfb8dfb80fb74fb71fb80fb95fbacfbc8fbd4fbd7fb;
    decBuf[1247] = 256'hd4fbc0fbaefb98fb84fb82fb8efba5fbcefbf5fb0ffc1cfc18fcf5fbccfb8efb;
    decBuf[1248] = 256'h44fb12fbd2fab9faa2fa8efa88fa82fa73fa6efa7bfa86fa98fac7faf7fa2ffb;
    decBuf[1249] = 256'h82fbcffb29fc96fcfdfc75fd08fe6afe0bff77ff00005900cb0032019001fd01;
    decBuf[1250] = 256'h8202ff02b2032904c0047105e70528068a06e40635079c07fa077f084409c609;
    decBuf[1251] = 256'h9c0a2c0be30b5a0cc60c280da50d170e7e0e110fc20f3810fb10b2112912eb12;
    decBuf[1252] = 256'ha213481436151416dd16c817a5183519ec19631afa1a841b241ce71c9e1da31e;
    decBuf[1253] = 256'h521f2f20f8207b2121228d22c8224523d7233a24da247225d4257526b626f126;
    decBuf[1254] = 256'h4a279b27c7274028b228fb288e29f129262a572a662a232a2f2a0e2af0291e2a;
    decBuf[1255] = 256'h572a7d2ac82afa2adf2ae72aa42a2d2adc297529fc28ab2861280428df279227;
    decBuf[1256] = 256'h1027b7264526a3253725ad240d247523ec2227227021ca200720511faa1ee81d;
    decBuf[1257] = 256'h651dbf1c271c9e1bd91a231a7c198e18b117e81631162c157d14a013d7122012;
    decBuf[1258] = 256'h1b1126100a0ffd0d090dec0be00a310a540951085d0780067d0589046c036002;
    decBuf[1259] = 256'h6c018e00c5ff0eff38fe6ffdb8fce2fb19fb62faecf929f9a6f830f8c3f73af7;
    decBuf[1260] = 256'he1f62ef6b7f520f56ff4c9f35df3fbf2c5f2b5f289f27bf26ff24ef208f2b6f1;
    decBuf[1261] = 256'h53f110f1a3f077f069f05df07ef0c4f004f13ef181f19df194f18df16bf14bf1;
    decBuf[1262] = 256'h2ff10bf1fdf002f1fef00ff132f149f167f191f1adf1c7f1f1f101f225f23cf2;
    decBuf[1263] = 256'h49f25df275f278f292f2c0f2dff228f382f3d7f324f492f4dcf41ef55bf57cf5;
    decBuf[1264] = 256'haef500f637f691f6fef648f7c0f732f87cf8f4f866f9b0f9f3f948fa69fa87fa;
    decBuf[1265] = 256'ha2fa89fa73fa5efa32fa21fa27fa2bfa49fa7bfa90faaffaaafa86fa53fa07fa;
    decBuf[1266] = 256'hadf958f90bf9d9f8acf8a3f89cf895f88ff867f839f801f8bef76bf734f7daf6;
    decBuf[1267] = 256'h9ef667f621f6cff598f552f524f5fbf4e4f4ddf4f0f401f510f515f5f7f4c5f4;
    decBuf[1268] = 256'h87f42cf4d7f3a0f36ef365f39ff3d4f311f44bf462f45bf42ff4dbf36ef324f3;
    decBuf[1269] = 256'habf25af22ef206f2e1f1d6f1b8f19df184f15ff13cf136f11af100f1f3f0c4f0;
    decBuf[1270] = 256'h8cf057f0feefc1efa0ef96ef9fefd9effeef3cf076f07ef077f064f031f01df0;
    decBuf[1271] = 256'h16f01cf040f07cf0b6f0eaf01af12df13ef158f15cf17af1b4f1ddf112f250f2;
    decBuf[1272] = 256'h69f27ff294f281f287f2aaf2c2f201f366f3c3f318f47bf4bef4e2f4edf4f7f4;
    decBuf[1273] = 256'h01f519f530f552f58af5b0f5d2f5f2f5f7f5f2f500f604f618f63ef658f66ff6;
    decBuf[1274] = 256'h8df689f68cf696f698f6b5f6eff64af7b7f73cf895f8e7f830f93ef94af929f9;
    decBuf[1275] = 256'hf7f8dcf8d3f8dbf8fdf835f96af9a8f9e2f907fa1cfa2efa29fa24fa28fa24fa;
    decBuf[1276] = 256'h28fa40fa5dfa8ffabffaf7fa3bfb7bfbb4fbf8fb26fc3efc46fc3ffc2cfc10fc;
    decBuf[1277] = 256'he2fbb6fb78fb4ffb2afb15fb1bfb37fb65fb9efbe1fb21fc4afc70fc84fc8bfc;
    decBuf[1278] = 256'h9cfcbffce9fc3dfddbfd9efe55ff5a000801e601af02fd027403e0031b049804;
    decBuf[1279] = 256'h0a058f0553060a07e007a9089409720a3b0bf20b980c2f0db90d5a0ef10e7a0f;
    decBuf[1280] = 256'h1b10b3108a111a120513a3136d14ef1496152d168f1630177117fa177718e918;
    decBuf[1281] = 256'h6e19eb195d1ac41a221b5e1bab1b191c631cdb1c6e1dd01d4d1e9e1eca1ef21e;
    decBuf[1282] = 256'hff1ef41efe1e2b1f541fc51f5720e120812119227b22d422e522f3220123f522;
    decBuf[1283] = 256'h00231e234b23642398239f2374234c23ff22862215229021ef208320d21f2c1f;
    decBuf[1284] = 256'h951ee41d3e1da61cf61b4f1bb81a071a321968187d176116541560148313b912;
    decBuf[1285] = 256'h02125c11f0103f10990fd70eeb0d0e0d450c250b190a6a098d08fd074607d006;
    decBuf[1286] = 256'h3806af050e054b049503bf02f6010a012d002aff36fe59fd90fcd9fb32fb70fa;
    decBuf[1287] = 256'hedf947f984f8cdf7f8f62ef678f572f4c4f3e7f21df29bf124f1b8f056f0fcef;
    decBuf[1288] = 256'habef44efe6ee91ee44eeeaed95ed48ed02ed9eec5beceeeba4eb61eb0debd6ea;
    decBuf[1289] = 256'hb8ea9ceaa4eabbeac2eae1eafdea0deb11eb0debeaeacaeaacea89ea84eaabea;
    decBuf[1290] = 256'hd9ea2aeba3eb15ec7cecdaec16ed63ed81ed9dedb5edf9ed39eeb5ee55efedef;
    decBuf[1291] = 256'h9df044f1dbf18cf232f39ef300f47df4cff418f576f59af5d1f517f633f65cf6;
    decBuf[1292] = 256'haef6e5f653f7d8f732f8a3f80bf94df95af97bf95df966f96ef984f9b5f906fa;
    decBuf[1293] = 256'h53fa99fad9fa02fb18fb1ffb0dfb07fb0cfbfefa0bfb1efb1bfb24fb2dfb20fb;
    decBuf[1294] = 256'h14fb12fbfcfae8fadafab7fa7efa59fa1bfae1f9bcf97ef955f93ef90ef9d6f8;
    decBuf[1295] = 256'ha1f848f8dbf774f7e0f67ef601f6b0f584f55cf537f516f5f8f4b8f45ef4f0f3;
    decBuf[1296] = 256'h89f311f3c0f258f215f2d9f1a2f15cf11cf1d2f078f03bf004f0e6efefefe7ef;
    decBuf[1297] = 256'hdfefe6efc7efa0ef7cef49ef19ef1fef30ef68efcaef42f0b4f01bf15ef19bf1;
    decBuf[1298] = 256'ha6f1b0f1a7f19ef197f1abf1cbf1f2f135f287f2d4f21af35af383f3a8f3cbf3;
    decBuf[1299] = 256'hc5f3caf3daf3e7f316f467f4b4f40ef57cf5c5f508f62df64ef658f661f669f6;
    decBuf[1300] = 256'h9df6e9f657f7dcf77df8e9f872f9ccf91dfa49fa71fa7dfab4fafafa4cfbaffb;
    decBuf[1301] = 256'h0dfc62fcc5fc08fd2cfd4dfd6bfd87fd9ffdb6fdcafdeafd06fe15fe23fe30fe;
    decBuf[1302] = 256'h43fe6afe98fec4fe0dff3fff7fff97ffaeffb5ffaeffa9ff99ff95ff99ffa5ff;
    decBuf[1303] = 256'hb6ffc6ffd4ffe7fff7ff060020003900550068007a0076006e00560040002c00;
    decBuf[1304] = 256'h1f00260039005600790090009d008a006a003300feffc0ff97ff90ff97ffb6ff;
    decBuf[1305] = 256'hddff01002100480061007800a700df0023017501d80136028b02d8021e037003;
    decBuf[1306] = 256'hbd0317049c043d05a9055a06d0063d079f07d407050831087408c9084209d409;
    decBuf[1307] = 256'h850a2b0bc30b250ca20cf30c3d0d9a0d200e790eeb0e700fc90f1a109f10d510;
    decBuf[1308] = 256'h6711f0116d122013f61386143d15e3154f168a16e316f3165b17b8173e180219;
    decBuf[1309] = 256'hed198c1a8e1b821ce11cab1df91d401eac1ee71e1d1f8f1f13206d201f219621;
    decBuf[1310] = 256'h0222b3222a239623f82375248524b224a42480245f2441240124092411241824;
    decBuf[1311] = 256'h5c248a24822489244b24e0237923e6223522be212721c5206b203b20d31fab1f;
    decBuf[1312] = 256'h561ff31eb11e431ea11d351dac1ce71b641b8f1aff194819a2183618d4175617;
    decBuf[1313] = 256'he5167d16ea15121549145e1341123511fb0fd40e140e660dc80cfe0b480b720a;
    decBuf[1314] = 256'ha90989083007eb05c404b8037e02ab01eb003d0060ffd0fe19fe43fd7afc8ffb;
    decBuf[1315] = 256'hb1fa22fa6bf995f805f84ef7a8f611f687f5e7f47af418f49bf329f3c2f24af2;
    decBuf[1316] = 256'hb8f12ef1b1f01ff095ef18efc7ee60ee02eec6ed79ed33ed05edcbec97ec67ec;
    decBuf[1317] = 256'h22ecd0eb83eb15ebadea50ea13eadce9e6e9efe908ea4cea79eab3ead8eadfea;
    decBuf[1318] = 256'hd9eadfeacfead4ea03eb2eeb83eb08ec85ecf7ec99ed05ee68eec1ee12ef3eef;
    decBuf[1319] = 256'h81efa6eff3ef39f079f0c3f031f198f110f282f2e9f262f3d4f300f443f47ff4;
    decBuf[1320] = 256'h8af4bcf4eaf403f546f586f5d0f516f668f69ff6e5f625f74ff774f7a4f7c3f7;
    decBuf[1321] = 256'hf6f726f852f890f8daf80cf95ef9c1f904fa59fabcfafffa3bfb72fb90fb9afb;
    decBuf[1322] = 256'hb2fbabfbb2fbc4fbbffbc4fbd2fbcefbd1fbd5fbccfbc3fbc0fbabfb97fb8afb;
    decBuf[1323] = 256'h66fb2efbf9faaefa54fa17facaf998f97df974f97cf990f997f986f962f91df9;
    decBuf[1324] = 256'h9bf81df8acf744f71cf710f71bf761f78ff7c9f7dff7d8f7b9f786f748f70ff7;
    decBuf[1325] = 256'he9f6c7f6c1f6ddf6ecf6faf618f71cf71ff722f71af712f70bf7f3f6ddf6c3f6;
    decBuf[1326] = 256'h9df66ff650f628f619f60bf607f60bf615f612f60ff607f6fbf5f1f5eff5e9f5;
    decBuf[1327] = 256'hf5f508f615f62bf64af657f67af69af6c1f6f9f62ef76bf795f7baf7cff7d5f7;
    decBuf[1328] = 256'hdbf7d6f7e3f701f834f87ff8c5f805f93ff946f932f9f9f8c5f887f85ef874f8;
    decBuf[1329] = 256'h97f8f4f852f9a7f9f4f926fa1dfa04fad0f99ff98df9a9f9ebf950fac8fa5afb;
    decBuf[1330] = 256'hbdfb16fc47fc73fc66fc59fc4efc58fc86fcc0fc12fd75fdeefd5ffea9feecfe;
    decBuf[1331] = 256'h29ff60ff7eff99ffb2ffd7ff15004f00a100ee00340162018b01a201a901af01;
    decBuf[1332] = 256'h9e01a301a801bd01e8010f023302530269026c02700273028d02c10214037703;
    decBuf[1333] = 256'hef036104e6043f0570059c05aa05ce0505067306da0688072e08c60828098109;
    decBuf[1334] = 256'hb209c109b309bf09e009120a770aef0a610bc80b0b0c2f0c240c1a0cff0be60b;
    decBuf[1335] = 256'hee0b1e0c560cb80c150d520d890da70d9e0da60d9f0d980db70df50d3f0ead0e;
    decBuf[1336] = 256'h320f8b0f1d108010d9102a117411b7110c128512f61299133014e11487151e16;
    decBuf[1337] = 256'h8016fe162e1720172d17391744177617c81715188318cd18f5180119ca185c18;
    decBuf[1338] = 256'hf5177d170b17fc1609172e177b17ad17b6179d174b17a616ff1568150615d014;
    decBuf[1339] = 256'hc014cf141215361541150f15ab1418146713c1125512f211e111d011fd11ef11;
    decBuf[1340] = 256'he311ac112a118910c70fdb0e3d0eae0d2b0de40ca30c410c0b0c990bf70a340a;
    decBuf[1341] = 256'h7e0978088407e6061d066605ef048304fa03a0030e035d02b701c900ecff5cff;
    decBuf[1342] = 256'ha5fe2ffec2fd88fd52fd01fd7cfcfffb6dfbbcfa16fa7ef9f5f8bff86ef842f8;
    decBuf[1343] = 256'h34f8f8f7abf729f788f6c5f50ef568f4d1f36ff339f329f31af30df3b8f255f2;
    decBuf[1344] = 256'hc2f111f16bf0a8ef26efdeeec9eeb5eeebee1bef2aef1defe0ee7dee05ee93ed;
    decBuf[1345] = 256'h0eedd9ecc8ecd7ec35ed8aededed4aee6fee64ee32eee0ed7ded3aed15ed20ed;
    decBuf[1346] = 256'h8eedf6ed89ee39efb0eff1ef05f0cfef9eef54ef2cef08ef29ef6fefc1ef24f0;
    decBuf[1347] = 256'h67f08bf080f04ef0fcefc5ef7fef64ef7defa2efe0ef3bf077f098f0b6f0adf0;
    decBuf[1348] = 256'ha5f0acf0c1f0f9f06af1fcf185f226f3bef320f49df4cef4faf422f546f593f5;
    decBuf[1349] = 256'hedf542f6bbf62df794f7d7f72cf84df87ff888f880f878f872f85ff84ef853f8;
    decBuf[1350] = 256'h4ef85bf87ef88cf8a1f8b5f8aaf894f886f85ef842f83df82ff83cf85ff876f8;
    decBuf[1351] = 256'h94f8aff8c0f8d0f8e4f8f7f811f945f96bf9a9f9e2f917fa2bfa4bfa3afa2afa;
    decBuf[1352] = 256'h1dfafff9ebf9e8f9e5f9e8f9f0f9e4f9d1f9b4f981f951f919f9d5f896f85cf8;
    decBuf[1353] = 256'hfaf79df730f7c8f66bf616f6dff5c1f5caf5c2f5baf598f553f501f59ef426f4;
    decBuf[1354] = 256'hb4f36af35df381f3cef328f495f41af573f5a4f5b3f5a5f599f58ef584f58df5;
    decBuf[1355] = 256'hc7f50bf65df6d6f627f78ef7d1f70ef819f837f81bf813f81bf814f81af836f8;
    decBuf[1356] = 256'h50f879f8a1f8baf8dbf8f0f803f915f931f94cf973f9a1f9c0f9f3f907fa1afa;
    decBuf[1357] = 256'h20fa1bfa16fa2bfa46fa7bfacdfa30fb8efbfbfb62fca5fccafcd5fcdffce8fc;
    decBuf[1358] = 256'hf0fc15fd53fdaefd1bfe82fefbfe4cffb3ffdbffe8ff0900130040007a00ae00;
    decBuf[1359] = 256'h08015d01aa01f0011d0247025d028d02ac02f6025003a40307048004d1041b05;
    decBuf[1360] = 256'h430567058805ce050e06690607079e074f08f508b7093a0ab10af20a540b890b;
    decBuf[1361] = 256'h9a0be30b410cae0c330dd40d400ec90e460f980fa60fb40f8f0f840f660f4b0f;
    decBuf[1362] = 256'h640f980fc80f26109f10cf1037115f11531148112a11fc10f4100a111f117011;
    decBuf[1363] = 256'hd3114b12bd1242139b13ed13191441147e149f14d11423158615c9154e16a716;
    decBuf[1364] = 256'hf9166017a317c717fe1730184b188518ba18c118ec18f218ce18c01891184018;
    decBuf[1365] = 256'h0918d71797177f176817381725170917c61699165f160d16d615a41576158f15;
    decBuf[1366] = 256'ha515ba15ff153e166816ab16d916e116f816f116d116cc16bc16a516bb16d616;
    decBuf[1367] = 256'he716161738173f1744171617b8165b16d5155815e71462140814d813ab136913;
    decBuf[1368] = 256'h44130d139f1238128a11b4102510390f5c0ecc0d150d9f0c5e0c230ced0bbd0b;
    decBuf[1369] = 256'h900b330bc60a410aa00909097f08de079d073b070607160707072f0754074907;
    decBuf[1370] = 256'h3f073607eb06910624069f052205b1042c04d20381033703f502d00299025302;
    decBuf[1371] = 256'hef015c01ab00d5ff0cff21fe44fdb4fcfdfb86fb45fb0afbf9fac8fa7efa3bfa;
    decBuf[1372] = 256'hcef967f9eef85cf8faf77df72cf7e2f69ff67bf670f666f65df665f66cf673f6;
    decBuf[1373] = 256'h86f675f647f61bf6d2f58cf54cf502f5e4f4dbf4e3f409f539f558f55ef56df5;
    decBuf[1374] = 256'h56f527f508f5caf490f46bf448f429f40df4f3f3dcf3d8f3ccf3d0f3ecf3fff3;
    decBuf[1375] = 256'h18f43af448f444f438f412f4e4f3d1f3c0f3c5f30af450f4c7f439f5a0f5fef5;
    decBuf[1376] = 256'h53f674f67ef699f680f688f68ff688f6a4f6bef6def6fcf627f743f767f790f7;
    decBuf[1377] = 256'h96f79bf797f779f746f716f7c5f68ef670f667f680f6b4f600f75af7aff7e6f7;
    decBuf[1378] = 256'h18f821f819f811f818f812f823f851f889f8dbf828f96ef9aef9f9f917fa44fa;
    decBuf[1379] = 256'h6dfa93faa8fac7fac1fabcfab7fa9afa77fa69fa5cfa58fa6afa6dfa70fa6dfa;
    decBuf[1380] = 256'h4afa07fac7f95cf9f5f897f82af8e0f7b8f794f75df73ff711f7d7f6a3f665f6;
    decBuf[1381] = 256'h2bf615f600f6faf50bf605f60af617f613f616f626f629f636f650f654f65df6;
    decBuf[1382] = 256'h66f659f651f654f64ef656f66ff680f696f6b0f6acf697f66bf627f6e7f59df5;
    decBuf[1383] = 256'h6bf54ff557f56ef59ef5d6f5edf501f6eff5bcf57ef534f5daf49df47cf472f4;
    decBuf[1384] = 256'h8ef4c7f40bf56ff5cdf522f685f6c8f6ecf623f741f74af763f788f7b9f70af8;
    decBuf[1385] = 256'h83f8f5f879f91afa86fa10fb69fb9afba9fbb6fbaafbb5fbbffbc8fbe1fb15fc;
    decBuf[1386] = 256'h45fc7efcb2fce2fc0efd35fd59fd83fdaafdcefde5fdfafdfefd02fefffd07fe;
    decBuf[1387] = 256'h29fe5cfea8fe16ff7dfff6ff6700cf002c0169018a01a801c301ec0112025e02;
    decBuf[1388] = 256'hb80225038c03ea035704a004e30438056f05a105e1051b06400670069c06b806;
    decBuf[1389] = 256'hd206e906070731076407a207ec0746089b08e8082e095c0974096d0958092d09;
    decBuf[1390] = 256'hfa08ca08ab08a508b408f0083b098109e509280a340a3f0a0d0abb096e091409;
    decBuf[1391] = 256'hbf089e08a808d60830098509e8092b0a500a450a270ae7098c094f090209d008;
    decBuf[1392] = 256'hb508ad08a5089e08a508940899088b087e088a0886087d0886087e0868085a08;
    decBuf[1393] = 256'h3d081a08160811081d084a088308c608060950096e099c0994098c0978096509;
    decBuf[1394] = 256'h3d0938092a0926093a094b095b0975098d09900993098609670949091709d908;
    decBuf[1395] = 256'hb0086c083f080508df07af0784075c0738070f07e706b9068d065b062b06ff05;
    decBuf[1396] = 256'hcc058e0555051105bf04880456042804100408040f042204270422041e04f703;
    decBuf[1397] = 256'hc90385034503fa02b40275023b0224020202fc01eb01d101b10182013d01eb00;
    decBuf[1398] = 256'h720000007cffdbfe43febafd61fdeffc88fc45fcf0fbcffb89fb49fbeefa99fa;
    decBuf[1399] = 256'h0afaa8f907f99bf839f8e0f78ff762f755f761f76cf776f77ff777f760f723f7;
    decBuf[1400] = 256'he9f696f633f6d6f581f534f516f5faf4f2f4faf40ef515f51af50bf5e1f4baf4;
    decBuf[1401] = 256'h6df420f4eef39cf365f347f32bf323f33af333f346f356f351f356f363f34ff3;
    decBuf[1402] = 256'h3ef32ef303f3d7f2bbf297f280f27cf278f28af2b2f2cef2e8f212f32ef33df3;
    decBuf[1403] = 256'h5df362f36df37ff375f378f385f37ef389f3a3f3b4f3ddf31bf455f498f4eaf4;
    decBuf[1404] = 256'h21f53ff56df565f55df549f529f524f529f537f55df595f5caf508f652f684f6;
    decBuf[1405] = 256'hc4f6edf604f718f71ef702f7e9f6d2f6abf69cf6aaf6b7f6e1f62af770f7c2f7;
    decBuf[1406] = 256'h0ff841f86ff888f871f85df83df816f811f81ff83df877f8c1f807f959f9a6f9;
    decBuf[1407] = 256'hd8f906fa2ffa45fa4cfa46fa35fa1cfa04fadef9d9f9e7f9fcf936fa91fae6fa;
    decBuf[1408] = 256'h33fb8dfbcafbebfbe1fbc5fbacfb78fb56fb36fb3cfb4bfb75fbbefbf0fb30fc;
    decBuf[1409] = 256'h6afc80fc87fc81fc59fc2bfc00fccdfb9dfb7efb56fb47fb4bfb47fb5bfb6cfb;
    decBuf[1410] = 256'h6ffb6cfb64fb41fb1dfbfdfad6fabdfaaffaa2faa6faa2fa99fa90fa83fa73fa;
    decBuf[1411] = 256'h68fa72fa89fab1faeffa3afb80fbbffbe9fbf0fbf7fbe4fbdffbdafbf1fb28fc;
    decBuf[1412] = 256'h7afcddfc56fde8fd4afea4fed4fe01ff29ff35ff2aff20ff29ff31ff48ff5cff;
    decBuf[1413] = 256'h95ffc9ff15005b009b00c400f8000d010701eb00d1009e007c00690063007d00;
    decBuf[1414] = 256'hb000ee004801b601ff015d02b202e902070334033d03440359036c039e03dc03;
    decBuf[1415] = 256'h26049404fc04740506066806c20613073f0732073e07490753078107ba070d08;
    decBuf[1416] = 256'h7008cd0822099b09ed09360a790ace0a050b4b0b8b0bb40bda0b0a0c1d0c440c;
    decBuf[1417] = 256'h5e0c750c9b0cde0c0b0d660dbb0d080e760ec00ee80e0c0f2d0f230f1a0f220f;
    decBuf[1418] = 256'h0c0f200f4c0f730fc00f3910ab103011ad11de1145126d12611256123812f811;
    decBuf[1419] = 256'hf011e811e1111a126c12cf124813b91303144614831478146e144014f613d813;
    decBuf[1420] = 256'haa1381139713ba13d9132d149a14e4145d15ae15bd15ca158d152a15cd146014;
    decBuf[1421] = 256'hf813b513a9139e13f81335148214dc140015f514d71497142c14e21385133013;
    decBuf[1422] = 256'hf912db12c012e912ff1206133e1355135c13621351130f13cf1284121612cd11;
    decBuf[1423] = 256'h8a114d114211381154116c1183117c1169112b11d11094103110ee0fb10fa60f;
    decBuf[1424] = 256'h880f7f0f770f520f2f0fea0e980e350ed80d830d4c0d1a0dec0cd30c9f0c610c;
    decBuf[1425] = 256'h270cd50b720b140ba70a220ac9095709f008ad08700839081b0812080a081208;
    decBuf[1426] = 256'hef07b70773070f0797062506a0052305f204c604d304f8041905370552053905;
    decBuf[1427] = 256'h1405d6046b04e6036903f70272021902e801bc01af01a3019801a20186015d01;
    decBuf[1428] = 256'h1901a300110087ffc3fe0cfe65fdcefc6cfc36fc06fcd9fbccfba8fb71fb2bfb;
    decBuf[1429] = 256'hb4fa22fa98f9f7f88bf802f8a9f757f72bf71ef712f707f7fdf6f3f6ebf6e4f6;
    decBuf[1430] = 256'hcff6b0f688f665f628f6eff5baf58af552f52cf518f505f50bf505f513f520f5;
    decBuf[1431] = 256'h24f512f5f6f4bcf461f40df4aaf34cf3f7f2c0f2a2f2bdf2e7f20cf358f376f3;
    decBuf[1432] = 256'h7ff387f353f315f3dbf289f252f234f218f220f255f277f2a3f2e1f20af330f3;
    decBuf[1433] = 256'h60f366f377f391f38cf390f394f38af38df3acf3c2f3fcf356f4abf4f8f466f5;
    decBuf[1434] = 256'hb0f5d8f5fdf5f2f5d4f5a6f56cf556f54ff555f571f5b4f5e1f52cf672f69ff6;
    decBuf[1435] = 256'hc9f6dff6caf6b8f69cf66df64ef649f639f65af699f6d9f623f77df7a2f7c3f7;
    decBuf[1436] = 256'hcdf7b1f788f754f708f7d6f6cdf6c5f6dbf60bf72bf747f760f75cf757f74cf7;
    decBuf[1437] = 256'h2cf720f714f702f7f3f6f0f6def6d2f6d4f6cef6d7f6eff607f72af74af757f7;
    decBuf[1438] = 256'h4bf73af70bf7dbf6a3f67df668f67bf697f6daf61af754f779f78ef76ef73cf7;
    decBuf[1439] = 256'h0cf7c7f699f691f699f6bbf6f3f637f777f7a0f7b6f7aff790f75ef720f7e6f6;
    decBuf[1440] = 256'hb1f68ff695f6a6f6caf606f72ff764f779f772f761f73ef701f7c8f6a2f68ef6;
    decBuf[1441] = 256'h94f6b0f6e8f62cf790f7d3f728f85ff87df886f88ef878f871f884f895f8b8f8;
    decBuf[1442] = 256'hfef858f9c5f92cfa8afadffa16fb48fb51fb49fb41fb3afb40fb51fb7ffbc4fb;
    decBuf[1443] = 256'h04fc5ffcb4fcebfc1dfd26fd2efd27fd20fd0dfd07fd17fd2efd54fd97fdd7fd;
    decBuf[1444] = 256'h21fe67fea7fee0fe06ff28ff54ff65ff7fffa8ffdbff19007300e1004801a501;
    decBuf[1445] = 256'hfa01470279029502ad02c402d902f8022a037603bc030e044504770493049b04;
    decBuf[1446] = 256'h840470045d04570467047e04a404c804df04f404f804ee04e404dc04cf04cc04;
    decBuf[1447] = 256'hd304d504e104ec04ee04f704fb0405051a05340553058205a105bd05cd05db05;
    decBuf[1448] = 256'hce05d205ce05d105f105170645067e06b206c706e606e006c706b00689065b06;
    decBuf[1449] = 256'h3c06200606060206fd05010605060e060506fe05e305b6057e053a05e8049b04;
    decBuf[1450] = 256'h69043b0444044b047b04b404d904ee04f404c10476041c04af0347030403e002;
    decBuf[1451] = 256'hd502070322035c038203890369033703eb0291023c02d9019601720167015d01;
    decBuf[1452] = 256'h66015e0165016c01590149011a01e2009f005f001500e3ffa3ff8aff73ff6dff;
    decBuf[1453] = 256'h66ff6cff67ff50ff32ff07ffd5fe97fe5dfe38fe15fe02fefdfdf8fdeafdddfd;
    decBuf[1454] = 256'hc2fd9bfd6dfd42fd0ffddffcb3fc97fc73fc65fc50fc35fc1cfcfafbc7fb97fb;
    decBuf[1455] = 256'h5ffb1bfbdbfa91fa4bfa1dfaf4f9def9e5f9f7f9fdf90cfa08faeaf9bff976f9;
    decBuf[1456] = 256'h1cf9e0f893f861f845f84df864f886f8b2f8cef8e8f8daf8b4f890f84af8f0f7;
    decBuf[1457] = 256'hb4f767f735f707f7fff606f71bf73af762f790f796f790f76df727f7cdf678f6;
    decBuf[1458] = 256'hfff5aef582f55af566f587f5a5f5d2f50cf605f6f0f5d1f588f542f502f5b8f4;
    decBuf[1459] = 256'h86f47cf464f47af49df4c8f4f0f428f54ef562f581f571f557f52df5fbf4cbf4;
    decBuf[1460] = 256'habf49af4a0f4c0f4def408f530f53ff531f51cf5e2f4a8f483f452f44cf45df4;
    decBuf[1461] = 256'h62f479f497f493f482f46cf441f421f41cf421f438f478f4a5f4dff405f519f5;
    decBuf[1462] = 256'h13f502f5def4d0f4d5f4e0f40ef546f58af5c9f503f629f64bf66af67bf69ff6;
    decBuf[1463] = 256'hc9f6e5f609f729f736f749f762f771f791f7c8f70cf84cf8a6f8e3f81af938f9;
    decBuf[1464] = 256'h41f928f912f9eff8e9f8faf814f947f992f9c4f904fa3efa72fa95fab4fabafa;
    decBuf[1465] = 256'hd3faeafaf7fa0afb23fb39fb5efb97fbdafb2cfc8ffcedfc42fd8ffdadfdb6fd;
    decBuf[1466] = 256'h9dfd69fd46fd40fd46fd7efdd0fd33feacfefdfe29ff51ff45ff24fff2fee9fe;
    decBuf[1467] = 256'he1fe06ff44ff8fffe9ff3d008a00bc00ea00030119012e014d0175019801c201;
    decBuf[1468] = 256'hf501250251028302b302f802380361038703a903af03aa03a503a003b503e003;
    decBuf[1469] = 256'h1e046804c2041705640582058b0572056b0556055c058405bc050f068806d906;
    decBuf[1470] = 256'h40078307c007e107ff070808310856087908be08fd0837098a09d7091d0a6f0a;
    decBuf[1471] = 256'hd20a150b6a0bb70be90b280c410c490c5d0c700c810caf0cf40c340d8e0de30d;
    decBuf[1472] = 256'h1a0e4c0e680e5f0e670e6e0e4f0e540e4f0e410e4e0e5a0e5d0e860ead0edb0e;
    decBuf[1473] = 256'h130f480f6a0f8a0f8f0f760f710f5c0f410f4b0f670f920fe60f3b107210b810;
    decBuf[1474] = 256'he610ee10f510ef10cf10ca10c510b710d410e010e410f310f610e910f510ff10;
    decBuf[1475] = 256'hfd1018111c1111110811e810b1108b105b103c1036103b1037105d1062105410;
    decBuf[1476] = 256'h50102d10fa0fd80fac0f850f800f7b0f6e0f7a0f6f0f4d0f3f0f2a0f070f0c0f;
    decBuf[1477] = 256'h180f1c0f3c0f490f450f410f2b0f000fe10ed00ec10ed80ee50ee80e010ff80e;
    decBuf[1478] = 256'hd20eae0e7b0e3e0e250e0e0efa0d000e060eec0dd50da60d550d1e0dd80caa0c;
    decBuf[1479] = 256'h910c8a0c830c890c8f0c800c720c540c220cff0bec0bd00bd50bd10bcd0be00b;
    decBuf[1480] = 256'hdc0bcd0bd00bd20bd50bf50b1e0c3a0c680c6f0c530c390cfd0bc30b9e0b890b;
    decBuf[1481] = 256'h8f0bb70bef0b140c370c3d0c0a0cda0b890b260bfe0ac10ab60aac0ac80abf0a;
    decBuf[1482] = 256'hc70aa50a790a460a080acf09b809b1099e09a40995096b093809fb08b0087e08;
    decBuf[1483] = 256'h510838083f0846084d08520843082208fc07c407800740070707d206b0067806;
    decBuf[1484] = 256'h43060506cb0588055a052105fb04d904a0046c042e04c3035c03e30271020a02;
    decBuf[1485] = 256'hc7018b016a014c0143013a012401f400c8008a0040000e00ceff84ff3efffefe;
    decBuf[1486] = 256'hb4fe5afe1dfed0fd9efd83fd6afd71fd5dfd3dfd00fda5fc1ffc7ffbe7fa37fa;
    decBuf[1487] = 256'hc0f954f919f907f917f908f9fbf8bef871f817f892f715f783f6f9f57cf52bf5;
    decBuf[1488] = 256'he1f49ef47af459f43bf444f43cf425f41ef4fff3d8f3b4f381f343f31af303f3;
    decBuf[1489] = 256'heff202f31ef342f37ef3a7f3dbf3fef304f4fef3f9f3e2f3bcf3a2f379f351f3;
    decBuf[1490] = 256'h2df30df3eff2ebf2e8f2ebf20bf317f31bf31ff3f6f2c4f293f242f20bf2edf1;
    decBuf[1491] = 256'hc0f1b7f1cef1e2f102f229f22ef23cf251f246f242f24cf249f251f26bf267f2;
    decBuf[1492] = 256'h71f27ff272f279f290f29af2bff2edf20cf334f358f35cf361f35df344f33bf3;
    decBuf[1493] = 256'h38f326f323f32ef324f322f324f313f30df317f319f327f345f352f365f370f3;
    decBuf[1494] = 256'h66f352f340f321f314f320f338f367f3cef336f4aef420f587f5caf507f63ef6;
    decBuf[1495] = 256'h5cf689f6b2f6e7f633f779f7cbf744f895f81af973f9c4f92cfa54fa60fa55fa;
    decBuf[1496] = 256'h37faf7f9cef9b7f995f99bf9b7f9d1f9faf917fa26fa18faf2f9aff96ff925f9;
    decBuf[1497] = 256'hdff8b1f8a9f8a2f8c4f8e3f80bf91af928f91bf908f9eff8d3f8c8f8c4f8c7f8;
    decBuf[1498] = 256'hdbf803f92af958f984f9b7f9e7f906fa22fa31fa36fa29fa1efa1afa1dfa37fa;
    decBuf[1499] = 256'h6cfaaffaeffa4afb86fba7fbb1fb96fb5cfb0afbbdfa8bfa82fa8afacdfa32fb;
    decBuf[1500] = 256'h8ffbfdfb64fca7fccbfcecfce2fcd9fce1fce9fc0bfd50fda2fd05fe7dfeeffe;
    decBuf[1501] = 256'h74ffcdff3f008900e6000b0116010c01f000c700b1008e0088009900b200e500;
    decBuf[1502] = 256'h23014c017201790166013301f6009b004600f9ffc7ffacffb4ffbbffdefffdff;
    decBuf[1503] = 256'h2400480072008e009d00ab00af00ac00a800a500a800bf00e2001e016801ae01;
    decBuf[1504] = 256'h00026302a602e3021a03380365037e0386039a03ad03a703a20394037f036403;
    decBuf[1505] = 256'h530349034c035e0374038e039f03960376033f03ec0289022c02d701a0018201;
    decBuf[1506] = 256'h8b01a401d80116023f02650287028e02880279026102440229020902f401e801;
    decBuf[1507] = 256'hec01fb0121024f027b02ad02d002d602c5028d023a02d70179010c01a5006200;
    decBuf[1508] = 256'h3e00490053005c0075008b00840072004a001200ceff8eff44ff12ffe5feccfe;
    decBuf[1509] = 256'hc4fee7fe12ff50ff8affceff0d0037003e004500320021001c00210036005900;
    decBuf[1510] = 256'h9500cf00210158018a01a601bf01d501ce01c801c201a9019201740149010b01;
    decBuf[1511] = 256'hd2008e003c000500bfff91ff58ff32fff4feaafe64fe12fec5fd7ffd2dfdf6fc;
    decBuf[1512] = 256'hb0fc82fc59fc24fc02fceffbeafbf9fb19fc40fc6efca6fccbfce0fce6fccafc;
    decBuf[1513] = 256'hb1fc90fc72fc67fc71fc9afcd8fc33fd87fdd4fd1afe36fe4ffe47fe32fe07fe;
    decBuf[1514] = 256'hdffdbbfd9bfd8efd92fda4fdc6fdf9fd29fe61fe87fe9bfe95fe6efe2bfed9fd;
    decBuf[1515] = 256'h8cfd46fd18fd10fd27fd57fd8ffdd3fd12fe2bfe33fe1efef2fdcbfda7fd87fd;
    decBuf[1516] = 256'h7afd7efd88fd98fdacfdaffdacfda2fd84fd66fd43fd10fde0fcb4fc76fc3dfc;
    decBuf[1517] = 256'h08fccafb91fb5cfb3afb0efbf2fac4fa98fa65fa35fafdf9d7f9c3f9bdf9c2f9;
    decBuf[1518] = 256'hdcf9fcf922fa32fa40fa44fa31fa2dfa2afa33fa4ffa7afab8fa02fb5cfbb1fb;
    decBuf[1519] = 256'hfefb44fc84fcbefcf2fc15fd34fd39fd3ffd3afd3efd42fd5bfd83fdc1fd0bfe;
    decBuf[1520] = 256'h65febafef1fefbfee0fea6fe36fec4fd5dfdfffcc2fccdfcebfc2bfd86fddbfd;
    decBuf[1521] = 256'h12fe44fe3bfe22fedefd8cfd3ffde5fcc1fca0fcbefcecfc36fd90fdfdfd47fe;
    decBuf[1522] = 256'ha4fee1feecfef6fedbfeb1fe8cfe5cfe49fe4ffe5efe7efeb6feeafe28ff51ff;
    decBuf[1523] = 256'h86ffa8ffc7ffcdffd2ffcdffc1ff9eff7dff4fff23ff12ff0dff24ff5bffaeff;
    decBuf[1524] = 256'h11006e00c300fa002c012301fa00d400a40085008b00af00f4006201e7016402;
    decBuf[1525] = 256'hd6023d039a03d703f80316041f0427042f0436043c044d0467048704a504d704;
    decBuf[1526] = 256'h0705330566058805a705ad059305730544050c05c8049b0461044a0444044a04;
    decBuf[1527] = 256'h7c04ba0405055f05b305000632064e06560640061d06fe05f805080631068606;
    decBuf[1528] = 256'h0b07ac074308f4086b09020a3d0a4f0a3f0a300aed09c909a8099e09b909030a;
    decBuf[1529] = 256'h710ad80a6c0bce0b270c370c290ce60b790bd60a6a0ae1098709570948097009;
    decBuf[1530] = 256'had09fa09180a330a2b0af609ab095109e4089a0857083308540872089f08d908;
    decBuf[1531] = 256'h1c093809510967096009730979097e099509aa09b609c009bd09a90997097809;
    decBuf[1532] = 256'h510942093409270933094c095b0975098709770963093b09f208ac086c082208;
    decBuf[1533] = 256'h0408e907f107170847087f08c208f008190921091a09ee08d2089a0865085108;
    decBuf[1534] = 256'h4a08450869089b08d90824096a09a909e309eb09e409c50987092c09d7087408;
    decBuf[1535] = 256'h1608f207d107c707e207eb0701080808e907ab075007cb064e06bb055905dc04;
    decBuf[1536] = 256'hab047f048d049904ba04c404df04e704d104ca04ab04830474045d0450046304;
    decBuf[1537] = 256'h75048504aa04c404d104e704f20404051a0528053a0550055805510549052e05;
    decBuf[1538] = 256'hfb04cb04870447040d04e703c503bf03c403ca03d703d303b8038b034603f402;
    decBuf[1539] = 256'h91023302de01a70175015a01520159017b019b01b701c601dd01d901d501bd01;
    decBuf[1540] = 256'ha1017e015d014001240121012401380160019201c201fb01110226021302ec01;
    decBuf[1541] = 256'h9f015201e4007c003a00e5ffc4ffbaffc3ffdcfff2ff07000000f0ffadff5bff;
    decBuf[1542] = 256'hf8fe9afe2dfee3fda0fd7cfd87fda5fdc0fdfafd2ffe51fe57fe52fe38fe0efe;
    decBuf[1543] = 256'hdcfdacfd80fd64fd54fd59fd66fd79fd8bfda1fda9fda7fd9bfd7ffd54fd22fd;
    decBuf[1544] = 256'hf2fcc6fc88fc5ffc39fc17fcf8fbdcfbb8fb97fb71fb43fb17fbe5fab4faa2fa;
    decBuf[1545] = 256'h86fa6cfa5efa51fa3efa25fa09fae6f9cff9baf9aef9b2f9cef9f1f92dfa77fa;
    decBuf[1546] = 256'hbdfafdfa37fb5cfb71fb84fb7efb6ffb6afb66fb6afb82fbb1fbeffb39fc7ffc;
    decBuf[1547] = 256'hbffcf9fc1efd33fd20fd04fdd6fc9efc69fc47fc34fc3afc53fc7dfcbbfcf5fc;
    decBuf[1548] = 256'h38fd54fd6cfd65fd42fd17fdcefc88fc48fc0efce8fbeffb02fc35fc80fcc6fc;
    decBuf[1549] = 256'h06fd2ffd37fd15fde9fc94fc40fcddfb9afb5dfb52fb5cfb8afbd4fb06fc46fc;
    decBuf[1550] = 256'h6ffc77fc54fc1cfcd8fb74fb31fbdcfabbfa9dfaa6fad0fa04fb50fb96fbd6fb;
    decBuf[1551] = 256'hfffb06fc0dfcfbfbdefbc5fbaefbb2fbc5fbe5fb1cfc60fc9ffcd9fc0efd30fd;
    decBuf[1552] = 256'h43fd54fd4ffd4afd46fd42fd3efd48fd45fd47fd4afd3ffd35fd33fd2bfd27fd;
    decBuf[1553] = 256'h30fd34fd3afd41fd35fd24fd09fdd5fca0fc70fc2cfcecfbc2fb9dfb96fb9cfb;
    decBuf[1554] = 256'ha2fbb1fbc8fbc4fbb9fb99fb62fb1efbdefa84fa47fa26fa08fa11fa2afa5efa;
    decBuf[1555] = 256'h81faadfac9facefac9faabfa81fa59fa36fa15fa08fa05fa16fa38fa62fa89fa;
    decBuf[1556] = 256'hc2faf6fa19fb44fb55fb65fb69fb5dfb49fb3ffb2ffb32fb44fb63fb9afbedfb;
    decBuf[1557] = 256'h3afc80fcd2fcf3fc11fd1afd01fddcfcbafc9afc89fc84fc92fcb8fcf1fc25fd;
    decBuf[1558] = 256'h55fd9afdb6fdcefdd6fdcffdbcfda0fd86fd66fd59fd4efd58fd68fd82fdaffd;
    decBuf[1559] = 256'hdbfd0efe4bfe75fe9afebdfec3fec8feb9fe99fe7bfe58fe41fe34fe38fe5ffe;
    decBuf[1560] = 256'h97fedafe3fff82ffbefff5ffebffd0ff86ff2cffd7fea0fe6efe77fea0fef3fe;
    decBuf[1561] = 256'h6cffddff4500a200df00ea00cc008c0052000000c9ffabffa2ffcbffffff5900;
    decBuf[1562] = 256'hc6002d018b01e001170221021802ee01ba0160012401ed00cf00c600ef003201;
    decBuf[1563] = 256'h8501e8012a026702720254021402b9014c01c8004a00f9ffafff87ff93ffb4ff;
    decBuf[1564] = 256'he6ff14003d0063005c003d00ffffb5ff5bffedfea4fe7cfe57fe62fe94fed4fe;
    decBuf[1565] = 256'h1eff78ffcdff0400360052005a0052003e001e00f7ffddffd0ffd4ffe7ff1500;
    decBuf[1566] = 256'h5900ac000f016c01c101f8010202e701ad015a01f700b5007800570061008f00;
    decBuf[1567] = 256'hc8000c01390163015b012b01e60082002400cfff98ff66ff5dff66ff7cff91ff;
    decBuf[1568] = 256'ha3ffb4ffafffabff95ff7aff69ff5fff57ff59ff5cff55ff4bff38ff1bfff1fe;
    decBuf[1569] = 256'hc9fe9bfe7cfe76fe7bfe92feb0fedbfef7fe11ff03ffe5feabfe61fe1bfedbfd;
    decBuf[1570] = 256'hb1fdaafdbffdeafd33fe79feccfe03ff35ff3eff35ff1fff0afff8fee7feecfe;
    decBuf[1571] = 256'hfafe0fff32ff5bff8effccff16005c009c00e600180134013c012501f500bd00;
    decBuf[1572] = 256'h7a003a00210019002e005a00a300e90017012f012801f8009a003c00b7ff3aff;
    decBuf[1573] = 256'he9fe81fe59fe4dfe58fe76fea4feddfe03ff18ff1eff0dffdffea7fe63fe23fe;
    decBuf[1574] = 256'he9fdb5fda0fda7fdcefdfcfd41fe93fee0fe12ff40ff58ff60ff4bff1fffedfe;
    decBuf[1575] = 256'haffe75fe50fe3bfe4efe75feb8fe0aff6dffcbff07003e0048002d00f3ffb0ff;
    decBuf[1576] = 256'h70ff36ff10ff0aff1cff4fff9bfff5ff49009600c800f600fe000601e300c400;
    decBuf[1577] = 256'h9200610036000e00f5fff9ff170049009500ef0044019101af01b8018f014b01;
    decBuf[1578] = 256'he7006f00fdff96ff53ff2eff39ff57ff97ffd1ff05001a001400ecffb4ff62ff;
    decBuf[1579] = 256'hfffea1fe4cfe15fe0bfe02fe1bfe4ffe7ffed1fe08ff4eff8dffa6ffbdffd1ff;
    decBuf[1580] = 256'hcbffbaffabff94ff87ff8bff8effa4ffcfff14006600c90027019401de012102;
    decBuf[1581] = 256'h450250023202e00193014d011f0106011d015b01c6012d02c00223037c038c03;
    decBuf[1582] = 256'h60031d0398021b028801ff00a60075008400ac0001014e01bc01050248025402;
    decBuf[1583] = 256'h3302ed01890111019f003800f5ffd0ffdbff21008600fe007001d7011a023e02;
    decBuf[1584] = 256'h1d02eb0199013601d9006b003f00170023005a00b4002101a60123027402be02;
    decBuf[1585] = 256'he602f202bb0275021102b3017701560160018d01e8016e02eb025c03c403ec03;
    decBuf[1586] = 256'hf803d70391032d03cf027a024302390242026b02af0201036403c20317044e04;
    decBuf[1587] = 256'h6c0475045c042704ea039f0359032c030203fb021d0349039203d80318044104;
    decBuf[1588] = 256'h49043404fc03b80354031103bc02850267025e0277029c02da0225036b039803;
    decBuf[1589] = 256'hb103c703b303940361032303e902c402af02a902c502f3021f03520374039303;
    decBuf[1590] = 256'ha403a9039b039703930390038d038f0388038a03880386039203a403be03ec03;
    decBuf[1591] = 256'h17043f046d0480048504760455042704fb03c80398038503800370037e038303;
    decBuf[1592] = 256'h8e039903a803b103b903c003be03b803a80388035f0337031303f302e602ea02;
    decBuf[1593] = 256'h0a03380364039703c703da03ea03d103a70369031f03d902990270024a024402;
    decBuf[1594] = 256'h4a0266029402cc02f2022203350324030a03ce0284023e02fe01c401ae01b501;
    decBuf[1595] = 256'hd40112024b028f02bd02e602ed02e602c702a00267022402e401bb0195018e01;
    decBuf[1596] = 256'h9501b101e9012d027f02b602fc020503fd02d7028c023202dd0190015e015501;
    decBuf[1597] = 256'h5d018201b201de0106020b02fd01d7019e015b011b01d1009f005f0046002000;
    decBuf[1598] = 256'h0c00f9ffffff180039005f009700cc00ee000d011301f900d900b30085005900;
    decBuf[1599] = 256'h48004d006e00a500e80028017201b801e601ee01d801b5017d012b01de009800;
    decBuf[1600] = 256'h6a00620069008c00c400f8002901480142011e01e20098003e00e9ff86ff5eff;
    decBuf[1601] = 256'h21ff00fff6feedfee5feddfed7fed0fed6fed1fed5fed1febefe97fe69fe24fe;
    decBuf[1602] = 256'he5fdabfd94fd8dfda0fdd3fd1efe78feb5feecfe0aff01ffc7fe93fe47fe01fe;
    decBuf[1603] = 256'hd3fdbbfdc2fde5fd1dfe60fea0fec9fefefe13ff19ff13fffafee2fecdfebafe;
    decBuf[1604] = 256'haffeacfebbfed2fef5fe1eff46ff69ff8affa8ffbbffbeffc2ffbfffb7ffabff;
    decBuf[1605] = 256'h98ff85ff75ff66ff60ff5eff6aff80ffa9ffd0fff4ff0b000f00fcffd5ff9dff;
    decBuf[1606] = 256'h5aff1affe0fec9feb5fec8fee4fe08ff1fff2bff28ff0fffe6feb4fe91fe72fe;
    decBuf[1607] = 256'h61fe5cfe6afe7ffe9afeacfebcfecafecdfed4fed6fed8fedafedbfeddfedefe;
    decBuf[1608] = 256'hdffee3fee4fee5fee9fef1fef4fef7fefafefbfefcfefefe01ff0eff24ff38ff;
    decBuf[1609] = 256'h55ff70ff7bff84ff81ff74ff68ff59ff4bff49ff4bff56ff62ff71ff77ff78ff;
    decBuf[1610] = 256'h7aff6fff66ff62ff5cff59ff59ff54ff53ff4fff47ff41ff42ff47ff50ff65ff;
    decBuf[1611] = 256'h79ff8cff97ff9eff94ff81ff64ff41ff17fff0feccfeacfe8efe7afe70fe60fe;
    decBuf[1612] = 256'h5dfe5bfe54fe52fe4cfe3ffe2afe0bfee4fdb6fd8afd63fd54fd58fd6efd90fd;
    decBuf[1613] = 256'hc3fde6fd05fe0bfe05fee5fdb6fd7efd59fd36fd23fd29fd38fd59fd7ffda3fd;
    decBuf[1614] = 256'hbafdc7fdd2fdcffdccfdcffdd7fddefdedfdfffd0ffe22fe35fe45fe58fe66fe;
    decBuf[1615] = 256'h71fe80fe8afe90fe98fe99fe98fe94fe8afe78fe63fe43fe1dfef9fdd9fdc3fd;
    decBuf[1616] = 256'hb8fdbbfdc5fddefdf7fd07fe15fe08fef2fdcdfd9ffd73fd57fd3dfd42fd57fd;
    decBuf[1617] = 256'h7afda4fdcbfde5fdf3fdf7fddcfdbcfd96fd72fd52fd45fd39fd44fd54fd68fd;
    decBuf[1618] = 256'h85fda0fdb8fdd4fdeffd01fe11fe19fe1cfe19fe1cfe1afe1bfe27fe34fe47fe;
    decBuf[1619] = 256'h5ffe6ffe77fe7ffe73fe5cfe46fe21fef3fdd3fda1fd7efd6cfd4ffd4afd46fd;
    decBuf[1620] = 256'h41fd4dfd58fd5bfd5efd5bfd4ffd3cfd2afd0ffdfefcf5fcf2fcfffc14fd28fd;
    decBuf[1621] = 256'h3bfd47fd3cfd26fd01fdd2fca7fc8bfc67fc62fc6ffc7afc9afcb8fccbfcddfc;
    decBuf[1622] = 256'he0fcddfcd0fcc9fcbefcc4fcd0fcdffcf9fc18fd2efd41fd52fd4ffd47fd34fd;
    decBuf[1623] = 256'h1afdfbfce5fccafcb2fca8fc94fc8cfc8afc84fc7afc7bfc77fc6ffc73fc77fc;
    decBuf[1624] = 256'h81fc93fca4fcb7fcc4fccbfcc5fcbffcabfc99fc8dfc82fc84fc94fca3fcb1fc;
    decBuf[1625] = 256'hc1fcbffcb5fc9afc68fc38fc0cfce5fbcbfbd0fbe5fb10fc42fc72fcabfcd0fc;
    decBuf[1626] = 256'he5fcdffccefcaafc89fc6cfc58fc55fc6bfc85fcabfcd9fc05fd21fd30fd35fd;
    decBuf[1627] = 256'h28fd15fdeefccbfcb3fc9efc9afcacfcc8fcebfc1efd40fd6cfd93fda3fda7fd;
    decBuf[1628] = 256'ha3fd9ffd95fd91fd89fd8bfd97fda2fdb4fdcefde0fdeffd03fe10fe1cfe27fe;
    decBuf[1629] = 256'h31fe3afe45fe4dfe53fe5cfe64fe73fe86fe99feb3fed2fef0fe13ff33ff51ff;
    decBuf[1630] = 256'h74ff82ff8eff9aff9eff8eff85ff7dff76ff70ff6eff70ff7bff89ff95ffa3ff;
    decBuf[1631] = 256'hadffb3ffaeffa3ff8fff75ff5cff40ff25ff1bff1eff2cff3eff5dff7bff96ff;
    decBuf[1632] = 256'hafffbeffc7ffc4ffb8ffaaffa0ff97ff98ffa3ffb5ffd4fffaff280047006f00;
    decBuf[1633] = 256'h9300a000ad00b100ae00a400a700aa00b100c800de0003012701480165018101;
    decBuf[1634] = 256'h8b018e018b017e01720163015d015c016101650171017d0184018b018f018e01;
    decBuf[1635] = 256'h8b0185017f017c017d017e018b019901a201b301bf01c601d001d101d001d401;
    decBuf[1636] = 256'hd301d401dc01e901f90110022602340247024e024802420235022a0228022f02;
    decBuf[1637] = 256'h3b02510273029402ba02d402e202e602e202d002c102ad02a0029d029f02ad02;
    decBuf[1638] = 256'hc102d802e802fc0209030b030903ff02ec02df02d302c802c602d302de02f502;
    decBuf[1639] = 256'h110324033d034c034f0357035503460340033a033203340338033c0344034703;
    decBuf[1640] = 256'h46034803470341034b035703660380039803ae03c203d503d703d503cf03c303;
    decBuf[1641] = 256'hbe03bf03c103d403eb0301042104360442044c04430429040904ec03c903b203;
    decBuf[1642] = 256'ha503a103b903d603f8032b044e046d047e0483046c04570434040a04f903e003;
    decBuf[1643] = 256'hdb03e803fb030d042f043d04410435042b040904e803c2039e03900383037803;
    decBuf[1644] = 256'h82039203a603c303e603fd031b04360439043c043a042c041c040d04ff03fa03;
    decBuf[1645] = 256'hfb0303041504250434043e04430438042e041e040804fa03ed03e103df03e903;
    decBuf[1646] = 256'hee03fa0304040804110419041604170416041104110411040a040404f903e503;
    decBuf[1647] = 256'hd803c303a3038e037b0362035f0368036a0380039403a103a803a60394038303;
    decBuf[1648] = 256'h68034d0342033f0342035f038203a203c003d303d703cd03b3038d0369034903;
    decBuf[1649] = 256'h2b031f031c032503330341033e033c032e031e030b03f902e802e602e802f102;
    decBuf[1650] = 256'hff0211031d032c032e032c0324031a030b03090307030c0319032d033f035003;
    decBuf[1651] = 256'h5a035403480330030903e502c502a70294029702ad02cd02f302210340035103;
    decBuf[1652] = 256'h4c033e032003f602ce02ab028a0286029202aa02c602e902090316031a030203;
    decBuf[1653] = 256'he502b30275023b021602e601e001e501f501150244026f028c029b02a0029302;
    decBuf[1654] = 256'h780251022d02160209020d0218022e024d0263026e0279026f0261024f023402;
    decBuf[1655] = 256'h1c020002ec01db01cb01c301b601b301b101b701b901c101cb01dd01e901f401;
    decBuf[1656] = 256'hf601f101df01c901af0197017b0167015d015a0157015a01650168016a016401;
    decBuf[1657] = 256'h590142012001f600da00b6009f009b009700a200ab00bf00cc00d300d100c700;
    decBuf[1658] = 256'hb4009700740054003f00240012000200f4ffecffe5ffd6ffccffc7ffbfffb4ff;
    decBuf[1659] = 256'hadffa5ff98ff86ff76ff63ff50ff44ff3eff40ff45ff54ff66ff77ff81ff87ff;
    decBuf[1660] = 256'h85ff81ff76ff67ff59ff4dff45ff40ff3fff3dff3fff40ff3fff3cff38ff32ff;
    decBuf[1661] = 256'h31ff2cff28ff25ff21ff17ff0eff00fff4fee8fedbfecffecdfecbfecafecbfe;
    decBuf[1662] = 256'hcffecefecbfec3feb7fea8fe96fe7cfe64fe54fe40fe38fe3afe3cfe42fe4ffe;
    decBuf[1663] = 256'h54fe58fe51fe41fe2efe16fe00feecfddffdddfde3fdedfdf2fdfafdfcfdf5fd;
    decBuf[1664] = 256'hecfddbfdc6fdb8fdb0fda9fdaffdb5fdbefdccfdcefdcdfdc5fdbafda8fd98fd;
    decBuf[1665] = 256'h89fd83fd88fd90fda1fdb4fdc1fdcdfdd7fdd1fdc2fdaefd97fd81fd73fd60fd;
    decBuf[1666] = 256'h59fd64fd6efd7dfd91fd9efda0fd9afd84fd6afd4afd24fd0afdf3fce7fce3fc;
    decBuf[1667] = 256'hedfcf7fc05fd12fd10fd05fdf7fcddfcc2fca2fc84fc71fc6efc64fc67fc6ffc;
    decBuf[1668] = 256'h71fc6ffc75fc70fc6bfc67fc5dfc54fc51fc4efc4bfc4cfc4dfc4efc50fc4afc;
    decBuf[1669] = 256'h46fc43fc3bfc34fc2ffc27fc21fc1efc1afc15fc18fc14fc0dfc0dfc03fcf9fb;
    decBuf[1670] = 256'hf3fbe9fbe2fbe6fbe7fbecfbf6fbfcfb03fc0bfc0afc03fc01fcf4fbeafbddfb;
    decBuf[1671] = 256'hcffbc5fbc3fbb8fbb0fbacfba6fba2fba5fba3fba2fba5fb9efb98fb92fb85fb;
    decBuf[1672] = 256'h77fb75fb6dfb69fb6afb70fb7dfb8ffb9afba5fbb3fbb1fbb0fba8fb99fb8bfb;
    decBuf[1673] = 256'h7ffb73fb6ffb70fb6ffb75fb80fb87fb94fba2fba4fba9fbb2fbb0fbaffbb0fb;
    decBuf[1674] = 256'hadfbaefbb2fbb5fbc0fbd2fbdefbf1fb03fc0ffc1afc1cfc1afc18fc14fc0afc;
    decBuf[1675] = 256'h01fcfefbf9fbf8fbfefb03fc0bfc1bfc27fc36fc48fc59fc63fc71fc7afc82fc;
    decBuf[1676] = 256'h8afc8bfc87fc8dfc90fc96fca3fcb1fcc1fcd8fceefcfdfc05fd02fd00fdf6fc;
    decBuf[1677] = 256'he3fccbfcbcfcadfca0fc9efca0fcaafcbdfcd5fcebfcfffc0cfd18fd1afd14fd;
    decBuf[1678] = 256'h04fdf5fce7fcdbfcddfce7fcf9fc1dfd40fd61fd87fda1fdaffdaafd9ffd8dfd;
    decBuf[1679] = 256'h77fd63fd5bfd59fd5ffd75fd95fdbbfddffd09fe25fe3efe56fe5afe56fe52fe;
    decBuf[1680] = 256'h49fe4cfe4ffe5afe72fe8efeb1fed1feeffe02ff0dff10ff07fffafeeefee4fe;
    decBuf[1681] = 256'hdafed8feddfeeafefafe09ff17ff23ff2fff39ff40ff4bff5cff6fff86ff96ff;
    decBuf[1682] = 256'haaffbdffc4ffc6ffc8ffc3ffbeffbcffbbffc1ffcbffd5ffdeffe5ffe8ffe8ff;
    decBuf[1683] = 256'he0ffd3ffc1ffb6ffabffa5ffa7ffafffc2ffdafff6ff19003000450059006300;
    decBuf[1684] = 256'h60005d005b0058005a006000700083009b00aa00b900c100c300c100b700b200;
    decBuf[1685] = 256'hb000b500c600dc00fb00190134015401690175017801750172017a017c017f01;
    decBuf[1686] = 256'h8d01a001b201c301cd01d301d201c301ad019901810165015a014f0152015b01;
    decBuf[1687] = 256'h72019501b501d301e601f801f501ec01df01ce01bf01bd01c601d501ef010e02;
    decBuf[1688] = 256'h2c023f024a0247023e022c0212020002ea01dc01d901d701d901e301ec01f401;
    decBuf[1689] = 256'hfb01fd01fe01ff01fe01fd01020208020a0216021b021f0221021d0215021202;
    decBuf[1690] = 256'h0802ff0100020602110224023c0252026b027602790270025e0249023a023202;
    decBuf[1691] = 256'h350248026a029402c602f60216033203370329031403f902d202c302b502b102;
    decBuf[1692] = 256'hc402dd02f9021c033c0349034d034903390325030803ed02dc02d202ca02d702;
    decBuf[1693] = 256'hec0206031f033b035603600364035b0353034c033d032f032a03250326032503;
    decBuf[1694] = 256'h21031e0319030f0308030003f802f702f402f002f102ee02e102d302c002a802;
    decBuf[1695] = 256'h98028a0282028e029d02b702d602f402080319031c0314030603ec02c602ac02;
    decBuf[1696] = 256'h950288028c029702b302d602ff0227034b0358035d03510332031403f102d102;
    decBuf[1697] = 256'hc402cf02e10203032d03540378038f039403800361033a030203dd02ac029a02;
    decBuf[1698] = 256'h8902840288029e02a902bb02c402cd02cf02c802b9029f028702710251024502;
    decBuf[1699] = 256'h3902350239024102540264026f02750277026e025e0247022a020f02f001db01;
    decBuf[1700] = 256'hcf01cb01c801d101e301f9010d022402340237023a0229021202f501da01c901;
    decBuf[1701] = 256'hb901b601b901c501d401e601f201f401ee01e501d301be01af01a2019b019d01;
    decBuf[1702] = 256'ha301ac01bb01c101c601ce01d201d101d201d101cc01cd01c901c301bc01b101;
    decBuf[1703] = 256'ha6019e0192018a0188018401850189018a0189018d0192019401970198019901;
    decBuf[1704] = 256'h990192018c0185017a017101670163015d0159015401500148013c012d012301;
    decBuf[1705] = 256'h10010301f700ec00e600dd00dc00d700d600d200cc00c900ca00cf00d100d400;
    decBuf[1706] = 256'hd300d600d500cf00c900c100b400a6009c008f008b0080007c007b007a007f00;
    decBuf[1707] = 256'h860091009d00ac00b600bb00b900af009d008700730061005a00600072008c00;
    decBuf[1708] = 256'hac00c100d400d800c800ae0088005a002200fcffdaffc7ffcdffe6ff07002400;
    decBuf[1709] = 256'h470068006c00600048001f00f8ffcaff9eff82ff7dff81ff96ffb2ffd8fffcff;
    decBuf[1710] = 256'h130017000c00ecffc6ff98ff6cff45ff2bff1dff19ff25ff36ff46ff54ff5cff;
    decBuf[1711] = 256'h63ff61ff5fff5aff52ff4aff40ff35ff2bff21ff16ff0eff0dff13ff22ff34ff;
    decBuf[1712] = 256'h49ff63ff75ff7eff7bff6eff54ff2dff09ffe9fecbfeb0feadfeb6fec4fedcfe;
    decBuf[1713] = 256'hf8fe1bff32ff47ff4bff41ff25fffafed3feaffe98fe8bfe87fe99feb5fed0fe;
    decBuf[1714] = 256'heffe05ff10ff0dfff7fed1fea3fe78fe50fe37fe29fe2dfe39fe51fe6dfe88fe;
    decBuf[1715] = 256'ha1feb7fec5fed2fed9fedbfed9fed4feccfec8febefeb5feb4feb7febafec5fe;
    decBuf[1716] = 256'hd0fedbfee2fee3fee0fed5febefea2fe87fe6efe52fe37fe26fe23fe25fe38fe;
    decBuf[1717] = 256'h52fe71fe8ffeaafec3feccfec9febcfea2fe7cfe62fe42fe35fe31fe3bfe51fe;
    decBuf[1718] = 256'h71fe8ffeaafeb4feb7fea9fe91fe75fe5afe50fe46fe4ffe67fe83fea6fecffe;
    decBuf[1719] = 256'hebfe05ff13ff17ff1bff10ff07fff9fef1feeafee3fee5fee4fee5fee4fee2fe;
    decBuf[1720] = 256'hdcfed6fecbfec4febdfeb7febafebffec5fed2fee4fef0fefbfe01fffffefefe;
    decBuf[1721] = 256'hfcfef5fef6fe01ff0dff1fff2fff3eff44ff46ff3eff30ff1dff0bfffffef4fe;
    decBuf[1722] = 256'heafee9fee7fee5feeafeedfeeefef3fefafefefe06ff0bff0eff13ff15ff13ff;
    decBuf[1723] = 256'h0dff08ff00fffbfef8fef7fefdfe08ff14ff21ff2eff2fff31ff32ff2cff26ff;
    decBuf[1724] = 256'h23ff1aff10ff07fffffe00ff03ff07ff14ff32ff50ff6bff84ff93ff9cff94ff;
    decBuf[1725] = 256'h84ff70ff5eff44ff39ff30ff33ff3bff50ff6aff83ff9fffaaffb5ffb8ffaaff;
    decBuf[1726] = 256'h97ff78ff5bff38ff21ff0bff07ff19ff3bff65ff98ffc8fff3ff10000a00fdff;
    decBuf[1727] = 256'hd6ffa8ff7cff55ff3bff40ff4dff68ff95ffc1ffddffedfffbffeeffdaffbbff;
    decBuf[1728] = 256'h95ff71ff50ff44ff38ff3cff45ff53ff6bff87ff9affacffc2ffcaffc8ffcaff;
    decBuf[1729] = 256'hbbffa5ff91ff7aff64ff55ff53ff55ff5bff6dff83ff9dffb5ffd1ffe5fff6ff;
    decBuf[1730] = 256'hf9fff1ffd9ffb7ff96ff79ff65ff62ff71ff9cffd5ff09004700700087008e00;
    decBuf[1731] = 256'h6e0047001900e1ffacff98ff91ffadffd1ff040034006d0083008a0084006800;
    decBuf[1732] = 256'h44002300fdffe3ffd6ffd1ffddffeeff04001e00370046004f004c0040002900;
    decBuf[1733] = 256'h1300f9ffe8ffdeffd6ffdeffeafff8ff06000f0017001c001d00210027002c00;
    decBuf[1734] = 256'h320038003a003a003200250017000900f9fff3fff1fff9ff08001a002f003e00;
    decBuf[1735] = 256'h40003e0038002a001a000f0009000b00100014001e00240028002f0035003700;
    decBuf[1736] = 256'h3a00390035002d001e0010000400f9fff4fff0fff4fffcff0700110018001e00;
    decBuf[1737] = 256'h240025002200230027002f0037003e00440047003f0030001e000900f5ffe8ff;
    decBuf[1738] = 256'he5ffe8fff6ff02001000160015000d00fcffe5ffcfffbbffaeffa6ffa4ffaaff;
    decBuf[1739] = 256'hb7ffc8ffdefff8ff0900190021001f000e00f7ffdbffb8ffa1ff8bff78ff7cff;
    decBuf[1740] = 256'h7fff93ffa5ffbbffc9ffd1ffcaffb7ff9fff89ff6fff5eff54ff51ff54ff5bff;
    decBuf[1741] = 256'h5dff63ff69ff71ff78ff82ff8dff98ff96ff90ff7fff60ff42ff20fffffeeafe;
    decBuf[1742] = 256'hdefee2fef1fe11ff2fff4aff62ff72ff7bff73ff62ff4bff35ff1bff0aff00ff;
    decBuf[1743] = 256'h03ff0bff25ff3eff60ff8affa6ffbfffcdffc9ffb6ff8fff61ff29ff03ffe1fe;
    decBuf[1744] = 256'hdbfeebfe05ff2fff61ff84ff96ffa7ff98ff8aff6cff49ff29ff14ff00fffdfe;
    decBuf[1745] = 256'h06ff1aff37ff5aff7bff98ffacffb6ffadff99ff77ff56ff30ff16fffffefbfe;
    decBuf[1746] = 256'hfffe09ff2cff43ff61ff6cff70ff6dff64ff57ff50ff4eff50ff5cff6aff78ff;
    decBuf[1747] = 256'h7eff7fff78ff76ff75ff74ff7dff88ff93ffa2ffacffb1ffacff9fff8fff7cff;
    decBuf[1748] = 256'h6aff59ff5bff61ff71ff88ffabffcbfff1ff0b0019002500290026001c001400;
    decBuf[1749] = 256'h0700fbfff9ffffff0e00260042005d006f007e0076006800530033001e001300;
    decBuf[1750] = 256'h0f00180032004b0067007a008c00950092009500970099009f00ac00b400bb00;
    decBuf[1751] = 256'hbf00bc00af00a100930083007d007b0087009500a300b000b800b600b200a700;
    decBuf[1752] = 256'h9900910089008d009400a200b100c000ce00db00e300e700eb00e500dd00d600;
    decBuf[1753] = 256'hcb00bc00b200b000b200ba00c300ce00dc00e100e000de00d700d100d200db00;
    decBuf[1754] = 256'he600fa00110121012a0132012a01240116010601000106011201240139014e01;
    decBuf[1755] = 256'h5b015d015201400126010701fa00ee00f200fb000a011c013101460148014b01;
    decBuf[1756] = 256'h4d0143013d0132012501180113010c010d0116011e012b013b0145014b014a01;
    decBuf[1757] = 256'h41013701280116010f0104010201070113011d01270130013301300126011d01;
    decBuf[1758] = 256'h160115011a012401300135013a013b0135012f012a01260128012b0131013b01;
    decBuf[1759] = 256'h4401480150015301500150014d01470142013b012e0126011f011a011e012201;
    decBuf[1760] = 256'h2d013d0150015d01690167015d014d0136011a010601fc00f900fc0009011e01;
    decBuf[1761] = 256'h380143014c014901410131012601180108010201fc00f700fb0003010a011801;
    decBuf[1762] = 256'h2b01380149014f0151014f014401330120010e01fd00f300f500fa0005011301;
    decBuf[1763] = 256'h1b0124012801210116010e010201f700f200e900e000da00d300cb00c800c500;
    decBuf[1764] = 256'hc400c700cd00d600db00d900d600cd00ba00a30093007f006c006a006c006e00;
    decBuf[1765] = 256'h7a00860093009c00a100a2009e009300860076006700550044003e0038003600;
    decBuf[1766] = 256'h42004f005f0069006f006e00660052003500220009000000fdff050016002d00;
    decBuf[1767] = 256'h3d004b00530050004600380028001d0013000e001300180019001d001e001d00;
    decBuf[1768] = 256'h13000a0003000000fbfffaff0000060012001d002200230022001c0013000800;
    decBuf[1769] = 256'hfafff2fff0ffeefff3fff9ff01000a000b000800fbffe7ffcaffafff97ff87ff;
    decBuf[1770] = 256'h84ff87ff9cffb6ffcfffe5fff3fff0ffe4ffd1ffbaffaaff96ff93ff96ffa5ff;
    decBuf[1771] = 256'hb3ffc6ffd3ffd5ffcfffbdffa8ff99ff82ff72ff6fff72ff79ff83ff8dff9aff;
    decBuf[1772] = 256'h9fffa0ff9fff9bff98ff95ff94ff93ff95ffa1ffa9ffb3ffc0ffc8ffc9ffc8ff;
    decBuf[1773] = 256'hbdffacff99ff91ff8aff84ff8aff96ffa5ffb7ffc3ffc9ffcbffc6ffbaffadff;
    decBuf[1774] = 256'ha1ff9fff9dffa4ffb2ffc5ffd2ffe3ffe9ffe7ffe6ffdaffcaffbbffb1ffa5ff;
    decBuf[1775] = 256'h9dff9bff97ff9bff9cff9dffa1ffa4ff9fff9dff98ff94ff8eff88ff85ff84ff;
    decBuf[1776] = 256'h83ff8aff91ff99ffa0ffa6ffa9ffa6ffa0ff98ff93ff90ff8bff8bff91ff99ff;
    decBuf[1777] = 256'ha0ffa5ffa6ffa2ff9cff96ff8aff7fff77ff79ff7dff84ff8fff9dffa9ffb5ff;
    decBuf[1778] = 256'hb9ffbdffb9ffb4ffadffa3ff9aff93ff94ff97ffa1ffb0ffbeffcaffd6ffdaff;
    decBuf[1779] = 256'hd6ffcdffbdffa7ff99ff8cff85ff87ff91ff9dffafffc4ffd3ffe0ffe2ffdcff;
    decBuf[1780] = 256'hd6ffcdffc2ffbaffb9ffbcffc4ffcdffd6ffdeffe1ffdeffdcffd6ffcfffc9ff;
    decBuf[1781] = 256'hc5ffc1ffc1ffc2ffc3ffc4ffc7ffc6ffc1ffc1ffbaffb8ffbaffc1ffc8ffd7ff;
    decBuf[1782] = 256'he5fff5ff04000e000c000400f6ffe3ffcbffbcffadffa6ffa8ffb3ffc5ffdaff;
    decBuf[1783] = 256'he8fff5fff8fff1ffdfffcaffb6ffa4ff93ff91ff9bffb2ffc7ffe7ff05001800;
    decBuf[1784] = 256'h23002c0023001100fcffe2ffd0ffc1ffb8ffbbffc2ffd1ffe3fff3fffeff0400;
    decBuf[1785] = 256'h0600fefff6ffe7ffd9ffd0ffcbffc7ffceffd9ffe3fff0fffeff000002000100;
    decBuf[1786] = 256'hfcfff0ffe8ffddffd1ffc5ffbeffbaffb6ffb3ffb2ffafffacffabffaeffafff;
    decBuf[1787] = 256'hb0ffadffacffabffa5ff9fff9bff96ff94ff8fff8dff8aff89ff85ff81ff7eff;
    decBuf[1788] = 256'h76ff6cff62ff5aff4fff49ff40ff3cff3bff39ff34ff37ff38ff34ff2fff2dff;
    decBuf[1789] = 256'h2cff2bff2cff2dff31ff32ff36ff3bff3bff39ff36ff30ff28ff20ff17ff11ff;
    decBuf[1790] = 256'h0eff0dff0fff15ff1aff1eff23ff1eff1aff17ff0eff04fffefef8fef5fef6fe;
    decBuf[1791] = 256'hf9fefbfefafefdfefefefbfef5feedfee8fee1fed9fed3fed2fecffec9fec5fe;
    decBuf[1792] = 256'hc2fec0febbfeb9febbfebafebbfebefec2fec3fec2fec1fec1febcfeb3feacfe;
    decBuf[1793] = 256'ha8fea2fe9ffea2fea6feaefeb8febcfec0fec1febcfeb4feadfea4fe9dfe98fe;
    decBuf[1794] = 256'h93fe92fe96fe9bfea2feaafeb3febcfec2febffebefebbfeb7feb1feacfea6fe;
    decBuf[1795] = 256'ha7feaafeabfeb1febafec4fecffed7fedefee4fee7fee4fee0fedafed4fecdfe;
    decBuf[1796] = 256'hc7fec5fecbfed8fee6fef2fe04ff15ff1fff21ff1cff17ff10ff06fffbfef6fe;
    decBuf[1797] = 256'hf5fefbfe08ff13ff1dff2dff33ff34ff33ff28ff1cff10ff06ff02ff03ff0bff;
    decBuf[1798] = 256'h18ff28ff37ff45ff4dff4fff4dff49ff41ff3bff3aff39ff43ff52ff60ff6cff;
    decBuf[1799] = 256'h77ff7cff7dff77ff6dff61ff55ff4eff4fff55ff5fff71ff82ff95ffa2ffa9ff;
    decBuf[1800] = 256'habffa9ffa1ff99ff97ff96ff99ffa4ffb0ffc2ffd7ffe6ffedfff5fff7fff1ff;
    decBuf[1801] = 256'hebffe3ffd9ffd7ffd9ffdaffe1ffecfff8ff02000c00120015001c0021002700;
    decBuf[1802] = 256'h2d003700430048004f0056005500520051004e00480049004d00510059006300;
    decBuf[1803] = 256'h700078007900750072006a005d0054004c004a005400640077009400af00c100;
    decBuf[1804] = 256'hd000d900d600cf00bc00af009e00940092009400a200b400ca00de00f000fc00;
    decBuf[1805] = 256'hfe00f800f300e700d700cc00c600c800d000e100f4000b0121013b0146014f01;
    decBuf[1806] = 256'h52014a01430138012e0122012001220126012f01400150015f0171017d018301;
    decBuf[1807] = 256'h850180017f0177016d016c017001750182019401a401b701ca01d101d701d901;
    decBuf[1808] = 256'hd101c801c101b701b101b001b101bb01c401cf01e001eb01ed01f201ed01e801;
    decBuf[1809] = 256'he401e101db01de01e201e801f60104020c02140219021a02190213020e020c02;
    decBuf[1810] = 256'h09020c02120216021c0228022d022e02320231022b022a022802220224022902;
    decBuf[1811] = 256'h2a023002360238023f0243024002450246024102440245024402460247024602;
    decBuf[1812] = 256'h4b024d024b024f025202510259025c025b026002640260025f025c0252025402;
    decBuf[1813] = 256'h53024d02520255025702610268026b02730274026e026f026c0261025c025802;
    decBuf[1814] = 256'h54025202530254025c026002630269026a02690266025e0254024d0242023802;
    decBuf[1815] = 256'h33022d0228022b02310237023f02440247024c0247023e02340221020f02fe01;
    decBuf[1816] = 256'hf401ea01eb01f001f8010c021b0223022a02280216020502f201da01c401b601;
    decBuf[1817] = 256'hae01b501c001ce01e501f401fd010502f901ea01d801be01a501900187017f01;
    decBuf[1818] = 256'h8b019601a801b801c301c101c301ba01a4018e017a0168015c01550153015901;
    decBuf[1819] = 256'h5d0165016c016d0165015c014c013d012f012301170113011201130116011701;
    decBuf[1820] = 256'h1801190115010d010501fc00f300ed00e600e200df00d900d300cb00bf00b400;
    decBuf[1821] = 256'ha9009a008c0083007b0074006f006c0066005f00570052004b00430036002e00;
    decBuf[1822] = 256'h2a0023001f00190016000f000200f7ffecffddffcbffbfffb0ffa6ffa5ffa3ff;
    decBuf[1823] = 256'h9fff98ff91ff8cff83ff75ff6cff5eff54ff4eff50ff55ff59ff5fff65ff6aff;
    decBuf[1824] = 256'h69ff63ff57ff49ff37ff26ff1bff0dff05ff00ff01ff05ff04ff05ff00fffafe;
    decBuf[1825] = 256'hf0fee4fed5fecbfebffeb7feb3feb4feb3feb6febdfebefebbfebefebbfeb3fe;
    decBuf[1826] = 256'ha9fe9dfe92fe87fe78fe6afe5efe52fe45fe39fe30fe2cfe28fe24fe23fe24fe;
    decBuf[1827] = 256'h20fe1bfe15fe0dfe05fefcfdf1fde7fde0fddefde0fde3fde9fdebfdf0fdf1fd;
    decBuf[1828] = 256'hecfde6fddbfdc9fdbdfdaefda0fd97fd92fd91fd98fd9efda4fdadfdb0fdb2fd;
    decBuf[1829] = 256'hb3fdacfda6fda0fd9afd96fd95fd90fd91fd97fd9afd9dfda3fda0fda3fda5fd;
    decBuf[1830] = 256'ha3fd99fd95fd8cfd82fd7efd73fd6bfd6afd66fd65fd6afd69fd6efd75fd79fd;
    decBuf[1831] = 256'h7afd79fd73fd6dfd67fd5ffd59fd56fd57fd5bfd65fd6cfd75fd7cfd7dfd7bfd;
    decBuf[1832] = 256'h78fd70fd64fd59fd51fd4dfd4efd4dfd50fd5bfd60fd5ffd63fd5ffd57fd4efd;
    decBuf[1833] = 256'h48fd3efd3dfd39fd3efd47fd4bfd53fd5afd57fd55fd50fd47fd3dfd34fd2dfd;
    decBuf[1834] = 256'h2cfd2efd2ffd33fd3afd3afd3bfd3afd33fd2bfd26fd20fd19fd19fd1bfd21fd;
    decBuf[1835] = 256'h2bfd35fd40fd47fd4bfd4ffd4efd4bfd4cfd4dfd48fd49fd4efd4ffd51fd52fd;
    decBuf[1836] = 256'h4ffd52fd55fd52fd51fd54fd4ffd4ffd53fd50fd4ffd50fd4efd4ffd4ffd4ffd;
    decBuf[1837] = 256'h53fd5dfd63fd6cfd76fd7afd81fd82fd7bfd75fd70fd65fd5dfd5bfd57fd5bfd;
    decBuf[1838] = 256'h63fd68fd71fd78fd77fd78fd75fd68fd5efd59fd51fd52fd56fd5dfd69fd78fd;
    decBuf[1839] = 256'h86fd8efd93fd92fd8bfd85fd7afd71fd6dfd6efd73fd7ffd8afd94fd9efda7fd;
    decBuf[1840] = 256'ha8fda7fda1fd97fd93fd8dfd8cfd93fd9cfdabfdbdfdc9fdd4fddafdd8fdd0fd;
    decBuf[1841] = 256'hc9fdbffdb9fdbafdbbfdc1fdcefddcfdecfdfbfd01fe02fe01fef9fdf0fde9fd;
    decBuf[1842] = 256'he4fde3fde9fdf1fd02fe12fe21fe27fe30fe2bfe27fe20fe17fe0ffe10fe11fe;
    decBuf[1843] = 256'h1bfe27fe36fe48fe53fe5afe60fe65fe63fe5ffe5bfe5cfe64fe6dfe78fe89fe;
    decBuf[1844] = 256'h93fe9dfea6fea8fea3fe9afe91fe89fe88fe8bfe8ffe97fea5feaffeb8fec4fe;
    decBuf[1845] = 256'hc8fec4fec0febbfeb6feb3feb4feb8fec5fed7fee8fef7fe05ff07ff05fffdfe;
    decBuf[1846] = 256'heefee0fed8feccfecbfeccfed5fee3fef5fe01ff10ff16ff18ff1aff15ff0eff;
    decBuf[1847] = 256'h0aff09ff10ff1dff2bff42ff58ff66ff79ff85ff87ff85ff80ff7bff70ff6cff;
    decBuf[1848] = 256'h6dff73ff78ff83ff8fff9cffa5ffadffb2ffb3ffafffaeffabffaeffb7ffc1ff;
    decBuf[1849] = 256'hccffdaffe9fff8fffeff040002000000fafff1ffebffe6ffe9ffeafff0fff6ff;
    decBuf[1850] = 256'hfafffdfffefff8fff0ffe8ffe1ffdbffdaffe2ffeefffdff0b001e0030003800;
    decBuf[1851] = 256'h420040003b0033002b00240026002b0034004200520065007200790077006d00;
    decBuf[1852] = 256'h640056004c00430045004c005e0073008d00a600bc00ca00cd00ca00c000b600;
    decBuf[1853] = 256'had00a500a600b000c000d700ed0001010f01160114010a01fa00eb00e100d800;
    decBuf[1854] = 256'hd700e400f40007011f01340143014b014d014701410134013001340138014801;
    decBuf[1855] = 256'h600176019001a101b101b901b701ab01a4019a01920193019b01a701bc01d001;
    decBuf[1856] = 256'he301f301fe0100020202fa01ef01eb01ef01f401010215022c0242025c026702;
    decBuf[1857] = 256'h76027902760274026e02640265026a026f027e0290029c02ab02b502b602bb02;
    decBuf[1858] = 256'hba02b602b702ba02b902c302d202e002f3020603160329033c03480352035c03;
    decBuf[1859] = 256'h62036d037703810391039c03a203ae03bd03c303cc03d403db03e503ee03f303;
    decBuf[1860] = 256'hfe0309040a0415042304280437044904550463047504810494049c04a304ae04;
    decBuf[1861] = 256'hb004ae04b304b504b604bc04c004c304d004d604d404d904dd04dc04dd04e104;
    decBuf[1862] = 256'he004eb04fa0404051a0530053f0556056c0575057d0589058b05910599059b05;
    decBuf[1863] = 256'ha905b805c305d505e605ec05fa05030601060606040603060b0616061d062f06;
    decBuf[1864] = 256'h4506530670068306870696069f069c06a306a606a006a806b406b806c706d106;
    decBuf[1865] = 256'hd706e206e606e006e306de06d106d206d406d006df06ed06f206070715071807;
    decBuf[1866] = 256'h240726072007220723071f07290734073b074d075e0764077207770773077107;
    decBuf[1867] = 256'h6a075a075c075a0758076a077b078a07a007ae07b107b807b1079f0798078e07;
    decBuf[1868] = 256'h7c077907800782079507a207a907b807c207af07a20791077507620751074107;
    decBuf[1869] = 256'h4a07510754076707790777077d0777076107510737071f070f070607fe060a07;
    decBuf[1870] = 256'h19071f0732073a072e072c0722070c07fc06f306e106e306ea06ec06fb060607;
    decBuf[1871] = 256'h0c0711070c07fc06f106df06c506bb06b106a906ab06ae06ac06b206a9069406;
    decBuf[1872] = 256'h85066e0652063e062d061d062006230620062b062906200618060406e205cb05;
    decBuf[1873] = 256'ha505810573056605630566056f056d056f055f0547052b050005d904b5049504;
    decBuf[1874] = 256'h880484048f049804ac04bf04c104bf04ad04890465043c041404fb03e403df03;
    decBuf[1875] = 256'heb03fc030c04150417040204e803c2038903550325030503f402ef02f4020903;
    decBuf[1876] = 256'h1d0327032a031c03fa02d0029d026d02350210020902020208020d021b021f02;
    decBuf[1877] = 256'h1402fb01d901a60176013e010901e700d400ce00d300d800e500e900de00cf00;
    decBuf[1878] = 256'haf0089005b002f001300f9ffe2ffdeffe2ffdeffdbffd8ffcbffb6ff96ff70ff;
    decBuf[1879] = 256'h42ff22fffbfed7fec9feb4fea8fe9efe8efe80fe68fe46fe1cfef5fdd1fdb1fd;
    decBuf[1880] = 256'h93fd78fd5ffd56fd42fd2ffd1ffd03fde0fcc0fc91fc65fc49fc30fc0ffc02fc;
    decBuf[1881] = 256'heffbe5fbd5fbc1fba4fb89fb5bfb30fb08fbe4fabbfaaafa90fa8cfa87fa7cfa;
    decBuf[1882] = 256'h71fa6efa54fa35fa17faecf9c5f9a1f98af975f969f95ff95bf95ef951f941f9;
    decBuf[1883] = 256'h2df906f9dff8b1f885f852f830f811f8f4f7eff7e1f7ccf7c8f7b0f794f780f7;
    decBuf[1884] = 256'h53f727f70bf7e7f6c7f6baf69ff68df684f676f668f65df63df61cf607f6e4f5;
    decBuf[1885] = 256'hbbf59ef57bf55af545f522f50bf5fef4dbf4c4f4b7f4a4f48cf488f474f467f4;
    decBuf[1886] = 256'h65f452f43ff438f41df409f4fff3e3f3cff3d3f3bdf3b4f3b2f3a1f38ef381f3;
    decBuf[1887] = 256'h5df339f322f3f3f2c8f2b7f29df28ff293f288f28bf2a1f293f286f283f263f2;
    decBuf[1888] = 256'h43f236f20cf2f0f1eaf1ddf1d8f1ecf1e8f1ebf1f4f1e2f1c3f1b6f17cf153f1;
    decBuf[1889] = 256'h3cf10cf1f9f0f4f0eef0fcf01af11ef121f137f123f111f105f1e5f0c5f0c0f0;
    decBuf[1890] = 256'ha5f0a2f0bef0c2f0d3f0f6f0f1f0edf0f1f0caf0a6f098f06af04af045f02bf0;
    decBuf[1891] = 256'h30f045f051f062f078f075f06df070f050f02ff02bf010f006f015f012f01ff0;
    decBuf[1892] = 256'h3ef043f04ef060f04af036f02ef00ff0faeff6efe4efe1effbefffef14f034f0;
    decBuf[1893] = 256'h30f034f045f036f027f02ff023f025f03bf044f056f07af089f097f0acf0a9f0;
    decBuf[1894] = 256'ha5f0a8f09af097f0a8f0a6f0b4f0cef0e9f0fbf01df122f126f131f120f11df1;
    decBuf[1895] = 256'h25f11ef129f149f157f16cf197f1a8f1b7f1cef1caf1c6f1d1f1c1f1c4f1dcf1;
    decBuf[1896] = 256'hdff1f9f11ff239f259f27ff285f292f2a8f29cf2a0f2aff2a7f2b4f2cef2e6f2;
    decBuf[1897] = 256'h02f32df349f363f38cf392f3a1f3aff3b4f3b7f3d0f3d9f3f9f31ff443f463f4;
    decBuf[1898] = 256'h92f4b1f4cef4f1f4fff40cf527f52bf534f54ef55ff57cf5a6f5c2f5e6f510f6;
    decBuf[1899] = 256'h2cf646f666f673f686f69ff6a8f6c2f6e1f6f7f619f74cf76ff79af7c2f7e6f7;
    decBuf[1900] = 256'h06f82cf83cf853f871f884f89cf8bff8d6f8fcf82af93df964f993f9b2f9d9f9;
    decBuf[1901] = 256'hfdf914fa3afa5efa75fa9cfac0fae0fa0ffb3afb57fb85fbb0fbcdfbfbfb26fc;
    decBuf[1902] = 256'h43fc66fc90fcacfcd0fcf0fc0efd29fd49fd67fd91fdb9fddcfd06fe2dfe5cfe;
    decBuf[1903] = 256'h87feaffed3fef3fe11ff2cff4bff69ff8cffacffdbff070039006a009500bd00;
    decBuf[1904] = 256'heb000a0126014001570175018801af01dd0108023b026b02a302d80208033403;
    decBuf[1905] = 256'h500374038b03a903c403dc03ff03320454048c04d004fd0437055d058d05ac05;
    decBuf[1906] = 256'hc805d705f8050d06200647067506a106df0629075b078907c207d907fb071a08;
    decBuf[1907] = 256'h15082e083c08520874089e08d1080f0948097d09ad09d909ea09030a110a0d0a;
    decBuf[1908] = 256'h200a400a550a870ac50aee0a320b720b9b0bd00be40bea0bf00bf50bf10b0e0c;
    decBuf[1909] = 256'h290c420c710cbc0cee0c2e0d580d6e0d900da30d9e0dad0dbb0dbf0dea0d110e;
    decBuf[1910] = 256'h3f0e840ec40eed0e220f440f4a0f5b0f560f480f5d0f690f730f9c0fcf0ff10f;
    decBuf[1911] = 256'h29105e1080109f10bc10ac10ba10be10b310cb10e710fb102f1164118611be11;
    decBuf[1912] = 256'he411f8110b121c120d121112161202121b1231123f1266129912ae12d912f512;
    decBuf[1913] = 256'hfb1208130d13f212fc12f912f0120d1328133a1369139913ac13d313ed13df13;
    decBuf[1914] = 256'he313d713b813b413b0139e13c113d813ed1318143f1444145b1457143c143114;
    decBuf[1915] = 256'h1514f213f713fb13f7131e14421450147e1491148014901478144a1437142614;
    decBuf[1916] = 256'h021407141414171437144c145014621465143f143a141a14eb13e513d413c513;
    decBuf[1917] = 256'hd213df13db13fb130814f413f813e813c313b3139c1376137b136d1360137413;
    decBuf[1918] = 256'h7013611369135c133d1331131d13f012e912d912b512b912ad1291129c128c12;
    decBuf[1919] = 256'h6d12681255122f121f121112eb11e611d811ba11b611a51183117e1169113e11;
    decBuf[1920] = 256'h2d111e11f410ef10df10b610b010a110771071104d102d1020100510df0fda0f;
    decBuf[1921] = 256'hcc0fae0faa0f990f700f6a0f460f1d0f0c0ff20ec90ec30eb40e930e8f0e830e;
    decBuf[1922] = 256'h640e570e340e010edf0dc00d820d690d530d300d370d260d160d1b0d060de30c;
    decBuf[1923] = 256'hc20c9c0c640c3e0c0e0cd60bce0bba0ba70bad0bb20ba40b970b7c0b480b130b;
    decBuf[1924] = 256'hd50a8b0a590a2b0af209ea09e309e909fa09f509e709d209a7096a091f09d908;
    decBuf[1925] = 256'h990860083a0826082c08310837084e0841082608f807b40761071407ba067e06;
    decBuf[1926] = 256'h5d063f0636063e0645064c06530636060806d0058d052805e504a90472045404;
    decBuf[1927] = 256'h5d0455046b0472046c045b042d04e803a8035e030403c70290025e0255024d02;
    decBuf[1928] = 256'h54025b026102510237020402c6017c013601e400ad008f006100590060006700;
    decBuf[1929] = 256'h6e0068004e002e00f7ffb3ff61ff14ffcefea0fe77fe61fe68fe6efe73fe79fe;
    decBuf[1930] = 256'h6bfe4dfe1bfeddfd92fd38fdfcfcaffc7dfc61fc59fc61fc68fc7afc75fc65fc;
    decBuf[1931] = 256'h3cfcfefbb4fb6efb1bfbcefa9cfa81fa79fa80fa87fa8dfa9efa85fa64fa2dfa;
    decBuf[1932] = 256'hdbf98ef948f9f5f8bef8a0f897f88ff8a6f8acf8b3f8adf87ff853f815f8cbf7;
    decBuf[1933] = 256'h85f757f71ef7f8f6f1f6ebf6f1f6f6f6f1f6dcf6c1f693f64ff621f6d7f5a5f5;
    decBuf[1934] = 256'h77f54ef537f530f52af519f514f5fdf4d7f4bdf48af45af43bf408f4d8f3d2f3;
    decBuf[1935] = 256'habf39bf397f379f35ef34cf31df3edf2cef29bf279f25af232f20ef201f2e3f1;
    decBuf[1936] = 256'hc8f1b6f18ef166f157f124f102f1eff0bcf0a8f0a1f085f076f071f053f038f0;
    decBuf[1937] = 256'h20f0f1efc1efa2ef6fef3fef2cef10eff6eefbeeddeed2eed5eeb3ee92ee7dee;
    decBuf[1938] = 256'h4bee1beefbedc9eda6edaded90ed96edadeda0ed9ceda0ed7ded5ded3fed05ed;
    decBuf[1939] = 256'hcbecb5ec85ec72ec83ec73ec78ec9eec8fec8aec8eec64ec3cec23ece7ebbdeb;
    decBuf[1940] = 256'hb6eba1eb9bebb7ebb2ebc0ebd5ebcaebb8ebb5eb8aeb6beb5aeb36eb1feb23eb;
    decBuf[1941] = 256'h17eb1beb37eb33eb37eb46eb2ceb1beb1eebfeeaf2eafdeaeceae9ea02ebf1ea;
    decBuf[1942] = 256'heeea02ebeaeadbeae3eac6eabbeacceac3eacceaf3eaf9eafeea1eeb11eb06eb;
    decBuf[1943] = 256'h09ebe7ead9eaddead2eae3ea0ceb1deb36eb69eb70eb76eb87eb63eb43eb3feb;
    decBuf[1944] = 256'h0cebf8ea0aeb10eb34eb79eb97ebd7eb11ec18ec1fec32ec0becf1ebe3ebc5eb;
    decBuf[1945] = 256'hc9ebe9ebfeeb30ec7cecaeecc9ec03edfcecf5eceeecbcec99ec93ec82ec87ec;
    decBuf[1946] = 256'hbaecddec15ed67ed88edbaede8edf0edf8edf1edd2edcceddbedd7edeced1eee;
    decBuf[1947] = 256'h41ee79eeaeeed0eee3eeffeeefeeebeef8eedceed9eeefeef7ee0fef3eef60ef;
    decBuf[1948] = 256'h80efbdefd6effcef2cf032f04ef072f077f094f0b7f0c5f0d2f0f5f0f9f00ff1;
    decBuf[1949] = 256'h32f136f154f17ff19bf1bff1e8f1f9f11df234f238f24cf264f267f27bf2a3f2;
    decBuf[1950] = 256'hcaf203f346f386f3c0f303f41ff448f45ef457f451f462f45df474f49af4bef4;
    decBuf[1951] = 256'hfaf445f577f5a4f5def503f618f62bf630f636f64df662f68df6caf604f748f7;
    decBuf[1952] = 256'h9af7d1f703f830f849f860f874f87bf88bf8a5f8c5f8f4f82cf952f990f9caf9;
    decBuf[1953] = 256'heff911fa31fa42fa65fa7dfaa3fad1fa09fb3efb89fbbbfbfbfb24fc3bfc50fc;
    decBuf[1954] = 256'h62fc73fc83fca3fcd2fcfdfc47fd8dfdccfd17fe49fe64fe6cfe74fe6dfe67fe;
    decBuf[1955] = 256'h78fe91fec4fe10ff6affd7ff3e008100be00df00e900cd00b4008f007a008100;
    decBuf[1956] = 256'ha800f5005801d0016202c5021e032e033d031503d802a10283027a029302e502;
    decBuf[1957] = 256'h5e03f103a10418058405bf05ad057c053305d50480045f04690497040205a405;
    decBuf[1958] = 256'h3c06ec066307a407df07a90758070e07b006740669068706eb067e072f08d508;
    decBuf[1959] = 256'h6d09cf09e109d00987090e09bd08560813081f086c08da087c093f0ac10a380b;
    decBuf[1960] = 256'h790b8d0b7b0b2a0bc20a650a400a1f0a510ab60a2e0be10b870cc80c2a0d3c0d;
    decBuf[1961] = 256'h2c0de20c9f0c320ce80bdb0bcf0b1c0c8a0cf10c840d0d0e430e940ea30e600e;
    decBuf[1962] = 256'h3c0e050ed30db70dc00de50d310e9f0ee90e610f920fbe0fe60fc20f8b0f6d0f;
    decBuf[1963] = 256'h3f0f260f2e0f420f6e0fc30f17104e109410c210ca10d210cb10ac10a610a110;
    decBuf[1964] = 256'h9c10c310e61007113e11641178119711921182117e1171115e116f117f118d11;
    decBuf[1965] = 256'hb511e711ee111a122b121b1220121312f81103120612fd112412411250127012;
    decBuf[1966] = 256'h86128212851276124a12441228120e12261232123e1272129812ad12cc12dd12;
    decBuf[1967] = 256'hcd12c912b312891278125e1247125412601263128c12a812ad12c412c0129d12;
    decBuf[1968] = 256'h98127b12481234122d121c122c12431258128b12ad12c012dc12e112c112b412;
    decBuf[1969] = 256'h91125e123c122912021207121512101233124112451259125512331225120712;
    decBuf[1970] = 256'hd511ce11bb11aa11c411e411f111231246124c125d1258122e121212ee11a911;
    decBuf[1971] = 256'h8b116f1146113f1146113f115b11751170117d11721152113d111a11f010df10;
    decBuf[1972] = 256'hd010b910ce10e210f3101c1138113d11421135110211e0109b105b102210fc0f;
    decBuf[1973] = 256'hcc0fd20fd80fd30ff30f081005100f10ff0fd40fb50f8e0f4b0f300f170f000f;
    decBuf[1974] = 256'h150f280f390f670f7a0f740f6f0f4e0f0f0fcf0e850e2b0e060ecf0d9d0da60d;
    decBuf[1975] = 256'hbf0dc70de90dfc0df60dfb0dd20d940d5a0d160dd70c9d0c860c720c840ca10c;
    decBuf[1976] = 256'hba0cdb0cf00cdc0cc40c950c2e0ce40b870b190bed0ac50aa10ac20ae00afb0a;
    decBuf[1977] = 256'h140b2a0b080be90aa00a460af1098e094b09260905090f093d0966097d099f09;
    decBuf[1978] = 256'h990966092809ce086108f9079c075f073e0734074f0779078f07a407b7079a07;
    decBuf[1979] = 256'h62071007ad064f06fa05ad058f0586058e05a505d505e805e205d305a9056005;
    decBuf[1980] = 256'h1a05b50458041b04fa03dc03e503ee03f5030a041004ff03db03a8035d031703;
    decBuf[1981] = 256'hd7028d025b023f0226021f0218021e0219020902e901c30195015c012801f800;
    decBuf[1982] = 256'hbf009a00780065005f00500039002c000900e9ffbaff8eff5cff1efff4fec0fe;
    decBuf[1983] = 256'h90fe64fe48fe24fe04feeefdd3fdb4fd96fd73fd4afd22fdfefcd5fcb9fc95fc;
    decBuf[1984] = 256'h6bfc4ffc2bfc0bfcedfbc2fb9bfb77fb44fb14fbe8fab6fa86fa5afa32fa04fa;
    decBuf[1985] = 256'he5f9bef99af979f94bf91ff903f9dff8b5f899f880f85ff84af827f807f8e9f7;
    decBuf[1986] = 256'hc6f79cf775f73df708f7e6f6aef679f664f639f611f602f6e2f5c4f5b0f58af5;
    decBuf[1987] = 256'h66f54ff520f5f4f4cdf49ff480f46ff44bf43df439f425f41bf412f4f2f3ccf3;
    decBuf[1988] = 256'hb2f376f33cf317f3d9f29ff289f274f261f267f262f266f273f258f23ff22af2;
    decBuf[1989] = 256'hfef1baf18cf163f12ef127f115f11af134f139f13df150f13ff11cf105f1c5f0;
    decBuf[1990] = 256'h86f04cf017f0f5efefefe9efeeef18f034f043f064f057f03cf02af0fbefb0ef;
    decBuf[1991] = 256'h92ef52ef39ef41ef3aef4def74ef83ef9aefb8efa5ef85ef70ef36ef0defe7ee;
    decBuf[1992] = 256'hc5eea6eeb6eebceedcee0bef1def3aef5def50ef43ef2feffbeec6eeb2ee86ee;
    decBuf[1993] = 256'h75ee85ee80ee95eeb8eec6eedbeef6eee5eed5eecdeea5ee89ee7aee63ee5eee;
    decBuf[1994] = 256'h79ee7dee93eebeeed1eee2eefbeee4eee0eedceebceea7eea3ee8bee88ee96ee;
    decBuf[1995] = 256'h93ee9beeb6eeb2eebdeed3eecaeecdeeddeed7eeddeef4eef7eeffee17ef14ef;
    decBuf[1996] = 256'h1def2fef28ef2eef44ef47ef54ef78ef7def94efa9efa5efa9efb9efa4ef9def;
    decBuf[1997] = 256'h9fef94ef9eefb9efcceff2ef2bf050f073f09ef0a4f0b3f0c1f0acf0a0f0abf0;
    decBuf[1998] = 256'ha2f0b0f0d2f0e9f018f150f176f1a6f1c5f1d6f1d1f1d5f1c0f1adf1b7f1a8f1;
    decBuf[1999] = 256'hb0f1d8f1fff12df27ef2b5f2e7f215f32ef335f34af32bf31af31ff311f31ef3;
    decBuf[2000] = 256'h41f361f398f3dcf31cf455f48af491f4a4f4a9f485f477f46bf457f462f484f4;
    decBuf[2001] = 256'haef4e0f42cf572f5b2f5ecf502f609f60ff6fef5eff5eaf5def5e2f50ff62ef6;
    decBuf[2002] = 256'h6cf6b6f6e8f628f762f779f77ff786f775f765f758f753f75ff77ef7a5f7ddf7;
    decBuf[2003] = 256'h21f84ef888f8cbf8d5f8edf804f9fdf8f7f8fcf8f7f805f92bf94ff982f9c0f9;
    decBuf[2004] = 256'he9f91efa4efa6dfa7efa8dfa7ffa84fa88fa84fa94fab3fad1fafcfa2efb5efb;
    decBuf[2005] = 256'h8afbb2fbd5fbedfb02fc06fc10fc20fc34fc4cfc6efc8efcbdfce9fc05fd29fd;
    decBuf[2006] = 256'h49fd5efd72fd83fd93fda7fdbffdd5fdfafd14fe34fe5afe74fe8bfea0febbfe;
    decBuf[2007] = 256'hcdfee9fe04ff2bff4eff78ff9fffceffedff0900230030003d00490053006900;
    decBuf[2008] = 256'h8900a700d9000901350167018a01a901ba01c901ce01d201d601e101f6011c02;
    decBuf[2009] = 256'h4a028202b702f5021e03430366036c0372036c0371036d0371038903ac03d503;
    decBuf[2010] = 256'h080446047f04b404d604e904fa04ff04f104e404e104dd04ed040c0533056b05;
    decBuf[2011] = 256'h9f05dd0507062c06410647064d063d062f0623061f06300653067306aa06df06;
    decBuf[2012] = 256'h0f0747076d0773077a0774075a07560749073d074f0765077f07ac07e4070a08;
    decBuf[2013] = 256'h2c084c085c08620866085908560852084f085d087a089508bc08ea0809093109;
    decBuf[2014] = 256'h4a094f095c095f095509520955094d095909680976099009ba09cb09ef09060a;
    decBuf[2015] = 256'h130a260a310a2e0a3c0a440a4b0a5a0a700a790a960ab10abb0ad70aeb0aee0a;
    decBuf[2016] = 256'h040b0d0b0f0b200b2b0b310b400b4f0b510b610b6c0b6e0b810b8e0b950bb10b;
    decBuf[2017] = 256'hcc0bdd0bf90b1c0c210c3f0c4a0c470c500c4d0c3b0c420c4d0c4f0c690c8c0c;
    decBuf[2018] = 256'h9a0cc80ce80ced0c070d0c0df60cf20ce80cd20cdb0ce80cef0c0f0d420d640d;
    decBuf[2019] = 256'h9c0dc20dc90dcf0dd50dbb0dad0d980d840d880d910d9a0dc10de90d020e2c0e;
    decBuf[2020] = 256'h480e4d0e5b0e570e430e400e300e220e2a0e3a0e410e5f0e850e940ebe0ecf0e;
    decBuf[2021] = 256'hd40ee20ede0ed20ecf0ec50eb10eb90ebb0eb50ecb0ed90ee10efb0e140f170f;
    decBuf[2022] = 256'h2b0f380f2c0f3b0f390f260f2e0f270f180f1e0f230f1b0f310f3b0f3e0f550f;
    decBuf[2023] = 256'h5f0f560f630f610f490f460f380f200f1d0f1a0f0d0f1e0f2d0f2f0f490f640f;
    decBuf[2024] = 256'h680f770f7a0f680f650f560f380f230f180ff80efc0e000ffd0e190f2c0f300f;
    decBuf[2025] = 256'h460f4e0f410f3f0f2c0f040ff30eda0eb90ebe0ec10ebe0ee00ef70e040f270f;
    decBuf[2026] = 256'h350f280f1d0f040fd50eb30e940e6c0e5d0e580e5c0e780e900ea60ec60ed20e;
    decBuf[2027] = 256'hc70ec30ea70e750e600e340e0d0e080e030eff0d1a0e330e3c0e560e590e4a0e;
    decBuf[2028] = 256'h3b0e190ee60dc40d980d660d510d4b0d450d540d620d670d820d850d6f0d670d;
    decBuf[2029] = 256'h4a0d1f0d030dd50ca90c980c890c720c760c7a0c6f0c730c700c580c4f0c350c;
    decBuf[2030] = 256'h0e0cf50bd40ba60b930b770b5d0b580b4c0b380b350b2b0b170b0f0bff0adf0a;
    decBuf[2031] = 256'hd10aab0a870a670a400a120af309d709b309a50998098509810978095e095409;
    decBuf[2032] = 256'h3e091e090009d608a308810855082e081e080708f207ee07e407ce07bf07a207;
    decBuf[2033] = 256'h78075c072307ef06bf06860661063f061f060e060906fb05ef05eb05d905b705;
    decBuf[2034] = 256'ha005710539051305d5049c047604460427041604fc03ee03ea03d703be03a203;
    decBuf[2035] = 256'h780345030703cd028a025c022202fd01e801e201dc01e201dd01d901c501a601;
    decBuf[2036] = 256'h6f012b01d9008c0046000600ccffa7ff92ff8cff92ff8cff88ff7bff50ff1eff;
    decBuf[2037] = 256'he0fe96fe3cfefffdb2fd80fd65fd5cfd64fd6bfd71fd6bfd5cfd32fd0bfdbefc;
    decBuf[2038] = 256'h5bfc18fcc3fb76fb30fb15fbfcfaf5fafcfaf5fafbfaecfacbfaa5fa62fa10fa;
    decBuf[2039] = 256'hc3f97df92bf9f4f8d6f8bbf8b3f8baf8b3f8c6f8aaf890f867f81df8d7f785f7;
    decBuf[2040] = 256'h22f7dff6a3f66cf64ef657f64ff656f65df64af639f616f6d9f5a0f55cf50af5;
    decBuf[2041] = 256'hd3f4a1f473f45bf462f44ef447f44df433f413f4f5f3bbf371f33ff3fff2c5f2;
    decBuf[2042] = 256'haff27ff26cf266f257f249f245f22af211f2fbf1d0f1a4f188f150f12af116f1;
    decBuf[2043] = 256'heaf0cef0bef095f079f069f040f024f014f0ebefceefbfef9fef81ef75ef4fef;
    decBuf[2044] = 256'h2bef14efe5eec6eeb5ee91ee71ee75ee5aee4fee59ee3fee2dee24eef9edcded;
    decBuf[2045] = 256'hb1ed79ed53ed3eed1fed0eed13ed0fed13ed26ed1ced19ed16edefecc7ecb8ec;
    decBuf[2046] = 256'h85ec63ec50ec34ec2fec46ec41ec45ec65ec58ec54ec58ec2fec08ecf8ebc5eb;
    decBuf[2047] = 256'ha3eb90eb74eb6feb86eb82eb95ebb5eba8ebacebb6eb94eb74eb67eb35eb12eb;
    decBuf[2048] = 256'h0cebf0eae0eaf8eaebeae7ea06eb02ebfeea10ebfaeaeceaf3ead0eab6eabbea;
    decBuf[2049] = 256'h95ea85ea93ea86ea8aeaaaeaa5eab9ead8ead4ead8eae9eacdeabaeab6ea8eea;
    decBuf[2050] = 256'h7dea82ea6bea78ea9beaa8eac6eaf9ea0deb20eb3ceb2deb1feb23ebf8eae8ea;
    decBuf[2051] = 256'hedeadfeaecea1eeb33eb5eeb9cebb5ebdaebefebe9ebd8ebddebb3eba3eba8eb;
    decBuf[2052] = 256'ha3ebb8ebebeb0dec45ec89eca4eccdecf3ececece6ecebecd2ecc4ecd1eccdec;
    decBuf[2053] = 256'hdeec0ded30ed5beda4edc2eddeed07eef1edf7edfeede2eddcedeaede6ed09ee;
    decBuf[2054] = 256'h3cee5eee96eedaeef5ee1fef44ef4bef51ef57ef47ef4cef61ef65ef85efbcef;
    decBuf[2055] = 256'he1ef12f056f072f09bf0cff0d6f0e9f005f115f12cf152f176f19ff1e9f11bf2;
    decBuf[2056] = 256'h48f292f2b0f2def218f32ef343f36ff38bf3aff3ebf314f449f479f4a4f4d7f4;
    decBuf[2057] = 256'h15f52ef562f592f5b2f5e4f514f640f673f6b1f6daf60ef73ef75ef785f7b3f7;
    decBuf[2058] = 256'hc6f7edf71bf847f86ff8a7f8ccf8fdf828f950f969f993f9a4f9bdf9def9fcf9;
    decBuf[2059] = 256'h26fa59fa89fac1faf6fa34fb5dfb91fba6fbc5fbe1fbf1fb11fc2ffc4afc77fc;
    decBuf[2060] = 256'hb0fce4fc14fd4dfd81fdb1fdd0fdedfd06fe27fe3cfe5ffe88febbfeebfe30ff;
    decBuf[2061] = 256'h70ffbaffecff2c0055007b008f00ae00bf00d90003012a016201a601e6011f02;
    decBuf[2062] = 256'h54028402b002cc02e602fd021a03360363038f03c103ff0339046e049e04c904;
    decBuf[2063] = 256'he604f5040c0519052c054c0569059405c705f7052306550678068a06a606ac06;
    decBuf[2064] = 256'hb006bd06c906e1060a07310769079e07ce0706082c0833085208580852086a08;
    decBuf[2065] = 256'h7f088a08b808f008250963099c09d109010a2d0a3e0a570a6e0a7b0a9e0ac80a;
    decBuf[2066] = 256'hef0a320b710bab0bef0b410c620ca80cd50cee0c140d360d550d7d0dab0dd70d;
    decBuf[2067] = 256'h140e4e0e740ebf0ef10e1f0f590f8d0fa20fce0ff50f0f102f10551065108510;
    decBuf[2068] = 256'hab10b010da100111111131114f115a1173118911801193119a118b1195119a11;
    decBuf[2069] = 256'h8b119d11a911a711c111d311d011de11e611d511d711cd11b311af11a5118f11;
    decBuf[2070] = 256'h9711a5119911b411c811c411da11e811db11e211dc11c211cd11c911bb11d311;
    decBuf[2071] = 256'hef11fa11211245125c1282129c129712a412a8129612a012a812a012c412e812;
    decBuf[2072] = 256'hf6122d13621368139413b013ab13b913bd13aa13b413be13bb13e2130a141914;
    decBuf[2073] = 256'h4c146e1468148f1495147414701464143e14391434141f143a144b144f146e14;
    decBuf[2074] = 256'h7b14681472146214371431141514e713ed13e713ce13ee13fb13f71310140c14;
    decBuf[2075] = 256'hf813f613e513c513b713a2138f13a013b013b313da130114071427142b141814;
    decBuf[2076] = 256'h22141f1405141714261435145c149a14c314071534154d1573157a1567156c15;
    decBuf[2077] = 256'h72155a158115a515bc15fb154e166f16b516d016d816e016cb169f168e167516;
    decBuf[2078] = 256'h54166a167d168816b616d916df16f016e116a4167b162916dc15961556151c15;
    decBuf[2079] = 256'h0615f114de14e414ca14a11479143714d21375132013a71255120c12ae11a211;
    decBuf[2080] = 256'h6b11391130110711c31095104b10f10fb50f520ff40ed00e990e670e4b0e320e;
    decBuf[2081] = 256'h1c0e150e020edb0dd60db50d870d740d4d0d1e0d180dfc0ce20ce70ceb0ce00c;
    decBuf[2082] = 256'hf80c020dff0c160d190d110d190d120dfe0cfc0cf00cdd0ce50ce20ce00cf60c;
    decBuf[2083] = 256'h050d0c0d220d250d1d0d1a0d070de50cce0ca80c7a0c670c400c260c180c030c;
    decBuf[2084] = 256'he80bdd0bc70b9c0b7d0b560b130be50a9b0a690a290a000abc09a10978094309;
    decBuf[2085] = 256'h21090209cf08ad08740831080308ca07860758071f07db06c006970671065c06;
    decBuf[2086] = 256'h3d062c061d060606f105dd05c505a2058b056d054b053d052705240527052a05;
    decBuf[2087] = 256'h3305400547054d0553054b053c052e051705fb04e804d604c704be04bb04be04;
    decBuf[2088] = 256'hc004ba04b504ad04990477044d041b04eb03a60366032c03f802c8029c026902;
    decBuf[2089] = 256'h39020102cc0181012701d2006f0011008cff0fffbdfe56fedefd8dfd43fde5fc;
    decBuf[2090] = 256'ha9fc46fce8fb93fb46fbc4fa6bfaf9f974f91bf9a9f85ff802f8c5f78ef75cf7;
    decBuf[2091] = 256'h2ef7f5f6cff691f658f623f6d7f591f564f52af505f5f0f4ddf4d8f4e7f4ecf4;
    decBuf[2092] = 256'hf8f413f517f51af51df50bf5faf4f8f4e6f4dff4f2f4faf414f541f561f588f5;
    decBuf[2093] = 256'hacf5c3f5d0f5dbf5d1f5bbf5b2f59bf58bf588f57bf57df58cf586f588f590f5;
    decBuf[2094] = 256'h7df565f54ff524f5ecf4c6f488f44ff429f4ebf3b2f38cf35cf324f3fef2c0f2;
    decBuf[2095] = 256'h87f261f223f2d9f1a7f167f11df1d7f085f038f006f0c6ef7cef5eef1eeff4ee;
    decBuf[2096] = 256'hedeecbeeabee9aee6cee41ee24eeecedb8eda3ed77ed66ed76ed71ed86eda9ed;
    decBuf[2097] = 256'hc0edd6edf1edededeaedededd0edbdedc0edb1edb9ede1edfded2bee70ee8bee;
    decBuf[2098] = 256'hb4eedaeee1eedaeee0eec6eea6eeaaee87ee83ee98ee94ee9feec1eebceeb0ee;
    decBuf[2099] = 256'hb3ee7fee4aee1aeebded5fed22edd5ec8fec62ec28ecf3ebdfeba7eb72eb42eb;
    decBuf[2100] = 256'he4ea87ea32eab9e947e9fde8a0e832e806e8c3e787e766e734e7f4e6dbe689e6;
    decBuf[2101] = 256'h3ce60ae6b7e56ae538e5f9e4cfe4d7e4b4e4bbe4d7e4d2e4e0e406e50be519e5;
    decBuf[2102] = 256'h37e53ae54ce57be58fe5afe5f8e516e656e6b0e6d5e622e77ce7b8e7efe749e8;
    decBuf[2103] = 256'h86e8bde817e954e98be9d1e9fee938ea8beaaceadeea30eb67ebadebffeb20ec;
    decBuf[2104] = 256'h52ec92ec9aeca1ecb6eca3ec92ec98ec80ec7cec90ec85ec8eecaeecaaeca6ec;
    decBuf[2105] = 256'ha9ec7bec4aec2becd7eb9aeb63eb1debf0eae7eac2eabbeac1eab0eaa1ea9cea;
    decBuf[2106] = 256'h65ea40ea0feacbe98be972e93ee929e93ce941e95be98ee9a2e9cee9f6e905ea;
    decBuf[2107] = 256'h0aea1fea1bea1eea41ea4fea75eac2ea0feb55ebcbeb1dec84ece2ec1eed55ed;
    decBuf[2108] = 256'hafedd4ed0bee51ee90eedbee49ef92ef0bf07df0e4f041f196f1e3f115f255f2;
    decBuf[2109] = 256'h7ef2a4f2d4f2f3f21bf35df38bf3b4f3f8f313f43cf462f469f47bf48cf47df4;
    decBuf[2110] = 256'h8bf498f484f488f497f489f48cf48ef47ff479f47bf469f462f464f452f44bf4;
    decBuf[2111] = 256'h4df43bf434f432f41cf419f41bf419f428f446f464f48ef4ccf4f5f439f579f5;
    decBuf[2112] = 256'ha2f5d7f507f626f659f696f6d0f614f778f7d6f743f8c8f821f993f9faf958fa;
    decBuf[2113] = 256'hacfaf9fa3ffb7ffbdafb2ffc92fc0afd7cfd01fe7efef0fe74ffceffffff4800;
    decBuf[2114] = 256'h8b00b000d100030130016a01ad01ed0138027e029902c202d902d202bf02ae02;
    decBuf[2115] = 256'h8a0273026602530257025a025d025f02580249022f020902db01a2016e013001;
    decBuf[2116] = 256'h0701d200b0009100740065004e0039001e00feffe0ffc5ffa6ff90ff7dff7aff;
    decBuf[2117] = 256'h70ff79ff86ff92ffa9ffbfffd3fff0ff13002a0050008900ae00ec0026016901;
    decBuf[2118] = 256'ha901e30126027902c6020c035e03c1031e047304ec043d05a50502065706ba06;
    decBuf[2119] = 256'hfd0652079f07f9074e089b0809095309b0091d0a670aaa0aff0a200b660b930b;
    decBuf[2120] = 256'hbd0bf10b210c410c7e0cb80cde0c0e0d460d5d0d7f0d9e0da40db30db80db40d;
    decBuf[2121] = 256'hc70dd10dce0de20dfa0d030e1d0e360e390e530e640e610e810e8e0e910eb80e;
    decBuf[2122] = 256'hdc0eea0e210f460f690fa10fd60ff80f301056106a10a310d710f9103e116c11;
    decBuf[2123] = 256'h9511e81135126712b912061338137813c213f41334146d149314df1425155215;
    decBuf[2124] = 256'h8c15c015e3150f162b1626163316381624162816251611161e161b1604160116;
    decBuf[2125] = 256'he715b2158d154115e714ab144814ea13ad1360131a13db12a1124e1201129311;
    decBuf[2126] = 256'h2c11b4102110980ff70e8b0e020e850d130dac0c690c140cb10b530be60a610a;
    decBuf[2127] = 256'h080a7609140996084508fb07d3079707760758073c071307ee06cb0686066b06;
    decBuf[2128] = 256'h42061c0615061c061606440670068c06c406f9061b0754078807aa07ef072f08;
    decBuf[2129] = 256'h5808ba0817095409b709150a510ab40a120b4f0bb20b0f0c640cc70c3f0d910d;
    decBuf[2130] = 256'hf80d560e920ef50e380f750fc20f08104810a210f7102e118811dd1114125a12;
    decBuf[2131] = 256'h88129012b512ca12d012ec12101327135f139313c313081436144e1474147b14;
    decBuf[2132] = 256'h68146e1469145114671482148c14bb140715251565158e15a415b915bf15ae15;
    decBuf[2133] = 256'hb415af159a15bd15dd15fb1535169016b41617173f1763178417a2179917a217;
    decBuf[2134] = 256'ha917a217c117de17ed1720184218481870187f1868186c1849180d18f517c017;
    decBuf[2135] = 256'h7417561729170017da16b8167f165a161c16d21578150b15a3142b1499130f13;
    decBuf[2136] = 256'h921200127711d6103e10b50f380fa60ef50d7e0dbc0c050c5f0b9c0ae5093f09;
    decBuf[2137] = 256'h7c08c5071f075c06da0534059c04ec037503dd022d02b601f3007100cbff33ff;
    decBuf[2138] = 256'haafe2dfebbfd54fdf6fc89fc3ffcfcfbc0fb89fb6bfb3dfb14fbeefaccfaadfa;
    decBuf[2139] = 256'h9cfa8cfa88fa9dfac0faeafa27fb72fbb8fb0afc57fc89fcc9fc02fd37fd67fd;
    decBuf[2140] = 256'hacfdecfd46feccfe49ffbbff5d00f4007e01fb016d02d40231038603d3032d04;
    decBuf[2141] = 256'h8204e5045e05f0057906f6068907eb076808b908e50828094d096e09a009df09;
    decBuf[2142] = 256'h2a0a980ae10a5a0bab0b120c550c7a0c9b0ca50cae0cb60cbd0cd20cf10c190d;
    decBuf[2143] = 256'h510d860dc30dfd0d230e450e580e5d0e6d0e710e650e700e7b0e840ea40ec20e;
    decBuf[2144] = 256'hd50efb0e150f230f380f440f470f510f4e0f3b0f390f260f090ffd0ee50ec90e;
    decBuf[2145] = 256'hbd0eac0e960e8d0e7b0e650e4c0e250ef70dbf0d6c0d1f0dc50c700c0d0cca0b;
    decBuf[2146] = 256'h5d0b140bd10a640a1a0aa1093009ab082e087b07d50612065b05b5041e046d03;
    decBuf[2147] = 256'hf6025f02ae013801a000f0ff1aff8afe9ffdc2fcf8fb0dfb6ffa6cf9bef820f8;
    decBuf[2148] = 256'h57f7a0f6f9f562f5b1f40bf449f392f2bcf12cf175f0cfef0cef8aee13eea7ed;
    decBuf[2149] = 256'h45edebec7aec30ecd2eb7deb30ebeaea98ea61ea2fea02eaf9e9f2e9ebe9fee9;
    decBuf[2150] = 256'h1aea29ea53ea7aea9eead1ea0feb49eb8cebf1eb4eecbbec23ed9bed0deeafee;
    decBuf[2151] = 256'h1befa4ef45f0b1f03bf1dcf148f2f8f29ff30bf494f435f5ccf556f6d3f645f7;
    decBuf[2152] = 256'hc9f747f8b8f83df9baf92cfab1fa2efba0fb07fc64fcb9fc06fd4cfd7afdb4fd;
    decBuf[2153] = 256'he8fd18fe5dfe8bfec4fef9fe29ff3cff58ff72ff76ff72ff76ff6bff68ff71ff;
    decBuf[2154] = 256'h79ff85ff98ffa5ffb1ffbbffadff9eff86ff64ff43ff26ff0bff00ff03ff06ff;
    decBuf[2155] = 256'h18ff33ff3dff40ff43ff2bff0fffecfec3fe90fe6efe5bfe4afe4ffe54fe50fe;
    decBuf[2156] = 256'h5bfe51fe3bfe1bfedcfd9cfd51fd0bfdb9fc82fc3cfcfcfbe4fbaffb71fb48fb;
    decBuf[2157] = 256'hf6fa93fa35fab0f932f9c1f83cf8bff74df7c8f64bf6faf575f5d4f468f4b8f3;
    decBuf[2158] = 256'h11f37af2a2f1d9f056f080eff1ee3aee94edd1ec4eeca8ebe5ea63ea8de9c4e8;
    decBuf[2159] = 256'h41e89be704e77ae6d9e542e5b9e43be4a9e347e3a6e23ae2d8e15be1e9e09fe0;
    decBuf[2160] = 256'h5ce020e0ffdfcddf9fdfa7df91df8adf9ddf97dfa7dfd9dfeedf26e088e0cbe0;
    decBuf[2161] = 256'h38e19fe117e289e22be398e321e4c2e459e5e3e583e61be7cbe772e834e9ebe9;
    decBuf[2162] = 256'hc1ea8aeb41ec17eda7ed5dee33efc3ef46f0ecf083f134f2daf271f322f4c8f4;
    decBuf[2163] = 256'h34f5bef53bf68cf6d6f619f73df774f7a6f7c2f7ebf72ef84af862f888f88ff8;
    decBuf[2164] = 256'h7cf876f834f8f4f7cbf778f741f70ff7e2f6b8f693f670f645f61df6d0f583f5;
    decBuf[2165] = 256'h3df5d9f496f441f4f4f3c2f3a7f38ef387f38ef37bf375f370f359f344f338f3;
    decBuf[2166] = 256'h20f316f325f337f35bf39df3ddf317f469f4a0f4d2f412f53bf561f59ff5c8f5;
    decBuf[2167] = 256'hfdf556f693f6f6f653f7a8f7f5f73bf869f892f8b7f8b1f8b7f8d3f8c4f8c8f8;
    decBuf[2168] = 256'he6f8e2f8edf802f9eef8dcf8c7f89bf83ef8fbf78ef709f7b0f63ef6d7f579f5;
    decBuf[2169] = 256'h0cf5a5f447f4daf355f3d8f246f295f11ef15cf0a5efffee67eedeed3dedd1ec;
    decBuf[2170] = 256'h47eceeeb5cebfaea7dea0beaa4e946e9c1e867e816e8cce789e765e75ae750e7;
    decBuf[2171] = 256'h6be784e7aae7e7e711e845e883e8bde800e952e99fe921ea9fea31ebe1eb88ec;
    decBuf[2172] = 256'h4aed01eea7ee6aef21f0f7f0c0f177f21df3e0f3cbf4a8f571f628f7fef7c7f8;
    decBuf[2173] = 256'hb2f990fa20fbd6fb7dfc14fd9dfd3efeaafe34ffb1ff02008700e00032015e01;
    decBuf[2174] = 256'ha101ad01ce01d801bc01b4019e016e0142011a01d80098005e000c00bfff65ff;
    decBuf[2175] = 256'hf8fe90fe33feadfd30fdbefc57fcdffb6dfb06fb8dfa3cfad5f977f93bf9eef8;
    decBuf[2176] = 256'ha8f868f83ff80af8e8f7c8f7b8f7b2f7caf7e7f712f850f8abf8fff84cf9baf9;
    decBuf[2177] = 256'h22fa9afa0cfb91fb0efca0fc29fdcafd8dfe44ff1900e3009a016f023903ef03;
    decBuf[2178] = 256'h960458050f06b5064d07fd0774083709b909600acc0a550bd20b440cab0cee0c;
    decBuf[2179] = 256'h430d640d960db10dba0db20d9e0d7e0d570d290df10cad0c6d0c230cc90b740b;
    decBuf[2180] = 256'hfb0a890a220a8f0906098808d6075f07c8063e06c1054f05cb047104ff039803;
    decBuf[2181] = 256'h3b03cd02660209029b0134010c01cf00ae00b800c200da00000130015c019a01;
    decBuf[2182] = 256'hd301f90144028a02dd025603c7034c04ed0484053506db069e072008f6088609;
    decBuf[2183] = 256'h3d0ab40a760b2d0cd30c6b0d1b0ec20e840f0710ad101911a311fc116e12b712;
    decBuf[2184] = 256'hfa124f138613b813e613ff1324142b1425141414f013c61388134f13fc12af12;
    decBuf[2185] = 256'h5512e811811123119e102110af0f0d0fa10e170e760ddf0c560cd80b460bbd0a;
    decBuf[2186] = 256'h400ace094909a8086708de0785073307cc06890665062e06fc050506fd05f505;
    decBuf[2187] = 256'h0a0629063a067206b606e4062e079c07e6075e08d0083709e5098b0af70aa80b;
    decBuf[2188] = 256'h4e0c110dc80d6e0e300fe70fbd104d1138121513df1395146b153416eb16c117;
    decBuf[2189] = 256'h51180819ae191a1aa31a211b921b171c701cc21c291d871dc31d101e421e5e1e;
    decBuf[2190] = 256'h871e8e1e6c1e661e3e1e061ed11d941d491d031db11c4e1c0b1cb61b3d1bec1a;
    decBuf[2191] = 256'h671aea195819cf182e18c21711176b16ff157515f81486141f14a7135613ee12;
    decBuf[2192] = 256'h76122512db1163113211e8108a10661045102710301038103110531066106c10;
    decBuf[2193] = 256'h90109d10a210c510dc10f1102b117511bb1120129812e9125113ae13eb132214;
    decBuf[2194] = 256'h54146f1488149e14a514c514ec1406152f15571570157e157a1557152415d814;
    decBuf[2195] = 256'h7e141114aa134c13df1296121d12cc1182110a119810f60f5e0f870ebd0dd20c;
    decBuf[2196] = 256'h340c310b830ae5091c09990822088b0701078406f2056905c804300480030903;
    decBuf[2197] = 256'h7202e801b301610118010a01fe00f300fd0006010f0125013a0133015b017f01;
    decBuf[2198] = 256'h9f01df0131027e0200037d030f0499043a05d10582062807bf077008e7087e09;
    decBuf[2199] = 256'h070aa80a140bc50b6b0c030db30d590ef10ea10f4810b41016116f11a011ea11;
    decBuf[2200] = 256'h2d1251128812ce120e135813b2130714541486148f14971472142614cc137713;
    decBuf[2201] = 256'hfe12ad1246120312c6118f115d113011f61095101c108a0fd90e330e700d850c;
    decBuf[2202] = 256'he70b570ba10a2a0abe095c09020990080c088f07dc0606063d055204b403ea02;
    decBuf[2203] = 256'h3302bd017c011a01e400b3006a002700d2ff43ffb9fe19fe81fdf8fc9efc4dfc;
    decBuf[2204] = 256'h21fc14fc20fc2bfc49fc52fc4afc33fcf5fbabfb65fb01fbbefa81fa4afa40fa;
    decBuf[2205] = 256'h49fa51fa68fa7dfa83fa88fa6ffa3cfafef9b4f95af905f9b8f85ef821f8eaf7;
    decBuf[2206] = 256'hb8f78bf751f7fef6c7f659f6f2f57af5e8f45ef4bdf326f39df21ff2aef146f1;
    decBuf[2207] = 256'he9f07cf014f0b7ef62efe9ee98ee13ee96ed24ed9fec22ecb0eb49eb06ebcaea;
    decBuf[2208] = 256'h93ea89ea80ea88ea8feab2eab8eac9eae2eae7eaf4ea0feb27eb56eba2ebfceb;
    decBuf[2209] = 256'h69eceeec6bedfdedaeee25efbcef45f09ff0f0f057f1b5f13af2b7f24af3d3f3;
    decBuf[2210] = 256'h98f44ef5f5f5b7f63af7b1f71df87ff8d8f809f953f97bf9d0f91dfa77fafcfa;
    decBuf[2211] = 256'h56fba7fb0efc36fc5bfc66fc48fc1afcf1fb9efb67fb35fb08fbeffaf6faeffa;
    decBuf[2212] = 256'he9fafafad6faadfa85fa38fabff94ef9c9f84cf8daf773f715f7d8f6a1f65bf6;
    decBuf[2213] = 256'h1cf6c1f56cf509f591f4fef39cf3fbf264f202f2a8f137f10af1c8f08bf054f0;
    decBuf[2214] = 256'h22f0e2efa8ef47efe9ee94ee31eeb9ed88ed21eddeecbaec83ec65ec5cec32ec;
    decBuf[2215] = 256'h1cec15ecf6ebdaebd4ebabeb83eb74eb4aeb3aeb34eb27eb2beb46eb57eb74eb;
    decBuf[2216] = 256'haeebc6ebddeb1bec23ec2bec31ec2bec1aec1fec08ec04ec1fec2aec4cec88ec;
    decBuf[2217] = 256'ha1ecc6ec04edfcec04ed18edf9ecddecd8ecaeeca8ecb8ecaaecbfece2ece7ec;
    decBuf[2218] = 256'hfcec08edf6ecdaecbfec8aec56ec41ec15ec05ec14ec19ec47ec80eca5ece3ec;
    decBuf[2219] = 256'h0ced23ed45ed64ed5fed6eed8eeda4edd6ed22ee68eeccee44ef96ef1af074f0;
    decBuf[2220] = 256'he6f04df1c5f116f29bf218f38af30ff48cf41ef5cff575f60cf796f737f8cef8;
    decBuf[2221] = 256'h57f9d5f946faaefa26fb77fbdefb57fca8fc0ffd88fdd9fd40fe9efedafe11ff;
    decBuf[2222] = 256'h43ff5fff78ff7fff78ff72ff6cff5dff58ff54ff41ff36ff2dff0dffe7fec3fe;
    decBuf[2223] = 256'h7efe38fee6fd83fd25fdd0fc83fc29fcecfbb5fb83fb56fb2dfbf8fad6faaafa;
    decBuf[2224] = 256'h77fa55fa1dfaf7f9d5f9b6f999f98af985f981f97df981f97ef986f989f98bf9;
    decBuf[2225] = 256'h92f998f9a7f9bbf9cdf9e7f90efa31fa5bfa8efabefaf6fa2bfb4dfb85fbabfb;
    decBuf[2226] = 256'hcdfbecfb08fc18fc26fc3bfc3ffc50fc60fc69fc7bfc90fc99fca6fcb7fcb5fc;
    decBuf[2227] = 256'hb3fcadfc9ffc8dfc81fc72fc64fc5ffc5afc5efc62fc64fc67fc64fc59fc4afc;
    decBuf[2228] = 256'h38fc1efc05fcf6fbe7fbe0fbddfbe4fbeefbfafb08fc1afc26fc35fc43fc53fc;
    decBuf[2229] = 256'h62fc80fc9efcc0fcf3fc23fd5cfd9ffddffd19fe5cfe9cfec5fe09ff49ff83ff;
    decBuf[2230] = 256'hc6ff060040009200df0025018a01cc013a02a102fe025303cc031e048504e204;
    decBuf[2231] = 256'h50059905f70534068106db0617077a07bd0712087508b8080d0944098a09b709;
    decBuf[2232] = 256'he109f709190a390a550a790a990ab70ad20ae30af30aea0add0ac30a960a6a0a;
    decBuf[2233] = 256'h2c0af209af096f0935090109b5086f082f08d40780071d07bf06520608069005;
    decBuf[2234] = 256'h3e05f504970442040b04c50373033c03e2028d0256021002d001a70182015f01;
    decBuf[2235] = 256'h5901530144014901550151016a0180019a01c701f30131027b02d5022a038d03;
    decBuf[2236] = 256'heb033f048c04e6043b058805e2051f066c06c606030750079607d5070f085308;
    decBuf[2237] = 256'h8008aa08de08f30812092e093d095509590955094a093b091b09fd08d308a008;
    decBuf[2238] = 256'h70083808f407b4077b072807db0695064306e00582052e05e10487043204fb03;
    decBuf[2239] = 256'hc9039b0382035d033a0328030c03f202e402d702bc02c002c902cc02e4020603;
    decBuf[2240] = 256'h1d0354038903b903fe033e047704bb040d0544059e05f30540069a0607075107;
    decBuf[2241] = 256'hae071b088308e00835098209c8091a0a510a830ac30aec0a120b340b540b700b;
    decBuf[2242] = 256'h890ba00bb60bba0bbd0bba0bb10b9a0b7e0b5b0b310b0a0bdc0ab00a880a650a;
    decBuf[2243] = 256'h320a020ac90986094609fc08a2084d08ea078c073707ea06a40677063d06f905;
    decBuf[2244] = 256'hcc0592054f050f05c4047e043f04f403c20395036b03550340032e0311030203;
    decBuf[2245] = 256'heb02c502a102770250022c02150208020c021d022d0258028402a002ce02ed02;
    decBuf[2246] = 256'h0a0323033a0347035a0373038303a803d603020440047904ae04ec0426054b05;
    decBuf[2247] = 256'h8905b205d805fa052606420670069c06c306f1062a074f077f07ab07c707eb07;
    decBuf[2248] = 256'hf907f507f107e607d007b607a507890775076b075507470734071a07fb06d406;
    decBuf[2249] = 256'h9c0668062a06f005ca059a0562054c05370524051f0519050205f604da04b404;
    decBuf[2250] = 256'h9a047a0454044404360432043e04560466049104bd04d90407053f0556059405;
    decBuf[2251] = 256'hbd05e20520065a069e06dd0628076e07ae07f8072a0857088108a608bb08da08;
    decBuf[2252] = 256'he008ef08fd080a0915092009230926091e091709ff08dd08b30881084308f907;
    decBuf[2253] = 256'h9f074a07fd06a3063606ec058e053905ec0492043e04db036203f0026c021202;
    decBuf[2254] = 256'h80011e01c50053000900c6ff8aff53ff21fff3fecafeb3fe91fe65fe49fe2ffe;
    decBuf[2255] = 256'h18fe14fe18fe1bfe37fe5afe7bfeb2fee6fe17ff4fff83ffb3ffdfff1d005700;
    decBuf[2256] = 256'h9a00da0014016601b3010d026202af02e10221035b038f03b203c503d503ef03;
    decBuf[2257] = 256'hfd0312041e042f043f0453046004630460045a044b042f040c04e303b0038003;
    decBuf[2258] = 256'h48031303e302b7028502540229020102c901940157011d01d900990060003a00;
    decBuf[2259] = 256'h0a00ebffcfffb5ffa7ff9aff87ff7dff67ff58ff41ff31ff23ff1bff1dff28ff;
    decBuf[2260] = 256'h36ff4dff69ff8cffa3ffc9ffe3fffaff06001a002b0041005b0074009c00c400;
    decBuf[2261] = 256'hf2002a015e019c01d601fc012c024b026702810298029c02a802ab02b502b702;
    decBuf[2262] = 256'hba02bc02c302c102bc02b302a3028c027602500222020302d001a00168013301;
    decBuf[2263] = 256'h0301cb00880048000e00bbff6eff14ffa7fe40fee2fd8efd2bfdcdfc78fc15fc;
    decBuf[2264] = 256'hb7fb63fb00fba2fa4dfaeaf9a7f93af9f0f893f856f809f8c3f795f75cf736f7;
    decBuf[2265] = 256'h22f7f6f6daf6caf6b3f6a6f69bf690f68df68af692f69ef6adf6bff6d9f6f2f6;
    decBuf[2266] = 256'h0ef738f760f798f7cdf70af855f89bf8dbf825f96bf9abf9e4f928fa56fa8ffa;
    decBuf[2267] = 256'hd3fa00fb3afb6ffb91fbbdfbe4fbfefb27fc44fc5dfc74fc92fc96fc99fca9fc;
    decBuf[2268] = 256'ha0fc99fc8dfc6dfc4cfc26fceefbb9fb89fb51fb1cfbecfab4fa80fa4ffa17fa;
    decBuf[2269] = 256'he3f9b3f96ef92ef9f4f8a2f855f823f8d1f79af768f728f7fef6d9f6a9f67df6;
    decBuf[2270] = 256'h6cf648f631f624f619f61cf61ff622f62ff645f64df660f67ff68bf6a7f6cdf6;
    decBuf[2271] = 256'he7f610f743f765f79ef7d2f710f84af87ef8aef8e7f82af958f981f9b5f9d8f9;
    decBuf[2272] = 256'hf7f92afa3efa51fa6dfa72fa80fa8dfa89fa8dfa96fa93fa96fa98fa89fa7bfa;
    decBuf[2273] = 256'h76fa5efa37fa1dfaebf9baf98ff951f907f9d5f895f84af818f8c6f779f747f7;
    decBuf[2274] = 256'h07f7bdf68bf64bf612f6ecf5bcf590f569f530f5fcf4ccf487f459f420f4ebf3;
    decBuf[2275] = 256'hc9f3b6f3a5f3a0f3a5f3b1f3c5f3ddf3edf301f413f416f420f42ef434f442f4;
    decBuf[2276] = 256'h58f46cf48ff4b8f4e0f418f54cf57df5b5f5f8f526f660f6a3f6d1f60bf74ef7;
    decBuf[2277] = 256'h8ef7c8f7fcf72cf858f88bf89ff8cbf8e7f8f7f80ef934f943f964f992f9a5f9;
    decBuf[2278] = 256'hcdf9fbf91afa41fa65fa7cfa89fa9cfa92fa95fa98fa80fa77fa74fa67fa69fa;
    decBuf[2279] = 256'h70fa72fa81fa99faa2fab1fabefabbfab9fab7faa0fa91fa82fa66fa52fa4ffa;
    decBuf[2280] = 256'h3ffa3cfa3ffa3cfa43fa4dfa4bfa50fa5dfa63fa75fa8afa9efabbfadefafefa;
    decBuf[2281] = 256'h1cfb37fb49fb5efb6dfb6ffb77fb79fb7ffb8bfba3fbc3fbf2fb2afc5efcaafc;
    decBuf[2282] = 256'hf0fc30fd6afdadfdc8fdf2fd17fe2cfe3ffe44fe54fe61fe7ffe93feabfed4fe;
    decBuf[2283] = 256'hfbfe1fff49ff70ff8affa1ffb6ffc2ffc5ffbcffb3ffa6ff91ff7cff6aff55ff;
    decBuf[2284] = 256'h41ff33ff1eff0afff8fee7fed8fec6feb5fea7fe99fe8cfe84fe7afe70fe65fe;
    decBuf[2285] = 256'h51fe3ffe2efe13fef8fdd8fdc3fdaffda5fda2fdb0fdcdfdf0fd1afe4cfe8afe;
    decBuf[2286] = 256'hb3fef7fe24ff3dff63ff85ff98ffb4ffceffeeff140042007b00be0010015d01;
    decBuf[2287] = 256'hb7010c025902b302f0023d038303c303fc03220452047e04a504c904e904ff04;
    decBuf[2288] = 256'h1a052b0541055505680582059a05b605d905fa0517063a065106670672066806;
    decBuf[2289] = 256'h58063e061806f405c1059105720555053c0537053b053f0558056e0576058905;
    decBuf[2290] = 256'h8b05800576056705470530051a05ff04f504f204ef040605230536055c058b05;
    decBuf[2291] = 256'haa05d105f50515063c0660066d068b06a606b806d406e706f20608071c072907;
    decBuf[2292] = 256'h43075c0771079d07c807f00728085d088d08d108ff0828094e09620969096e09;
    decBuf[2293] = 256'h690952093d0922090909fa08f108ee08fa080d0920093f095409670979098809;
    decBuf[2294] = 256'h80097d09710951093a091409e608c708aa087c085d0841082708190815080208;
    decBuf[2295] = 256'h050808080608130810080a080c080308eb07e007ca07a50796077f0769076507;
    decBuf[2296] = 256'h69076c078607a507c307f607260851088408b408d308060928092f0956096509;
    decBuf[2297] = 256'h73098909a409b509e409140a400a890acf0a0f0b6a0bbf0bf60b3c0c7b0ca50c;
    decBuf[2298] = 256'hd90cee0c010d110d210d1c0d200d2c0d220d310d3a0d3c0d4d0d5c0d620d750d;
    decBuf[2299] = 256'h820d850d8f0d890d730d630d430d0c0de70ca90c5e0c180cd90b7e0b410b0a0b;
    decBuf[2300] = 256'hc40aa90a800a4b0a360a240afc09e309cc09a5098c096b0934090f09de08a608;
    decBuf[2301] = 256'h8108510818080208ed07ce07d407d907dd070408270848087708a208b308d708;
    decBuf[2302] = 256'hee08f20806091009130928093a094b096a099d09cd09060a3a0a6a0aa30ad70a;
    decBuf[2303] = 256'h070b330b4f0b5e0b760b7a0b6e0b6b0b550b350b200b050be50ad90abd0aac0a;
    decBuf[2304] = 256'ha90a9a0a8d0a8b0a800a6a0a560a2f0afc09cc0987094709fd08a3084e080108;
    decBuf[2305] = 256'ha70752070507bf06800646062006f005dd05c105a8059a058505690551053505;
    decBuf[2306] = 256'h0205e004b40482045f0440042404150419041d043104490465049004b704d104;
    decBuf[2307] = 256'hfb0422053c055c057a058d05ad05c205d505ee05fd0512062906450660068e06;
    decBuf[2308] = 256'hba06e10619074e0770079c07b807c807d507d107b607a5078207590731070307;
    decBuf[2309] = 256'hd706bb0697068006620647062f061906f905d305af057c053e05f4049a044504;
    decBuf[2310] = 256'he2036a03f80291021902c70160010201c6008f0049000900cfff8cff4cff12ff;
    decBuf[2311] = 256'hc0fe73fe2dfedafd8dfd47fd08fdbdfc8bfc4bfc12fcecfbbcfb9dfb8cfb7dfb;
    decBuf[2312] = 256'h78fb7cfb80fb99fba8fbbcfbc9fbd5fbdcfbe2fbdcfbd8fbd9fbdafbdefbeffb;
    decBuf[2313] = 256'h04fc1efc45fc73fc9ffcd1fcf4fc2cfd51fd66fd85fd96fda6fdaafdaefda3fd;
    decBuf[2314] = 256'h91fd88fd74fd61fd56fd42fd35fd2efd1ffd11fd09fdf3fcdafcbafc8bfc60fc;
    decBuf[2315] = 256'h22fcd7fb7dfb41fbdefa80fa2bfab2f961f9faf89cf847f810f8caf778f757f7;
    decBuf[2316] = 256'h11f7e4f6baf686f648f60ef6bcf56ff515f5c0f45df41af4c5f38ef35cf32ef3;
    decBuf[2317] = 256'h26f31ff326f32cf33df34cf351f366f362f36df37cf37ff387f3a1f3acf3c1f3;
    decBuf[2318] = 256'hedf3fff31bf43ff456f474f4a7f4bbf4e7f41af53cf55bf58ef5a2f5c2f5e9f5;
    decBuf[2319] = 256'heef5eaf5f6f5e3f5d1f5cef5aff599f596f576f561f55df544f535f532f515f5;
    decBuf[2320] = 256'hfaf4e8f4baf47cf452f400f4b3f359f304f3a1f243f2eff18cf149f10cf1d5f0;
    decBuf[2321] = 256'ha3f075f03cf025f0e7efaeef79ef3beff1eebfee7fee35ee17eed7ed9ded78ed;
    decBuf[2322] = 256'h48ed1ced00eddcecbbecb7eca4ec99eca9ecacecbeece2ecf1ecffec1ded21ed;
    decBuf[2323] = 256'h2bed41ed38ed3bed50ed53ed66ed89edadedd7ed20ee52ee92eeccee00ef30ef;
    decBuf[2324] = 256'h68ef8eefb0efdcefe2eff1ef1bf02cf03bf06ef082f0a2f0d4f0f7f016f154f1;
    decBuf[2325] = 256'h6df183f1b3f1b9f1bff1d9f1cbf1c7f1caf1c0f1c3f1ccf1bff1c1f1d0f1c6f1;
    decBuf[2326] = 256'hc1f1c5f1b2f1a0f19df186f176f17ff172f16ff17af16cf167f165f14ff12cf1;
    decBuf[2327] = 256'h15f1e6f0bbf09ef07bf06df071f06df07ff0a7f0c3f0ddf007f123f132f149f1;
    decBuf[2328] = 256'h3cf140f144f141f144f151f158f16ff19ef1c0f1e0f11ef247f27bf2b9f2e2f2;
    decBuf[2329] = 256'h17f355f37ef3b3f3e3f302f435f465f484f4b7f4e7f412f545f575f594f5c7f5;
    decBuf[2330] = 256'h05f61ef652f682f6aef6d5f60ef724f747f77ff795f7aaf7bdf7c2f7c8f7ccf7;
    decBuf[2331] = 256'hbff7c3f7d5f7d8f7ecf70ef825f854f88cf8a3f8c5f8e4f8eaf8eff8f4f8dff8;
    decBuf[2332] = 256'hd3f8c8f8b9f8b6f8bef8c5f8d4f8eef8fff81bf937f948f964f97ff998f9b4f9;
    decBuf[2333] = 256'hcff9eff90cfa37fa53fa77fa97faadfacffae7fafcfa1ffb3ffb65fb93fbbffb;
    decBuf[2334] = 256'hf2fb30fc69fc9efcdcfc16fd4afd7afdb2fdd8fd08fe34fe50fe7efeaafec6fe;
    decBuf[2335] = 256'hf4fe20ff52ff90ffcaff0e006000ad00f30033016c01a101c301e201ff010e02;
    decBuf[2336] = 256'h1c0231024c026c029202c002ec022a0363038903b903f1031704390458047504;
    decBuf[2337] = 256'h8e04a504b204cd04df04e204f004f804fa04050513051f0538055e057805a105;
    decBuf[2338] = 256'hd405e9051406310640064e065b064f0652064f064c064f0656065d0673068c06;
    decBuf[2339] = 256'h9e06c006ea0606072a07540770079e07ca07da07fe0715082208360840083d08;
    decBuf[2340] = 256'h5108630874089408be08e5081d0952097409ac09e109030a3c0a610a830aaf0a;
    decBuf[2341] = 256'hcb0ae50a050b230b2f0b4e0b630b670b800b9c0baf0bd60b040c300c6e0ca70c;
    decBuf[2342] = 256'hcd0cfd0c290d450d540d590d4c0d480d370d1b0d170d1a0d110d250d370d3e0d;
    decBuf[2343] = 256'h5e0d880d990dbd0dd40de10d030e1b0e1f0e3a0e440e3b0e3e0e360e1c0e180e;
    decBuf[2344] = 256'h0f0efb0d030e130e160e340e6b0e810ebf0ef90e0f0f400f6b0f7c0f960fa40f;
    decBuf[2345] = 256'h9f0fb30fc40fc10fdb0ff40ffd0f221046105d108c10c410db10191142116711;
    decBuf[2346] = 256'h8a11a911af11be11cc11b711bb11b711a111a411a711a011b311c011b911d011;
    decBuf[2347] = 256'hd911d111d911d611bf11c211ae11911185116d1144112811fa10c2108d105d10;
    decBuf[2348] = 256'h0c10eb0fb90f790f710f5a0f460f4c0f520f420f470f320f070feb0ebd0e840e;
    decBuf[2349] = 256'h500e200ee80dc20da00d800d7b0d760d680d750d800d7d0d990da40da80db80d;
    decBuf[2350] = 256'hc00db30dbf0db40d9a0d970d870d6d0d6a0d670d580d6b0d800d890db00dd70d;
    decBuf[2351] = 256'he70d070e1c0e200e320e350e210e190e040ee40dd70dbc0d960d860d660d400d;
    decBuf[2352] = 256'h3a0d2d0d170d1b0d180d0e0d170d1a0d040d010de40cb20c900c570c050cce0b;
    decBuf[2353] = 256'h880b480b1f0bf90ac90ab60ab10a970a930a860a720a680a5f0a3f0a320a170a;
    decBuf[2354] = 256'hf109d709b709900977094d0926090c09ec08ce08c208b808b508c908d608e208;
    decBuf[2355] = 256'h020922092f094a0954095809600953093e09350923090d09ff08ed08d708d408;
    decBuf[2356] = 256'hd708d508e808fa080b092609410953095c095f094d0937091209da08a5086708;
    decBuf[2357] = 256'h2e080808d807ac07900776075f075b07480728070a07e006ad066f063606e305;
    decBuf[2358] = 256'h96055005ec04a90454040704c1036f032203f002b002760251022102f501cd01;
    decBuf[2359] = 256'haa01800159012a01f200be00800036000400c4ff8aff64ff34ff09fff8fedefe;
    decBuf[2360] = 256'hd9fedefee2feecfe02ff10ff23ff38ff46ff4eff55ff53ff4dff45ff39ff32ff;
    decBuf[2361] = 256'h30ff34ff3cff4bff62ff85ffa5ffc3ffdefff6ff060014001700190013000500;
    decBuf[2362] = 256'hf5ffe6ffd4ffbaffa9ff8dff72ff59ff3dff22ff09ffe7fec7febafe9ffe7ffe;
    decBuf[2363] = 256'h6afe3ffe18feeafdb2fd6efd2efde4fc9efc5efc14fccefba0fb77fb51fb3dfb;
    decBuf[2364] = 256'h2afb24fb15fb10fb04fbf0fadffabcfa9cfa76fa48fa1cfa00fadcf9cef9c1f9;
    decBuf[2365] = 256'hc5f9d0f9e6f9fff926fa54fa73fa9bfab4fad5faeafaf6fa00fb09fb0cfb14fb;
    decBuf[2366] = 256'h25fb2bfb31fb48fb51fb60fb77fb81fb89fba1fba4fbb2fbc5fbc7fbc9fbd3fb;
    decBuf[2367] = 256'hcbfbbcfbb2fb98fb65fb43fb0bfbc7fa9afa4ffa1dfaf0f9b6f990f96ef942f9;
    decBuf[2368] = 256'h1bf901f9cef89ef873f829f8e3f7a4f749f7f4f6a7f64df6f8f5c1f57bf54df5;
    decBuf[2369] = 256'h24f5f0f4cdf4bbf49ef485f46ef450f435f41cf4faf3e3f3c5f3a2f382f36df3;
    decBuf[2370] = 256'h51f340f33df334f337f347f352f36cf393f3b6f3e0f313f443f47bf4b0f4d2f4;
    decBuf[2371] = 256'hf1f419f51ef52cf549f545f550f566f574f58cf5b4f5d1f5fff543f671f69af6;
    decBuf[2372] = 256'hdef6f9f622f739f740f746f74cf732f71bf717f7fcf6e3f6daf6c6f6b8f6bbf6;
    decBuf[2373] = 256'hacf6a2f69df684f66cf65cf631f612f6eaf5bcf584f55ff52ef503f5e7f4aef4;
    decBuf[2374] = 256'h7af465f42df407f4e5f3c6f39ef38ff378f363f35ff34df344f347f334f328f3;
    decBuf[2375] = 256'h26f314f308f302f3f4f2f2f2faf2fff214f333f351f383f3c1f3eaf31ff45df4;
    decBuf[2376] = 256'h97f4cbf4fbf41af542f570f58ff5abf5cff5f0f50df640f662f68ef6c0f6f1f6;
    decBuf[2377] = 256'h1cf75af783f7a9f7d9f7ecf7fdf716f812f816f81af808f8f9f7f0f7d8f7c3f7;
    decBuf[2378] = 256'hbaf79df78af77ff75df746f739f70ef7f2f6d9f6aff67cf65af62ef6f0f5c7f5;
    decBuf[2379] = 256'h84f544f51af5d7f4a9f480f45bf438f425f409f4faf3f5f3e0f3d4f3caf3b4f3;
    decBuf[2380] = 256'ha0f393f374f35ff353f349f345f34ef351f36bf391f3abf3d5f312f43cf470f4;
    decBuf[2381] = 256'haef4d7f40cf54af573f598f5c9f5e8f50ff63df669f690f6c9f6fdf62df772f7;
    decBuf[2382] = 256'hb2f7ecf72ff86ff8a9f8ecf81af954f988f9abf9caf9fdf911fa24fa35fa3afa;
    decBuf[2383] = 256'h48fa4cfa48fa4cfa55fa52fa5ffa70fa7bfa8dfaa2faa5fab2fabefaaffa9dfa;
    decBuf[2384] = 256'h8cfa6cfa43fa27faf9f9cdf9b1f98df976f971f966f95bf958f950f94df94bf9;
    decBuf[2385] = 256'h3cf932f925f90df9fcf8e6f8ccf8b3f8aaf896f889f88bf88df89bf8aef8c6f8;
    decBuf[2386] = 256'he8f812f92ef95cf988f9a4f9c8f9f2f903fa26fa47fa5cfa77fa97fab4fad7fa;
    decBuf[2387] = 256'h01fb28fb56fb8ffbc3fb01fc3bfc7efcbefc08fd3afd7afdb4fddafdfcfd1bfe;
    decBuf[2388] = 256'h2cfe3bfe49fe56fe5afe6bfe7bfe89fea6febafed2feeefe02ff1aff2aff2dff;
    decBuf[2389] = 256'h2aff28ff19ff03ffeffed2feb7fe97fe79fe5efe46fe2afe0ffefdfde7fdd3fd;
    decBuf[2390] = 256'hc6fdb1fd9cfd8ffd7afd66fd4efd32fd17fdfefce2fccffcb6fca7fc9efc91fc;
    decBuf[2391] = 256'h8ffc95fc97fcaafcc2fcd8fcf7fc15fd38fd58fd7ffd98fdb9fdd6fdeafdfbfd;
    decBuf[2392] = 256'h0bfe1ffe37fe59fe79feb1fee5fe23ff6dffb3ff050052009800d80012013801;
    decBuf[2393] = 256'h5a0179018a01a401b201c701e201fa011d023d025b028602ad02d102f1020f03;
    decBuf[2394] = 256'h2a0343035203610368036b0364035e03520340032b031703ff02e902d502c802;
    decBuf[2395] = 256'hc102b202b402b902bb02bf02c602c502c602bf02b202a00286026d0251023e02;
    decBuf[2396] = 256'h1e0212020602fc0105020e0220023f025d0278029702b502c802e102f002f302;
    decBuf[2397] = 256'h0003030301030b031703220339035b037c03a203d003fc032e046c049504ca04;
    decBuf[2398] = 256'hfa0426054d0571059105af05c305cd05dd05eb05f305ff0512061f0639065906;
    decBuf[2399] = 256'h7606a906cb06f7062a074c076b078707a107a607aa07a6078d07840770075807;
    decBuf[2400] = 256'h4907400733073a073c073e0751075f076a0779078307820786077c0767075f07;
    decBuf[2401] = 256'h470725070e07f806dd06cc06c206b406b706b906bb06c906d206d306e406f306;
    decBuf[2402] = 256'hf106f606fb06f906fe06fa06ed06f206f406ed06f80600070407170733074707;
    decBuf[2403] = 256'h6d079107b207d807060819084008640869088608920895089f08a708aa08bb08;
    decBuf[2404] = 256'hce08db08ff082209430969098d09ad09d409f709050a230a2f0a2b0a350a320a;
    decBuf[2405] = 256'h250a270a210a170a180a170a0f0a1e0a280a2e0a430a510a590a6e0a770a740a;
    decBuf[2406] = 256'h7b0a790a670a600a510a370a2d0a170a030afb09f409e509ef09f409f309030a;
    decBuf[2407] = 256'h120a140a240a2e0a2c0a3c0a3e0a300a350a310a230a250a1d0a0c0a130a190a;
    decBuf[2408] = 256'h130a220a340a3b0a570a6a0a7c0a980aa30aa70abd0ac00ab80abf0abd0ab30a;
    decBuf[2409] = 256'hb40ab30aab0aba0ac40aca0ae20a020b0e0b390b550b640b850b9a0ba60bb70b;
    decBuf[2410] = 256'hc10bb80bc00bb90bae0bb00bb20ba60bb70bc60bcc0be30bff0b0a0c2a0c480c;
    decBuf[2411] = 256'h530c730c880c8c0ca40ca70c9f0cac0caa0c960c940c880c750c6d0c610c4a0c;
    decBuf[2412] = 256'h4d0c4a0c420c4e0c500c4a0c5a0c5c0c4e0c500c410c230c0e0cf30bbe0ba80b;
    decBuf[2413] = 256'h850b4d0b370b220bf60af10ae10aca0ac60aba0a9b0a960a830a5d0a4d0a360a;
    decBuf[2414] = 256'h070ae809cc09a80991097c0959094b093e092b092e092b092309300932093009;
    decBuf[2415] = 256'h420944093e0948094a0942094c094b093f09440945093f094509480949095609;
    decBuf[2416] = 256'h64096c098509a409b109d409eb09f8090b0a160a130a150a0e0af809f009dd09;
    decBuf[2417] = 256'hc309b909af09a109a309a6099f09a909a40996099409840964094d092f090409;
    decBuf[2418] = 256'he808ba0882085c082c080108d907ab077f0763073507fd06e606b6068a066e06;
    decBuf[2419] = 256'h40062106fa05d605ac059005620536050f05e104b5048d046a0440042f041504;
    decBuf[2420] = 256'hfe03f203e603db03df03dc03d403d603d003be03b703ac039e03950390038c03;
    decBuf[2421] = 256'h90039903a503ba03d403ed0309041c042e0444045204550460045a0458045a04;
    decBuf[2422] = 256'h55044d044f044b0441043d0434042804230415040604fb03e903d803c103ab03;
    decBuf[2423] = 256'h9103790350032903fb02c2027f023f02f501af016f012501df009f0054000e00;
    decBuf[2424] = 256'he1ffa7ff64ff36ffecfebafe68fe31fed7fd9afd4dfd07fdb5fc68fc22fcf4fb;
    decBuf[2425] = 256'hbafb86fb56fb2afb0efbeafacafaacfa91fa78fa5cfa49fa30fa1afa06faf4f9;
    decBuf[2426] = 256'he8f9e2f9dcf9ddf9dff9e1f9eaf9f5f906fa19fa2bfa3cfa5cfa73fa80fa9bfa;
    decBuf[2427] = 256'hacfabcfad0fad8fadffaeafaecfae7faebfae4fae3fae9fae5fae4faecfaebfa;
    decBuf[2428] = 256'he8faedfadffad1fac9fab0fa8afa70fa3dfa0dfae1f9a4f96af944f906f9cdf8;
    decBuf[2429] = 256'ha7f869f830f80af8daf7a2f77cf73ef705f7dff6a1f667f633f6f5f5abf579f5;
    decBuf[2430] = 256'h39f5fff4daf49cf473f44df41df4fef3edf3d3f3bcf3b8f3a4f39af39df394f3;
    decBuf[2431] = 256'h8df398f38ef38cf398f393f395f3a9f3acf3b4f3d3f3e0f3fbf321f445f466f4;
    decBuf[2432] = 256'h94f4b4f4d0f4fef411f52df546f554f569f585f588f598f5acf5b4f5c4f5e0f5;
    decBuf[2433] = 256'he4f5f5f50bf608f610f621f616f60cf611f6f9f5daf5c4f5a1f578f55cf523f5;
    decBuf[2434] = 256'heff4daf4a2f46df44bf413f4edf3cbf39ff36df34af31ef3ecf2c9f291f25df2;
    decBuf[2435] = 256'h2df2f4f1c0f190f157f123f1f3f0c7f094f080f054f038f033f01cf00ff013f0;
    decBuf[2436] = 256'h08f0ffef08f005f007f012f010f015f024f026f036f051f05df075f09ef0baf0;
    decBuf[2437] = 256'hdef01af143f169f1a7f1d0f1f5f133f25df282f2b2f2d1f2f9f227f33af361f3;
    decBuf[2438] = 256'h99f3b0f3d2f30bf421f443f47cf492f4a7f4dff4e7f4fbf41af520f525f53cf5;
    decBuf[2439] = 256'h38f534f538f528f525f523f50df505f507f5f2f4e9f4ecf4e0f4d5f4d7f4c8f4;
    decBuf[2440] = 256'hc1f4bff4a8f493f48af46df45af44ff433f420f415f4fff3fcf304f4fdf308f4;
    decBuf[2441] = 256'h1ef421f433f44df45ff475f48ef4a0f4b6f4d5f4ebf406f52cf546f570f597f5;
    decBuf[2442] = 256'hbbf5eef51ef64af687f6c1f6f6f634f76df7a2f7edf733f861f89bf8def80cf9;
    decBuf[2443] = 256'h46f97af9aaf9d6f914fa3dfa63faa1facafaeffa1ffb4bfb73fb96fbb7fbd5fb;
    decBuf[2444] = 256'hf7fb05fc12fc25fc29fc2cfc35fc32fc39fc40fc3efc3ffc44fc43fc47fc50fc;
    decBuf[2445] = 256'h4cfc4bfc4afc42fc3dfc34fc26fc1dfc12fcfefbf7fbebfbdcfbd2fbcdfbc8fb;
    decBuf[2446] = 256'hc9fbcdfbd1fbdbfbedfbf9fb10fc26fc35fc51fc6dfc85fc9bfcb5fccdfce9fc;
    decBuf[2447] = 256'h05fd24fd42fd65fd85fdb4fde0fd07fe3ffe74fea4fedcfe11ff41ff79ffaeff;
    decBuf[2448] = 256'hdeff090031005f008b00b200d600000127014b017e01a001cc01f30121024102;
    decBuf[2449] = 256'h68028c02ac02ca02dd02f6020c031a032c033d0348035603650370037a038603;
    decBuf[2450] = 256'h8e039903a803b203be03cd03db03e403ef03f703fd030604030406040c040804;
    decBuf[2451] = 256'h07040d040f041604210429043d0454046404780490049f04b904cb04da04ee04;
    decBuf[2452] = 256'h010508051f052f053d05550571057d059505b705cf05ec050f0626064d067006;
    decBuf[2453] = 256'h9106b706db06f20618073c07530771078c079e07b407c807d507ea07fe070608;
    decBuf[2454] = 256'h2008320841085b086d087c089108a308aa08b908c308c108cd08ce08c708d008;
    decBuf[2455] = 256'hd308cc08d408d808d108d508d408c908ca08c608b408ad08a208900889087a08;
    decBuf[2456] = 256'h6c0867085c084e0849084108330835082d082208260820081608220824081d08;
    decBuf[2457] = 256'h2c0836083708460850084b0859085f085e0866086d0869087708800881089508;
    decBuf[2458] = 256'ha208ae08c508db08e408fb080b0914092609320938094a095b095d096f097b09;
    decBuf[2459] = 256'h7d098f099b099909a309a8099d09a409a009920994098f097f097c0976096709;
    decBuf[2460] = 256'h65095f094f0948093e0928091e091609fe08ee08e008c808bf08b6089f089c08;
    decBuf[2461] = 256'h8d087b086f0864084e0846083308230818080a08f707f407e807de07e007db07;
    decBuf[2462] = 256'hcf07d407d007c407c907c507b707c007be07b707c307c807c607d507df07de07;
    decBuf[2463] = 256'hf007f707f907070809080708110810080708110813080f08150814080e081208;
    decBuf[2464] = 256'h0e080008fe07f607e707e107d507c307c107b207a0079d07930781077a076607;
    decBuf[2465] = 256'h4f07450737071a07ff06e706ca06af0697066e06520638060f06f305cf05a505;
    decBuf[2466] = 256'h89056505450527050c05e504cc04b50497048b0473045d044f043c042c041d04;
    decBuf[2467] = 256'h0b04f503e703da03c403bc03a90399038e03840374037203680360035e035903;
    decBuf[2468] = 256'h5303560353035003560359035a03610367036c037703800384038b038f039203;
    decBuf[2469] = 256'h9b039f03a003a503a2039c039b0395038a037e03710361034e033c0322031003;
    decBuf[2470] = 256'hf402d902c702b102980286026a024f0236021a02ff01e001c2019f017f015001;
    decBuf[2471] = 256'h2401fd00cf00a3007b004d002200faffccffa0ff79ff55ff2bff04ffe0fec0fe;
    decBuf[2472] = 256'ha2fe7ffe68fe4afe2ffe17fe07feedfddcfdccfdbefdb6fdaffda4fda6fda8fd;
    decBuf[2473] = 256'ha6fdabfdb4fdbbfdc2fdc9fdd0fdd7fde2fde6fde9fdeffdf4fdfcfd04fe0ffe;
    decBuf[2474] = 256'h1cfe25fe30fe41fe4cfe56fe65fe70fe7afe8afe90fe92fe9bfe9cfe9bfe9cfe;
    decBuf[2475] = 256'h96fe8efe87fe7afe64fe56fe39fe1efe05fee9fdc6fdaffd89fd65fd4efd28fd;
    decBuf[2476] = 256'hf9fcdafcb3fc8ffc65fc3efc10fce4fbbdfb8ffb6ffb48fb1afb07fbe0fac6fa;
    decBuf[2477] = 256'haffa91fa7efa65fa43fa2cfa0efaebf9d4f9bff9a4f992f983f96ef967f964f9;
    decBuf[2478] = 256'h62f960f969f971f97bf98bf995f9a8f9bff9d5f9eff90ffa24fa3ffa5ffa74fa;
    decBuf[2479] = 256'h8ffaaefabbfad6faeffaf8fa0cfb1ffb2ffb3efb54fb5dfb6ffb85fb87fb95fb;
    decBuf[2480] = 256'ha5fba7fbadfbb3fbaefbacfbb0fba8fba2fba5fb9afb8efb90fb81fb6ffb63fb;
    decBuf[2481] = 256'h4bfb2ffb1cfbf5fac7faa8fa81fa52fa27fafff9c7f9a1f971f946f91ef9f0f8;
    decBuf[2482] = 256'hc4f8a8f87af85bf83ff81bf8faf7eef7d3f7c1f7b1f79df78bf77ff76cf75af7;
    decBuf[2483] = 256'h4ef73bf72df726f71cf716f717f719f721f72df738f74cf763f773f787f7a4f7;
    decBuf[2484] = 256'hb7f7d0f7f2f709f827f852f879f89df8d0f8f2f82bf95ff981f9adf9e0f902fa;
    decBuf[2485] = 256'h21fa49fa6dfa84faa2fabdfad5faebfaf9fa0cfb1cfb27fb31fb3dfb3ffb43fb;
    decBuf[2486] = 256'h4afb47fb48fb4dfb45fb3ffb40fb37fb30fb29fb19fb08fbf9fadffac7fab1fa;
    decBuf[2487] = 256'h91fa73fa58fa39fa1bfa00fae0f9c3f9aff990f97af967f94ff939f92af918f9;
    decBuf[2488] = 256'h0cf90af900f9fef803f908f911f921f930f94af963f97ff99af9baf9d7f9faf9;
    decBuf[2489] = 256'h1bfa41fa65fa8efaaafacefaf8fa1ffb43fb6dfb94fbc2fbeefb15fc44fc7cfc;
    decBuf[2490] = 256'ha1fcd1fc0afd3efd6efda7fdccfdfcfd28fe44fe72fe91feaefebdfeddfeeafe;
    decBuf[2491] = 256'hf6fe00ff0aff0cff0fff0dff0bff05fff5feeafedcfec9feb7fea6fe8ffe79fe;
    decBuf[2492] = 256'h65fe52fe42fe2efe1cfe10fe01feeffddffdd4fdc2fdb1fd9efd8cfd80fd69fd;
    decBuf[2493] = 256'h53fd44fd32fd1dfd0efd01fdf5fcebfce1fcd8fcdafcd8fcdcfce5fceffcfefc;
    decBuf[2494] = 256'h14fd28fd45fd60fd80fd9efdc0fde1fd07fe2bfe4bfe72fe95febffedbfe09ff;
    decBuf[2495] = 256'h29ff45ff73ff92ffb9ffddfffeff1b00460062008600b000cc00f00010013601;
    decBuf[2496] = 256'h500170018e01b101d101ef011202320250026b0284029a02ae02bb02c702cd02;
    decBuf[2497] = 256'hd702d502d402d502ce02c802c202bb02b502af02ab02aa02a702a502a4029f02;
    decBuf[2498] = 256'h9d029f02a0029f02a402a602a602ad02b302b602be02c402c502cc02d202d302;
    decBuf[2499] = 256'hdd02e602e502ed02f802fc020603110319032b033b0346035c03700382039d03;
    decBuf[2500] = 256'hbc03d103f40315043204550476049304b604d704f4040f05280538054c055e05;
    decBuf[2501] = 256'h6a0575057b0583058b058d058e05900593059205910592058f058e058c058705;
    decBuf[2502] = 256'h8705820580057f05790571056b05620557054c053d052b051b050305e704d404;
    decBuf[2503] = 256'hbb049f048c046c0457043c0423040104ea03d503b903a80392037e0371036503;
    decBuf[2504] = 256'h5a0358035703550359035b0357035f0360035a035b0355034b0347033e033203;
    decBuf[2505] = 256'h2d0325031c031d031a0315031703180315031a031c031d0327032e032f033903;
    decBuf[2506] = 256'h46034a035b03660370037f038a039403a003ac03ad03b903c203c303c703cd03;
    decBuf[2507] = 256'hcc03d303d403d203d803d903d403d903dd03de03e603ee03f303000412041e04;
    decBuf[2508] = 256'h35044b045f0477048c049b04b804cb04d604eb04fa0402050e0518051e052705;
    decBuf[2509] = 256'h2f05310537053b053c0547054f0553055c05680570057e058a059205a305ad05;
    decBuf[2510] = 256'hb305bf05c805cc05d605d905db05e205e205e005e205e205db05db05d305c405;
    decBuf[2511] = 256'hba05aa05970585056b055205430529051005fa04e604d404c804b904ab04a204;
    decBuf[2512] = 256'h970489048404760468045b044d043b042a041304fd03e903d103b5039a037a03;
    decBuf[2513] = 256'h5d03410322030403f102d102b402a0028f027902650258024702380226021a02;
    decBuf[2514] = 256'h1002fe01f201e701d901cd01c101b401a4019a018801770164014c0136012201;
    decBuf[2515] = 256'h0b01ee00d300bb009f0084006b005500410029001a000600f3ffe3ffd4ffc6ff;
    decBuf[2516] = 256'hbaffaeffa1ff94ff89ff79ff6aff5cff45ff2fff1bfffefee3fec3fea6fe83fe;
    decBuf[2517] = 256'h6cfe4efe33fe1afe0bfef7fde9fdd9fdcafdc4fdb8fdb0fda8fd9efd98fd95fd;
    decBuf[2518] = 256'h94fd91fd96fd9cfda2fdadfdb9fdc3fdcffdd8fde2fdecfdf4fdfafd03fe0cfe;
    decBuf[2519] = 256'h16fe20fe2dfe3dfe50fe63fe78fe92feb1fecffeeafe0aff30ff54ff74ff9aff;
    decBuf[2520] = 256'hbeffe8ff0f0033005d008400a800c800de00f900110121012f0142014e015801;
    decBuf[2521] = 256'h620172017d01870193019b01a501af01b301b801bb01bb01ba01b901b401ae01;
    decBuf[2522] = 256'hac01a6019f0198019001830176016801560140012c010f01f400dc00c0009d00;
    decBuf[2523] = 256'h7c005f00440024000600ebffccffaeff93ff7aff64ff56ff44ff38ff29ff23ff;
    decBuf[2524] = 256'h1aff15ff0bff01fff8feeafedcfec9feb6fea1fe8dfe75fe65fe51fe3ffe2efe;
    decBuf[2525] = 256'h1ffe11fe05fefafdeffde0fdd2fdc6fdb7fda9fd9afd8bfd81fd74fd66fd60fd;
    decBuf[2526] = 256'h54fd42fd3bfd2cfd16fd02fdeafccefcb3fc93fc6dfc53fc2afc02fce9fbbffb;
    decBuf[2527] = 256'h98fb74fb4afb23fbf5fac9faa2fa7efa54fa2dfa09fae8f9c2f9a9f991f974f9;
    decBuf[2528] = 256'h60f948f92cf918f9f9f8dbf8c0f8a0f883f868f848f82af80ff8f7f7e7f7d9f7;
    decBuf[2529] = 256'hc6f7bff7bdf7b7f7b9f7bef7bff7c9f7d7f7e3f7f8f712f82af846f869f88af8;
    decBuf[2530] = 256'hb0f8d4f8fdf825f953f97ff9b1f9e1f90dfa4bfa74faa9fae7fa20fb55fb93fb;
    decBuf[2531] = 256'hcdfb01fc4dfc7ffcbffcf8fc3cfd7cfdc6fd0cfe4cfe96fedcfe1cff66ffacff;
    decBuf[2532] = 256'hecff26005a008a00c300f7001a0145016d019101ba01d601f001100226024102;
    decBuf[2533] = 256'h52026802760289029502a402b202be02c602d302dc02e802ef02f602fa02fd02;
    decBuf[2534] = 256'hfa02f902f702ed02e602dd02d102c902be02b202a7029c029002840277026402;
    decBuf[2535] = 256'h560246023702290219020a020002f801ef01e801e401e001dd01d801d201ca01;
    decBuf[2536] = 256'hc001b301a5018f017a01630147012c010c01ee00cb00ab008500610037001000;
    decBuf[2537] = 256'hecffb9ff89ff5dff36fffefec9fe99fe61fe2cfeeefdb5fd80fd42fd08fdc5fc;
    decBuf[2538] = 256'h85fc3bfc09fcb7fb6afb38fbe6fa99fa53fa13fac8f982f930f9f9f8b3f873f8;
    decBuf[2539] = 256'h29f8f7f7b7f77ef749f719f7edf6c6f698f678f65cf643f62cf61ff60bf601f6;
    decBuf[2540] = 256'hfef5f5f5f3f5f5f5f3f5fdf509f60ef621f639f649f668f68ff6b2f6dcf60ff7;
    decBuf[2541] = 256'h3ff777f7bbf7faf745f88bf8cbf825f97af9c7f921fa76fad9fa37fb8cfbeffb;
    decBuf[2542] = 256'h4cfcb9fc03fd7bfdcdfd34fe92fefffe66ffc4ff31007a00f3004401ab010902;
    decBuf[2543] = 256'h5e02c1021e037303d60334048904d60444058e05eb0540067706d1060e075b07;
    decBuf[2544] = 256'h8d07df071608480875089f08d308f60815093c09600977099509b009c209de09;
    decBuf[2545] = 256'hf109fc090b0a1a0a210a2d0a380a3a0a430a480a430a440a3e0a300a2a0a160a;
    decBuf[2546] = 256'hff09ef09cf09b209970970094c092c09fd08d108aa087c0850081d08ed07b507;
    decBuf[2547] = 256'h72073207f806b40675062a06e40592054505ff04ad0460040604b10364030a03;
    decBuf[2548] = 256'h9d023602d8016b010401a6003900b4ff5bffe9fe82fe0afe98fd31fdb8fc46fc;
    decBuf[2549] = 256'hdffb82fb14fbadfa50fae2f97bf91ef9b0f867f809f89cf752f7f5f6a0f653f6;
    decBuf[2550] = 256'h0df6bbf56ef528f5e8f4aef46af43df414f4dff3bdf39df381f368f35af34df3;
    decBuf[2551] = 256'h41f33ef33bf343f351f35cf378f393f3acf3d4f307f429f462f496f4d4f40ef5;
    decBuf[2552] = 256'h51f591f5ecf528f675f6cff63df786f7e4f751f8b8f816f983f9eaf97dfae0fa;
    decBuf[2553] = 256'h5dfbeffb78fcf5fc88fd11fe8efe20ffaaff4b00e2006b01e9017b0204038103;
    decBuf[2554] = 256'h3404ab044205cc054906db0664070508710822099909300ab90a130ba50b070c;
    decBuf[2555] = 256'h840cf60c5d0dd60d270eac0e050f560fbe0f00105510a210d41014115e117c11;
    decBuf[2556] = 256'haa11d311ea11fe11111217122612221215120912f811d511be118f1164113111;
    decBuf[2557] = 256'hf310b91085103910df0fa30f560fe80e9e0e260eb40d4d0dd40c620cde0b610b;
    decBuf[2558] = 256'hce0a450ac8093609ac080b087407eb064a06b20529058804f1036703c6022f02;
    decBuf[2559] = 256'ha60105016d00e4ff43ffacfe22fe82fdeafc88fce7fb50fbeefa4dfae1f957f9;
    decBuf[2560] = 256'hdaf868f8e4f767f7f5f68ef615f6c4f55df5e4f493f42cf4e9f394f347f301f3;
    decBuf[2561] = 256'hd3f289f257f22af200f2ccf1a9f18af163f149f132f114f109f1f7f0e8f0eaf0;
    decBuf[2562] = 256'he3f0e5f0f8f000f115f135f153f176f1a8f1cbf103f238f275f2c0f206f346f3;
    decBuf[2563] = 256'ha0f3f5f342f4b0f417f575f5e2f549f6c2f654f7b6f733f8c6f84ff9f0f987fa;
    decBuf[2564] = 256'h11fbb1fb49fcd2fc73fd36feb8fe5fff2100d8007e011602c6029c032c04e304;
    decBuf[2565] = 256'hb80582063907df07a1085809ff09c10a440bea0bad0c2f0dd60d6d0ef60e730f;
    decBuf[2566] = 256'h06108f100c119e1101127e12ef123913b21303144d148f14cc14ed141f153a15;
    decBuf[2567] = 256'h4315591560155a155f1546152f151115e614b41484143f14ed13a0134613f112;
    decBuf[2568] = 256'h8e121512a4111f11a2101010860fe50e4e0ec50d240d8c0c030c3e0b870a110a;
    decBuf[2569] = 256'h4e09970820085e07a70601066905b904120450039902f3013001ad00070045ff;
    decBuf[2570] = 256'hc2fe1cfe84fdfbfc5afcc3fb39fbbcfa4afac6f949f9d7f870f8f7f785f71ef7;
    decBuf[2571] = 256'hc1f653f6ecf5a9f53cf5f2f4b0f45bf424f4def39ef375f331f303f3daf2a6f2;
    decBuf[2572] = 256'h76f24af222f2f4f1d5f1b9f195f17ef169f155f152f148f14bf153f15af165f1;
    decBuf[2573] = 256'h7bf189f19cf1bbf1d0f1ebf10af228f24bf275f29cf2caf202f337f375f3bff3;
    decBuf[2574] = 256'h05f445f4a0f4f5f458f5b5f50af66df6e5f637f7bbf739f8aaf812f98af91cfa;
    decBuf[2575] = 256'ha6fa23fbb5fb3efcbbfc4efdfefd75fe0cffbdff3400f60079011f02b7026703;
    decBuf[2576] = 256'hde03750426059d053406e5065c07f3077c08f9088c09150a920a240bae0b070c;
    decBuf[2577] = 256'h790cfe0c570dc90d130e700ead0efa0e2c0f6c0f950fc90fec0f0b101c103610;
    decBuf[2578] = 256'h43104810531050104010381025100210e80fb50f850f4d0f090fb70e800e260e;
    decBuf[2579] = 256'hd10d840d160dcc0c6f0c020c7d0b240bb20a2d0ad4094109b8085f08cc074307;
    decBuf[2580] = 256'hc60613069c0505057c04ff036c03e3024202d6014d01cf003d00b4ff37ffc5fe;
    decBuf[2581] = 256'h40fec3fd31fda7fc2afcb9fb34fbdafa48fae6f969f9f7f890f832f8c5f75ef7;
    decBuf[2582] = 256'h00f7abf648f6ebf596f549f503f5b1f44ef40bf4cef381f33bf3fbf2b1f27ff2;
    decBuf[2583] = 256'h52f218f2e3f1b3f187f16bf147f127f11af1fff0e7f0d7f0c3f0b6f0aff0a0f0;
    decBuf[2584] = 256'h96f098f093f094f0a3f0a9f0bdf0dff0f6f014f146f168f194f1d2f1fbf13ff2;
    decBuf[2585] = 256'h7ff2b8f2fcf23cf375f3c8f315f45bf4adf4faf440f5a4f502f66ff6d6f634f7;
    decBuf[2586] = 256'ha1f708f881f8f3f85af9d2f944fac9fa22fb94fb19fc96fce7fc6cfde9fd5bfe;
    decBuf[2587] = 256'hc2fe3affacff3100ae0020018701ff017102d8023603a3030a046804bd042005;
    decBuf[2588] = 256'h7d05d2051f067906ce061b076107a107eb0731087108bb08ed082d0967098c09;
    decBuf[2589] = 256'hbd09e809040a280a490a5e0a6a0a7b0a7e0a870a8f0a8c0a8a0a880a7f0a770a;
    decBuf[2590] = 256'h6a0a5a0a4b0a310a190afd09d209ab097c0944091009e0089b085b081108cb07;
    decBuf[2591] = 256'h8b074107e706aa065d060306ae054b05ed0499043604bd036c0305038c021b02;
    decBuf[2592] = 256'hb3012001be004100cfff68fff0fe7efef9fd7cfd0afda3fc2bfcb9fb52fbd9fa;
    decBuf[2593] = 256'h67fae3f989f9f7f895f818f8a6f75cf7e4f672f628f6cbf55ef514f5b6f461f4;
    decBuf[2594] = 256'h2af4d0f394f35df317f3d7f29df269f239f20df2daf1b8f199f171f158f14af1;
    decBuf[2595] = 256'h3df131f12ef12bf12ef13bf142f151f16bf17cf192f1b7f1d1f1f1f118f23cf2;
    decBuf[2596] = 256'h65f298f2baf2f2f227f365f39ff3e2f322f46cf4b2f4f2f43cf596f5d3f536f6;
    decBuf[2597] = 256'h79f6cef61bf775f7b1f714f857f8acf80ff952f9a7f90afa67fabcfa1ffb7dfb;
    decBuf[2598] = 256'hd2fb35fc92fce7fc34fd8efde3fd46fea4fee0fe43ffa1fff6ff43009d00f200;
    decBuf[2599] = 256'h5501b20107026a02c8021d038003c30330047a04d7042c057905bf0511065e06;
    decBuf[2600] = 256'ha406f60643077507c707fe0744088408cf08010940097a09af09df090b0a320a;
    decBuf[2601] = 256'h600a7f0a9b0ab50acc0ae10aed0af80afb0a030b010bfe0af80aea0ada0acb0a;
    decBuf[2602] = 256'hb10a990a7d0a520a1f0afd09b8098b094009fa08bb0870081608c10774071a07;
    decBuf[2603] = 256'hc60679060b06c1056305f6048f043104c4033f03e6027402ef0196010401a200;
    decBuf[2604] = 256'h2500b3ff4cffd3fe61fefafd82fd10fda9fc4bfcdefb94fb37fbcafa80fa22fa;
    decBuf[2605] = 256'hcdf980f926f9eaf89df857f817f8ddf7a9f778f74df725f701f7e1f6ccf6b1f6;
    decBuf[2606] = 256'ha6f697f688f686f67ef681f687f68cf694f6a4f6aff6c9f6e2f6fef621f741f7;
    decBuf[2607] = 256'h67f795f7cef7f3f731f86bf89ff8ddf817f94bf997f9c9f909fa53fa99fac7fa;
    decBuf[2608] = 256'h11fb57fb97fbd1fb14fc54fc9efce4fc36fd83fdc9fd1bfe68fec2fe17ff64ff;
    decBuf[2609] = 256'haafffcff49008f00e2002f017501c70114025a02ac020f035203a703f4033a04;
    decBuf[2610] = 256'h8c04d9041f057105be05040644069e06db0628076e07ae07e8073a087108b708;
    decBuf[2611] = 256'hf70841098709c709010a440a840aae0af10a1f0b480b7c0bad0bcc0bf30b170c;
    decBuf[2612] = 256'h2e0c4c0c5f0c710c870c950ca20cae0cb90cbb0cc30cc20cba0cb60ca80c950c;
    decBuf[2613] = 256'h880c6e0c4e0c310c060cdf0bb10b780b440b140bcf0a8f0a550a030ab6098409;
    decBuf[2614] = 256'h1f09dd0888082508c70772070f07b2064406dd05650514058f043504c4035c03;
    decBuf[2615] = 256'hff0292022a02cd017801ff00ae004600e9ff7cff32ffd4fe67fe1dfec0fd6bfd;
    decBuf[2616] = 256'h08fdc5fc70fc23fcf1fbb1fb78fb43fb05fbdcfab6fa94fa81fa65fa4cfa3efa;
    decBuf[2617] = 256'h31fa25fa22fa1ffa1cfa24fa2bfa35fa43fa5afa70fa8afaa9fad0fae9fa1cfb;
    decBuf[2618] = 256'h3ffb6afb9dfbcdfbf9fb37fc60fca3fcd1fc0bfd4efd8efdc8fd0bfe5efe95fe;
    decBuf[2619] = 256'hdbfe2dff64ffaafffcff49008f00e10018015e019e01d8011b025b029502c902;
    decBuf[2620] = 256'h070330036503a303cc0300043e0468049c04da040305380576059f05c405f405;
    decBuf[2621] = 256'h200648066b068c06aa06cc06e4060a0723073b07580773078c07a207bc07cd07;
    decBuf[2622] = 256'he307f7070408150824082a083a084408460852085b085f0866086c086d087408;
    decBuf[2623] = 256'h7708730873087108670866085b084a083b0829080f08fe07db07bb079d077207;
    decBuf[2624] = 256'h4b072707fe06cb06a90670063c060c06e005a20579053505f504bc0478043804;
    decBuf[2625] = 256'hee03a80356030903af025a020d02b3015e01fb009e004900e6ff88ff33ffd0fe;
    decBuf[2626] = 256'h73fe1efebbfd5dfdf0fca6fc49fcdbfb92fb34fbdffa92fa38fafcf9aff969f9;
    decBuf[2627] = 256'h29f9eff8abf87ef844f810f8edf7c1f79af776f74df730f717f700f7f3f6e7f6;
    decBuf[2628] = 256'hd6f6d3f6d6f6ddf6eef601f719f735f760f787f7abf7def70ef846f87bf8b8f8;
    decBuf[2629] = 256'hf2f836f976f9c0f906fa46faa0faddfa2afb84fbd9fb26fc80fcd5fc22fd7cfd;
    decBuf[2630] = 256'hd1fd1efe78fecdfe1aff74ffc8ff15005b00ae00fb0055019101de0124026402;
    decBuf[2631] = 256'hae02f40234036e03a203d3030b043f0462048104b404c804e704040513052105;
    decBuf[2632] = 256'h36054905540564056c057405800582058c05910593058e058a0584057a056e05;
    decBuf[2633] = 256'h5f0551053e0521050d05ee04d004b504960478045d0436041204f203cc03a803;
    decBuf[2634] = 256'h87036a033f031803f402ca02a3027f0255022e020002d401ad017f0153012b01;
    decBuf[2635] = 256'hfd00d2009f006f0043001000d3ff99ff64ff34ffeffec2fe78fe46fe06febbfd;
    decBuf[2636] = 256'h75fd36fdfcfcb8fc78fc3ffcfbfbbbfb82fb4dfb0ffbc5fa93fa53fa09fad7f9;
    decBuf[2637] = 256'h85f94ef908f9c8f87ef84cf80cf8c1f78ff750f716f7e1f6a3f67af646f616f6;
    decBuf[2638] = 256'heaf5cef5aaf589f56cf551f538f528f50ff504f5fbf4f2f4eff4f2f4f0f4faf4;
    decBuf[2639] = 256'h09f514f526f540f552f56ef591f5b1f5d7f505f631f664f694f6ccf601f73ff7;
    decBuf[2640] = 256'h89f7cff70ff859f8b3f808f955f99bf9fff95dfab2fa15fb58fbc5fb2cfc6ffc;
    decBuf[2641] = 256'hdcfc26fd83fdd8fd3bfe7efeebfe35ff78ffcdff1a007400b000fd0043019501;
    decBuf[2642] = 256'hcc01120252028c02c102fe0238035e038e03ad03d403ee030e04240437044904;
    decBuf[2643] = 256'h52045b04620465046304610454044604380425040d04f703dd03be03a0037d03;
    decBuf[2644] = 256'h5d0336031303e902c2029e02740241021f02e701c1019101650133010301d700;
    decBuf[2645] = 256'h990070003b000b00d3ff9eff6eff43ff10ffe0feb4fe81fe51fe26fefefddafd;
    decBuf[2646] = 256'hb1fd89fd70fd46fd1ffd05fde5fcc7fcacfc8cfc6ffc53fc34fc16fcfbfbe3fb;
    decBuf[2647] = 256'hc6fbb3fb9bfb7efb6bfb4cfb36fb23fb0afbf5fae0fac9fab3faa5fa8dfa77fa;
    decBuf[2648] = 256'h69fa56fa41fa33fa25fa10fa07fafaf9e5f9dcf9cff9bff9b4f9aaf99af990f9;
    decBuf[2649] = 256'h82f975f96df960f953f94ff947f940f93cf939f93af93df93ef944f94ff957f9;
    decBuf[2650] = 256'h62f976f985f997f9acf9c1f9d8f9f4f908fa27fa45fa68fa88faaefad2faf3fa;
    decBuf[2651] = 256'h21fb4dfb75fbadfbe1fb12fc3dfc70fcaefce8fc1cfd5afd94fdc8fd14fe46fe;
    decBuf[2652] = 256'h86fed0fe16ff44ff8effd4ff01004c009200bf000a013c017b01b501f9012602;
    decBuf[2653] = 256'h60029502c502f0022303450371039903bc03dd03030427043e045c0477048804;
    decBuf[2654] = 256'h9e04b204c004cb04d204dc04e104e304de04d704d404c704b904af04a2048d04;
    decBuf[2655] = 256'h79046704510437041f040304ef03d003b203970378035a033f031803f402dd02;
    decBuf[2656] = 256'hb70293027c0256023c021c02fe01e301c301ae018b017d016001440133011d01;
    decBuf[2657] = 256'h0301f200e200ce00bc00b000a100930087007b0074006d006700630060005f00;
    decBuf[2658] = 256'h6200650065006a006c0073007c00830089008f0094009c00a800b000b800c100;
    decBuf[2659] = 256'hca00d400e100ec00fa00060111011f012701330140014d0155015f0169016f01;
    decBuf[2660] = 256'h75017c01840189018c019101970199019c019f019f01a001a301a601a501a001;
    decBuf[2661] = 256'h9e019901970192018c0184017f0176016d0167015e01560150014b0143013b01;
    decBuf[2662] = 256'h36012e012b01260122011f011901130112010f010b0108010701050106010a01;
    decBuf[2663] = 256'h0b010a010e0116011e0125012b013501410149015701670171017f018b019a01;
    decBuf[2664] = 256'hac01bd01cc01de01ee01fd0117022902380252026b0280029a02b302c202dc02;
    decBuf[2665] = 256'hf5021103240336034c036603770387039b03b203c203d003e303f30302041404;
    decBuf[2666] = 256'h2004330440044c045b0465046a047904830485049004950496049c04a204a104;
    decBuf[2667] = 256'ha404a604a504aa04a904a404a704a804a404a804a7049f049e049b0497049804;
    decBuf[2668] = 256'h93048b048f048e0488048c048d0488048f04960498049f04a504a704b404c204;
    decBuf[2669] = 256'hc404d304e504e704f60400050905170525052b053d054d055405660576058105;
    decBuf[2670] = 256'h9305a305ae05c005cc05db05ed05f405fa050806150616061e0622061e062106;
    decBuf[2671] = 256'h20061e061d0613060406fa05ee05d905ca05b80599058405610541052305f804;
    decBuf[2672] = 256'hd104ad047a044a041e04ec03ae03850350031203d802950267021d02eb01ab01;
    decBuf[2673] = 256'h61011b01db00a1004f001800d2ff80ff49ff03ffb1fe7afe34fef4fdbafd85fd;
    decBuf[2674] = 256'h48fd0efdd9fca9fc7dfc4bfc28fcfdfbd5fbb1fb9afb7dfb61fb50fb47fb32fb;
    decBuf[2675] = 256'h25fb1efb1cfb1efb20fb28fb32fb3ffb51fb66fb7afb92fbaefbd1fbf1fb0ffc;
    decBuf[2676] = 256'h3afc61fc85fcb8fce8fc14fd51fd8bfdc0fdf0fd35fe74feaefef2fe32ff6bff;
    decBuf[2677] = 256'hafffefff28005d009b00d500180146017f01b401f2011b0250028002b802ec02;
    decBuf[2678] = 256'h0f033b036d039d03bd03ef0312043104580472048904a704ca04e104ed040905;
    decBuf[2679] = 256'h1a052a0538054505510560056a05730578058205860585058805870585058605;
    decBuf[2680] = 256'h85057f057e05780571056f056a05640563055a0550054f0547053c0535052505;
    decBuf[2681] = 256'h17050f05f604e504d504bb04a3048d046d04500434041504ef03d503ab038403;
    decBuf[2682] = 256'h6a0338031503e902b70287025b022802f801c0017c013d010301bf007f003500;
    decBuf[2683] = 256'hefff9dff50fff6feb9fe6cfe12febefd5bfdfdfcc0fc5dfc00fcabfb5efbf0fa;
    decBuf[2684] = 256'ha6fa48faf4f991f94ef9e1f897f854f8fff7b2f76cf72cf7e2f6b0f65ef627f6;
    decBuf[2685] = 256'hf5f5c7f58df559f537f517f5f0f4ccf4bef4a0f495f48af487f48af492f49ef4;
    decBuf[2686] = 256'hadf4cbf4e8f40bf535f55cf58af5c3f5f7f535f67ff6c5f605f760f79df700f8;
    decBuf[2687] = 256'h5df8b2f8fff86df9d4f932fa9ffa06fb64fbd1fb38fcb1fc22fd6cfde5fd56fe;
    decBuf[2688] = 256'hbefe36ff87ffeeff6700b8001f017d01ea0134029102e60233038d03e2031904;
    decBuf[2689] = 256'h5f049f04c8040c05390563058805ab05ca05e60500060d0623062e0632063506;
    decBuf[2690] = 256'h380635062e06230615060606f305db05b905a1057b0557052e050605d804a004;
    decBuf[2691] = 256'h7a043d040304dd039f0366032203e202a90274023602ec01ba017a013001fe00;
    decBuf[2692] = 256'hac0075002f00efffb5ff72ff32ffe7feb5fe63fe2cfefafda8fd71fd2bfdebfc;
    decBuf[2693] = 256'hb2fc6efc2efce4fb9efb5efb24fbe1faa1fa67fa24fae4f9aaf967f927f9edf8;
    decBuf[2694] = 256'hb8f86df83bf8fbf7d2f79df752f720f7f2f6a8f676f648f60ef6daf5aaf571f5;
    decBuf[2695] = 256'h3df51bf5eff4bcf49af46ef447f42df40df4eff3dcf3c3f3adf3a5f392f38bf3;
    decBuf[2696] = 256'h8df383f388f391f398f3aaf3bbf3c9f3e7f30ef427f451f478f4a6f4d2f410f5;
    decBuf[2697] = 256'h4af58df5cdf507f659f6a6f6ecf63ff7a2f7e4f752f8b9f816f984f9ebf948fa;
    decBuf[2698] = 256'hcefa27fb99fb1efc9bfcecfc71fdeefd60fec7fe3fffb1ff1800910002016a01;
    decBuf[2699] = 256'hc70134029c02f9024e03b1030f044b049804f2042f057c05c205f00529065e06;
    decBuf[2700] = 256'h8006ac06d306e306fa060f07230726072907260719070d07fa06e306c606a406;
    decBuf[2701] = 256'h7a0653062406ec05b8057a054005fd04bd0472042c04da038d033303de029102;
    decBuf[2702] = 256'h3702e30196013c01e70084002600d1ff6eff11ffbcfe59fefbfda6fd43fd00fd;
    decBuf[2703] = 256'habfc48fc06fcb1fb64fb0afbcdfa80fa3afafaf9c0f97df93df903f9def8aef8;
    decBuf[2704] = 256'h75f850f820f8f4f7cdf7a9f788f76bf748f731f71bf708f7f0f6e6f6d2f6c5f6;
    decBuf[2705] = 256'hbef6aff6a9f6abf6a3f6a1f6a8f6a4f6a8f6b5f6b6f6bef6d2f6dff6ebf6fef6;
    decBuf[2706] = 256'h10f726f73af74cf76bf789f79cf7bcf7daf7edf713f837f84ef875f8a3f8c2f8;
    decBuf[2707] = 256'he9f818f937f969f99af9c5f903fa2cfa61fa9ffad9fa0dfb4bfb85fbb9fb05fc;
    decBuf[2708] = 256'h37fc77fcc1fc07fd47fd91fdc3fd15fe62fea8fee8fe32ff78ffb8ff13005000;
    decBuf[2709] = 256'h9d00e30035016c01b20104023b029502d10208034e038e03d9030b044a048404;
    decBuf[2710] = 256'hc804f5042f0564058605be05e405060625064d06660687069c06af06c106d006;
    decBuf[2711] = 256'hdf06e706e906eb06ed06eb06e706df06d006c206b2069b0685066b064c062e06;
    decBuf[2712] = 256'h0b06e105ba059605630533050705e004a804730443040b04d60398035f033903;
    decBuf[2713] = 256'hfb02c1028d024f021502e101b101780144010601dd00a800780040001a00eaff;
    decBuf[2714] = 256'hbfff97ff73ff4aff2eff0affe9fed4feb9fe99fe8dfe72fe60fe57fe48fe3bfe;
    decBuf[2715] = 256'h39fe37fe31fe36fe38fe39fe45fe54fe5efe6efe81fe8efea3febdfed6feecfe;
    decBuf[2716] = 256'h0bff21ff43ff64ff82ffa4ffceffeaff1800440060008400b700d90005013801;
    decBuf[2717] = 256'h5a018601b801db0107022e025c027b02ae02d002fc0223033d0367038e03a803;
    decBuf[2718] = 256'hc803e603010420043e045204710486049a04b204c804d604e904f90404051205;
    decBuf[2719] = 256'h1e05260531053d05420547054b054c054f0552055005520553054b054a054705;


    $display("Done initializing");

  end

  //---------------------------------------------------------------------------------------
  // test bench implementation
  // global signals generation
  always @(posedge clk) begin
    mCtr <= mCtr + 1;

    if (testCount >= TESTS_TO_RUN) $finish(1);

    case (mainState)
      MAIN0: begin
        rst <= 1;

        inDone <= 0;
        encDone <= 0;
        decDone <= 0;

        if (mCtr >= 2) begin
          $display("");
          $display("IMA ADPCM encoder & decoder simulation");
          $display("--------------------------------------");
          mCtr <= 0;
          mainState <= MAIN1;
        end
      end

      MAIN1: begin
        rst <= 0;

        mCtr <= 0;
        mainState <= MAIN2;
      end // case: MAIN1

      MAIN2: begin
        if (inDone && encDone && decDone) begin
          $display("Test %d done!. mCtr: %d", testCount , mCtr);

          testCount <= testCount + 1;
          mCtr <= 0;
          mainState <= MAIN0;
        end
      end

    endcase // case (mainState)
  end

  //------------------------------------------------------------------
  // encoder input samples read process
  always @(posedge clk) begin
    iCtr <= iCtr + 1;
    if (rst) inState <= IN1;

    case (inState)
      IN0: begin
        iCtr <= 0;
      end

      IN1: begin
        // clear encoder input signal
        inSamp <= 16'b0;
        inValid <= 1'b0;
        // clear samples counter
        sampCount <= 0;
        inBytesRead <= 0;

        // binary input file
        inIdx <= 0;

        if (!rst) begin
          iCtr <= 0;
          inState <= IN2;
        end
      end // case: IN1

      IN2: begin
        if (iCtr >= 50) begin
          // read input samples file
          intmp <= inBuf[inIdx][(BUFFER_BYTES << 3) - 1:(BUFFER_BYTES << 3) - 8];
          inBytesRead <= inBytesRead + 1;

          $display("inBuf[%d] = %h%h%h%h%h%h%h%h", inIdx,
                   inBuf[inIdx][255:224],
                   inBuf[inIdx][223:192],
                   inBuf[inIdx][191:160],
                   inBuf[inIdx][159:128],
                   inBuf[inIdx][127:96],
                   inBuf[inIdx][95:64],
                   inBuf[inIdx][63:32],
                   inBuf[inIdx][31:0]);


          iCtr <= 0;
          inState <= IN3;
        end
      end // case: IN2

      IN3: begin
        // Stop looping through inputs if eof
        if (inBytesRead >= TOTAL_IN_BYTES) begin
          $display("Reached eof of input");

          iCtr <= 0;
          inState <= IN5;
        end

        else begin
          if (iCtr == 0) begin
            // read the next character to form the new input sample
            // Note that first byte is used as the low byte of the sample
            inSamp[7:0] <= intmp;

            case (inBytesRead % BUFFER_BYTES)
              1:  inSamp[15:8] <= inBuf[inIdx][247:240];
              3:  inSamp[15:8] <= inBuf[inIdx][231:224];
              5:  inSamp[15:8] <= inBuf[inIdx][215:208];
              7:  inSamp[15:8] <= inBuf[inIdx][199:192];
              9:  inSamp[15:8] <= inBuf[inIdx][183:176];
              11: inSamp[15:8] <= inBuf[inIdx][167:160];
              13: inSamp[15:8] <= inBuf[inIdx][151:144];
              15: inSamp[15:8] <= inBuf[inIdx][135:128];
              17: inSamp[15:8] <= inBuf[inIdx][119:112];
              19: inSamp[15:8] <= inBuf[inIdx][103:96];
              21: inSamp[15:8] <= inBuf[inIdx][87:80];
              23: inSamp[15:8] <= inBuf[inIdx][71:64];
              25: inSamp[15:8] <= inBuf[inIdx][55:48];
              27: inSamp[15:8] <= inBuf[inIdx][39:32];
              29: inSamp[15:8] <= inBuf[inIdx][23:16];
              31: inSamp[15:8] <= inBuf[inIdx][7:0];
              default: $display("Unexpected number of bytes read for inSamp");

            endcase // case (inBytesRead % BUFFER_BYTES)

            // until next clock tick, inBytesRead is still previous value
            inBytesRead <= inBytesRead + 1;
          end // if (iCtr == 0)

          if (iCtr == 1) begin
            // sign input sample is valid
            inValid <= 1'b1;

            if ((inBytesRead % BUFFER_BYTES) == 0) begin
              inIdx <= inIdx + 1;

              $display("inBuf[%d] = %h%h%h%h%h%h%h%h", inIdx + 1,
                   inBuf[inIdx][255:224],
                   inBuf[inIdx][223:192],
                   inBuf[inIdx][191:160],
                   inBuf[inIdx][159:128],
                   inBuf[inIdx][127:96],
                   inBuf[inIdx][95:64],
                   inBuf[inIdx][63:32],
                   inBuf[inIdx][31:0]);

            end // if ((inBytesRead % BUFFER_BYTES) == 0)

            // Prepare for next state
            iCtr <= 0;
            inState <= IN4;

          end // if (iCtr >= 1)

        end // else: !if($eof(instream))

      end // case: IN3


      IN4: begin
        // update the sample counter
        if (iCtr == 0) begin
          sampCount <= sampCount + 1;
        end


        // wait for encoder input ready assertion to confirm the new sample was read
        // by the encoder.
        if (inReady) begin
          //$display("Sample count: %d, iCtr: %d", sampCount, iCtr);

          // read next character from the input file
          case (inBytesRead % BUFFER_BYTES)
            0:  intmp <= inBuf[inIdx][255:248];
            2:  intmp <= inBuf[inIdx][239:232];
            4:  intmp <= inBuf[inIdx][223:216];
            6:  intmp <= inBuf[inIdx][207:200];
            8:  intmp <= inBuf[inIdx][191:184];
            10: intmp <= inBuf[inIdx][175:168];
            12: intmp <= inBuf[inIdx][159:152];
            14: intmp <= inBuf[inIdx][143:136];
            16: intmp <= inBuf[inIdx][127:120];
            18: intmp <= inBuf[inIdx][111:104];
            20: intmp <= inBuf[inIdx][95:88];
            22: intmp <= inBuf[inIdx][79:72];
            24: intmp <= inBuf[inIdx][63:56];
            26: intmp <= inBuf[inIdx][47:40];
            28: intmp <= inBuf[inIdx][31:24];
            30: intmp <= inBuf[inIdx][15:8];
            default: $display("Unexpected value");

          endcase // case (inBytesRead % BUFFER_BYTES)


          // use sampCount because you inReady occurs at an unknown time count
          inBytesRead <= (sampCount << 1) + 1;

          iCtr <= 0;
          inState <= IN3;
        end

      end // case: IN4

      IN5: begin
        // sign input is not valid
        inValid <= 1'b0;

        if (iCtr >= 1) begin
          inDone <= 1;

          iCtr <= 0;
          inState <= IN0;
        end
      end // case: IN5

      default: inState <= IN0;
    endcase // case (inState)

  end // always @ (posedge clk)


  // encoder output checker - the encoder output is compared to the value read from
  // the ADPCM coded samples file.
  always @(posedge clk) begin
    eCtr <= eCtr + 1;
    if (rst) encState <= ENC1;

    case(encState)
      ENC0: begin
        eCtr <= 0;
      end

      ENC1: begin
        // clear encoded sample value
        encCount <= 0;
        encBytesRead <= 0;

        // open input file
        encIdx <= 0;


        // wait for reset release
        if (!rst) begin
          enctmp <= encBuf[encIdx][(BUFFER_BYTES << 3) - 1:(BUFFER_BYTES << 3) - 8];
          encBytesRead <= encBytesRead + 1;

          $display("encBuf[%d] = %h%h%h%h%h%h%h%h", encIdx,
                   encBuf[encIdx][255:224],
                   encBuf[encIdx][223:192],
                   encBuf[encIdx][191:160],
                   encBuf[encIdx][159:128],
                   encBuf[encIdx][127:96],
                   encBuf[encIdx][95:64],
                   encBuf[encIdx][63:32],
                   encBuf[encIdx][31:0]);


          eCtr <= 0;
          encState <= ENC2;
        end
      end // case: ENC1

      // encoder output compare loop
      ENC2: begin
        if (encBytesRead >= TOTAL_ENC_BYTES) begin
          $display("Reached eof of encryption file");
          eCtr <= 0;
          encState <= ENC4;
        end

        else begin
          encExpVal <= enctmp;

          // wait for encoder output valid
          if (encValid) begin
            if (!decReady) $display("Encoder output too quickly into decoder!!!");


            eCtr <= 0;
            encState <= ENC3;
          end
        end // else: !if($eof(encstream))

      end // case: ENC2

      ENC3: begin
        // compare the encoded value with the value read from the input file
        if (encPcm != encExpVal) begin
          // announce error detection and exit simulation
          if (eCtr == 0) begin
            $display(" Error!");
            $display("Error found in encoder output index %d.", encCount + 1);
            $display("   (expected value 'h%h, got value 'h%h). encIdx: %d, inIdx: %d, decIdx: %d", encExpVal, encPcm, encIdx, inIdx, decIdx);            

          end

          // wait for a few clock cycles before ending simulation
          if (eCtr >= 20) $finish();
        end // if (encPcm != encExpVal)

        else begin
          //$display("encoder output correct. expected %h, got %h", encExpVal, encPcm);

          // update the encoded sample counter
          if (eCtr == 0) encCount <= encCount + 1;

          // delay for a clock cycle after comparison
          if (eCtr == 1) begin
            // read next char from input file
            case (encBytesRead % BUFFER_BYTES)
              0:  enctmp <= encBuf[encIdx][255:248];
              1:  enctmp <= encBuf[encIdx][247:240];
              2:  enctmp <= encBuf[encIdx][239:232];
              3:  enctmp <= encBuf[encIdx][231:224];
              4:  enctmp <= encBuf[encIdx][223:216];
              5:  enctmp <= encBuf[encIdx][215:208];
              6:  enctmp <= encBuf[encIdx][207:200];
              7:  enctmp <= encBuf[encIdx][199:192];
              8:  enctmp <= encBuf[encIdx][191:184];
              9:  enctmp <= encBuf[encIdx][183:176];
              10: enctmp <= encBuf[encIdx][175:168];
              11: enctmp <= encBuf[encIdx][167:160];
              12: enctmp <= encBuf[encIdx][159:152];
              13: enctmp <= encBuf[encIdx][151:144];
              14: enctmp <= encBuf[encIdx][143:136];
              15: enctmp <= encBuf[encIdx][135:128];
              16: enctmp <= encBuf[encIdx][127:120];
              17: enctmp <= encBuf[encIdx][119:112];
              18: enctmp <= encBuf[encIdx][111:104];
              19: enctmp <= encBuf[encIdx][103:96];
              20: enctmp <= encBuf[encIdx][95:88];
              21: enctmp <= encBuf[encIdx][87:80];
              22: enctmp <= encBuf[encIdx][79:72];
              23: enctmp <= encBuf[encIdx][71:64];
              24: enctmp <= encBuf[encIdx][63:56];
              25: enctmp <= encBuf[encIdx][55:48];
              26: enctmp <= encBuf[encIdx][47:40];
              27: enctmp <= encBuf[encIdx][39:32];
              28: enctmp <= encBuf[encIdx][31:24];
              29: enctmp <= encBuf[encIdx][23:16];
              30: enctmp <= encBuf[encIdx][15:8];
              31: enctmp <= encBuf[encIdx][7:0];
              default: $display("Unexpected value when filling in enctmp");

            endcase // case (encBytesRead % BUFFER_BYTES)

            encBytesRead <= encBytesRead + 1;

          end // if (eCtr == 1)

          if (eCtr == 2) begin
            // This only happens because encBytesRead 
            if ((encBytesRead % BUFFER_BYTES) == 0) begin
              $display("Reading more enc bytes");
              encIdx <= encIdx + 1;

              $display("encBuf[%d] = %h%h%h%h%h%h%h%h", encIdx + 1,
                   encBuf[encIdx][255:224],
                   encBuf[encIdx][223:192],
                   encBuf[encIdx][191:160],
                   encBuf[encIdx][159:128],
                   encBuf[encIdx][127:96],
                   encBuf[encIdx][95:64],
                   encBuf[encIdx][63:32],
                   encBuf[encIdx][31:0]);

            end

            // Prepare next state
            eCtr <= 0;
            encState <= ENC2;

          end // if (eCtr == 2)
        end // else: !if(encPcm != encExpVal)
        
      end // case: ENC3

      ENC4: begin
        encDone <= 1;

        eCtr <= 0;
        encState <= ENC0;

      end

      default: encState <= ENC0;

    endcase // case (encState)

  end // always @ (posedge clk)


  // decoder output checker - the decoder output is compared to the value read from
  // the ADPCM decoded samples file.
  always @(posedge clk) begin
    dCtr <= dCtr + 1;

    if (rst) decState <= DEC1;

    case (decState)
      DEC0: begin
        dCtr <= 0;
      end

      DEC1: begin
        // clear decoded sample value
        decCount <= 0;
        dispCount <= 0;

        decBytesRead <= 0;

        // "open" input file
        decIdx <= 0;

        // wait for reset release
        if (!rst) begin

          // decoder output compare loop
          dectmp <= decBuf[decIdx][(BUFFER_BYTES << 3) - 1:(BUFFER_BYTES << 3) - 8];
          decBytesRead <= decBytesRead + 1;
          
          $display("decBuf[%d] = %h%h%h%h%h%h%h%h", decIdx,
                   decBuf[decIdx][255:224],
                   decBuf[decIdx][223:192],
                   decBuf[decIdx][191:160],
                   decBuf[decIdx][159:128],
                   decBuf[decIdx][127:96],
                   decBuf[decIdx][95:64],
                   decBuf[decIdx][63:32],
                   decBuf[decIdx][31:0]);


          dCtr <= 0;
          decState <= DEC2;
        end
      end // case: DEC1

      DEC2: begin
        if (decBytesRead >= TOTAL_DEC_BYTES) begin
          $display("Reached eof of dec file");
          dCtr <= 0;
          decState <= DEC4;
        end

        else begin
          // read the next char to form the expected 16 bit sample value
          if (dCtr == 0) begin
            // display simulation progress bar title
            //$display("Simulation progress: ");
            
            decExpVal[7:0] <= dectmp;

            case (decBytesRead % BUFFER_BYTES)
              1:  decExpVal[15:8] <= decBuf[decIdx][247:240];
              3:  decExpVal[15:8] <= decBuf[decIdx][231:224];
              5:  decExpVal[15:8] <= decBuf[decIdx][215:208];
              7:  decExpVal[15:8] <= decBuf[decIdx][199:192];
              9:  decExpVal[15:8] <= decBuf[decIdx][183:176];
              11: decExpVal[15:8] <= decBuf[decIdx][167:160];
              13: decExpVal[15:8] <= decBuf[decIdx][151:144];
              15: decExpVal[15:8] <= decBuf[decIdx][135:128];
              17: decExpVal[15:8] <= decBuf[decIdx][119:112];
              19: decExpVal[15:8] <= decBuf[decIdx][103:96];
              21: decExpVal[15:8] <= decBuf[decIdx][87:80];
              23: decExpVal[15:8] <= decBuf[decIdx][71:64];
              25: decExpVal[15:8] <= decBuf[decIdx][55:48];
              27: decExpVal[15:8] <= decBuf[decIdx][39:32];
              29: decExpVal[15:8] <= decBuf[decIdx][23:16];
              31: decExpVal[15:8] <= decBuf[decIdx][7:0];
              default: $display("Unexpected number of bytes read for decExpVal");

            endcase // case (inBytesRead % BUFFER_BYTES)

            decBytesRead <= decBytesRead + 1;
          end // if (dCtr == 0)

          // This could be problematic bc what if decValid happens at dCtr 0?
          if (dCtr == 1) begin
            if ((decBytesRead % BUFFER_BYTES) == 0) begin
              decIdx <= decIdx + 1;

              $display("decBuf[%d] = %h%h%h%h%h%h%h%h", decIdx + 1,
                   decBuf[decIdx][255:224],
                   decBuf[decIdx][223:192],
                   decBuf[decIdx][191:160],
                   decBuf[decIdx][159:128],
                   decBuf[decIdx][127:96],
                   decBuf[decIdx][95:64],
                   decBuf[decIdx][63:32],
                   decBuf[decIdx][31:0]);
            end
          end

          // wait for decoder output valid
          if (decValid && dCtr >= 1) begin

            dCtr <= 0;
            decState <= DEC3;

          end
        end // else: !if($eof(decstream))

      end // case: DEC2

      DEC3: begin
        // compare the decoded value with the value read from the input file
        if (decSamp != decExpVal) begin
          if (dCtr == 0) begin
            // announce error detection and exit simulation
            $display(" Error!");
            $display("Error found in decoder output index %d.", decCount+1);
            $display("   (expected value 'h%h, got value 'h%h)", decExpVal, decSamp);
          end

          
          // wait for a few clock cycles before ending simulation
          if (dCtr >= 20) $finish();

        end // if (decSamp != decExpVal)

        else begin
          //$display("Dec correct! expected: %h, got: %h", decExpVal, decSamp);

          // delay for a clock cycle after comparison
          if (dCtr == 1) begin
            // update the decoded sample counter
            decCount <= decCount + 1;

            //// check if simulation progress should be displayed
            //if (dispCount[31:13] != (decCount >> 13))
            //  $write(".");
            // update the display counter
            //dispCount <= decCount;

            // read next char from input file
            case (decBytesRead % BUFFER_BYTES)
              0:  dectmp <= decBuf[decIdx][255:248];
              2:  dectmp <= decBuf[decIdx][239:232];
              4:  dectmp <= decBuf[decIdx][223:216];
              6:  dectmp <= decBuf[decIdx][207:200];
              8:  dectmp <= decBuf[decIdx][191:184];
              10: dectmp <= decBuf[decIdx][175:168];
              12: dectmp <= decBuf[decIdx][159:152];
              14: dectmp <= decBuf[decIdx][143:136];
              16: dectmp <= decBuf[decIdx][127:120];
              18: dectmp <= decBuf[decIdx][111:104];
              20: dectmp <= decBuf[decIdx][95:88];
              22: dectmp <= decBuf[decIdx][79:72];
              24: dectmp <= decBuf[decIdx][63:56];
              26: dectmp <= decBuf[decIdx][47:40];
              28: dectmp <= decBuf[decIdx][31:24];
              30: dectmp <= decBuf[decIdx][15:8];
              default: $display("Unexpected value");

            endcase // case (inBytesRead % BUFFER_BYTES)


            decBytesRead <= decBytesRead + 1;

          end // if (dCtr == 1)

          if (dCtr == 2) begin
            dCtr <= 0;
            decState <= DEC2;
          end // if (dCtr == 2)
        end // else: !if(decSamp != decExpVal)
      end // case: DEC3

      DEC4: begin
        // "close" input file

        // when decoder output is done announce simulation was successful
        $display(" Done");
        $display("Simulation ended successfully after %d samples", decCount);

        decDone <= 1;

        dCtr <= 0;
        decState <= 0;
      end // case: DEC4

      default: decState <= DEC0;

    endcase // case (decState)
  end // always @ (posedge clk)

/* */
  //------------------------------------------------------------------
  // device under test
  // Encoder instance


  ima_adpcm_enc enc
    (
     .clock(clk),
     .reset(rst),
     .inSamp(inSamp),
     .inValid(inValid),
     .inReady(inReady),
     .outPCM(encPcm),
     .outValid(encValid),
     .outPredictSamp(/* not used */),
     .outStepIndex(/* not used */)
     );



  // Decoder instance
  ima_adpcm_dec dec
    (
     .clock(clk),
     .reset(rst),
     .inPCM(encPcm),
     .inValid(encValid),
     .inReady(decReady),
     .inPredictSamp(16'b0),
     .inStepIndex(7'b0),
     .inStateLoad(1'b0),
     .outSamp(decSamp),
     .outValid(decValid)
     );

endmodule

test t(clock.val);
