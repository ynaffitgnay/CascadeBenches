//---------------------------------------------------------------------------------------
//  Project:  ADPCM Encoder / Decoder 
// 
//  Filename:  tb_ima_adpcm.v      (April 26, 2010 )
// 
//  Author(s):  Moti Litochevski 
// 
//  Description:
//    This file implements the ADPCM encoder & decoder test bench. The input samples 
//    to be encoded are read from a binary input file. The encoder stream output and 
//    decoded samples are also compared with binary files generated by the Scilab 
//    simulation.
//
//---------------------------------------------------------------------------------------
//
//  To Do: 
//  - 
// 
//---------------------------------------------------------------------------------------
// 
//  Copyright (C) 2010 Moti Litochevski 
// 
//  This source file may be used and distributed without restriction provided that this 
//  copyright statement is not removed from the file and that any derivative work 
//  contains the original copyright notice and the associated disclaimer.
//
//  THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, 
//  INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND 
//  FITNESS FOR A PARTICULAR PURPOSE. 
// 
//---------------------------------------------------------------------------------------

include ima_adpcm_enc.v;
include ima_adpcm_dec.v;

module test;
//---------------------------------------------------------------------------------------
// internal signal  
reg rst;        // global reset 
reg [15:0] inSamp;    // encoder input sample 
reg inValid;      // encoder input valid flag 
wire inReady;      // encoder input ready indication  
wire [3:0] encPcm;    // encoder encoded output value 
wire encValid;      // encoder output valid flag 
wire [15:0] decSamp;  // decoder output sample value 
wire decValid;      // decoder output valid flag 
integer sampCount, encCount, decCount;
integer infid, encfid, decfid;
integer intmp, enctmp, dectmp;
reg [3:0] encExpVal;
reg [15:0] decExpVal;
reg [31:0] dispCount;

  reg [2785279:0] infile;

initial begin
  infile = 2795280'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000ffff000000000000000000000000ffff00000000000000000000ffffffff000000000000000000000000000000000000ffff000000000000000000000000000000000000ffff0000000000000000000000000000ffff00000000ffffffff00000000000000000000ffff0000000000000000000000000000000001000000000000000000000000000000000001000100000000000100000000000000000000000000010000000000000000000000000000000000000000000000ffffffff000001000000000000000000ffff0000010001000000000000000000ffff0000000000000000000000000000000000000000000000000000ffff000000000000000000000000000000000000ffff00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff000001000100ffffffff000000000000000000000000ffff0000000000000000010000000000ffff000001000100000000000000000000000000000000000000010000000000000000000000000001000000ffff00000000ffff000000000000000000000000000000000000000000000000ffff0000010001000000000000000000ffff0000010001000000ffff01000100000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000010001000000000000000000010000000000000000000000000000000000000000000000ffff000000000000000000000000ffffffff0000010000000000000000000000000000000000000000000000ffff0000010000000000000000000000010001000000000000000000000000000000000001000100ffffffff00000000ffffffff0000000000000000000000000000ffff0000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000ffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffff0000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000010000000000000001000000ffff0000000000000000000000000000000000000000ffffffff00000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000ffff000000000000ffff000000000000ffff000000000000000000000000000000000000ffff0000010001000000ffff00000000000000000000000001000000000000000000ffff000001000100000001000000ffff00000000010000000000000000000000ffff00000000000000000000000000000000ffffffff00000000000000000000000000000000000000000000ffffffff00000100000000000000000000000000ffffffff00000100000000000000ffffffff000001000000000000000000000000000000000000000000000001000000000000000000ffff0000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000ffff0000000000000000010001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffff000001000000ffffffffffff0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000ffffffff000000000000ffff000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000ffff0000010001000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000ffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000ffffffff00000000ffffffff00000000000000000000000000000000ffff000000000000000000000100010000000000000001000000000000000000000001000100000000000000ffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffff00000000ffffffff010001000000ffff000000000000000000000000000000000000000000000000000001000000ffffffff000000000000010000000000ffffffff0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000ffff00000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000ffff00000000000000000000000000000000ffffffff0000ffff000001000000000000000000ffffffffffffffffffff000000000000000001000000ffff00000100ffffffff00000000000000000000000001000100ffffffff000000000000000001000000000000000000ffffffff00000000000001000100010000000000ffff00000000ffff000000000000010000000000ffff00000100000000000000010001000000ffff000001000100000000000000ffffffff00000000000000000000000000000000000000000000000000000000ffff000001000000ffff00000000000000000100000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000ffffffff00000100000000000000ffffffff000000000000ffffffff00000000000000000000000000000000000000000100fffffffffffffefffbfffbff00000d0019001200f7ffe9fff8ff0000ecffdfffedfffcff02000f0019000a00f4ffeffff9ff03000b000f000c0009000a000c000f001a0027002e002a001600ffff0a002e002800f0ffd1ffe2ffedffe3fff8ff250032002200240033002d0015000600040009000e000700f8fff2fff7fffcfff9ffe7ffcbffc3ffd5ffd5ffbeffceff0b0028001c002d0048001900c1ffb6fff0ff0300d9ffb2ffaaffb4ffcaffe0ffe8ffeaffebffe2ffdaffe4fff9ff140031002400e0ffb1ffcefff9ff0e00470083005800030023007600370091ff58ffaaff020025002a00190008000f0012000400fdfff0ffc4ff9fff9aff8cff95ff00005900280007005b004400a2ffc0ff6000d1ff46ff220287078d0aec093e09120a4e0a6b093609bb099e094909b709220abd0949092909b6080108ba079a072f070507590771072b072d075207ee064506eb05a50546055805f0056706770664063f0610062006680688068406a406cb06d20608079b074e080209bb092d0a270afa09ec09e209e609390ac50a4d0bc80b260c3b0c360c5f0c790c3b0cea0bc30b880b3a0b450b9b0bc30bb60bba0ba90b540bfb0abe0a640afb09c409a1095e092f0938092d09ee08b5087808ff0773072207ff06e906f6061b072b07340754076d076b0776078c078207640767077d079407cf073a08a108f8085d09bb09ee09090a1e0a1d0a0a0a0f0a3c0a800ad50a330b780b960b9a0b810b430b030be30ad70ad00ad50adf0ad00aa50a740a420a0b0ada09b809920963093a091409e708bc0894085e081008bc076e07330723073e07610770076c0757072907f006cd06ca06dc06ff062d075607720786079807a807bd07d707ed07fe070f081f082f08410854085e08620864086308630870088b089f089e0886084c08eb0778071607d706b806af06ad069b066f062606c4055405ee049b045f043b042b04220413040204f403e203cc03b6039c037403470326031c032b0350038103ab03be03b903a6039803a103c603ff0344048704b804d204e004ec0409053c057605ae05d805ed05ee05e305d305c105ad058e0559051005b80464042104f303d103ac036e03100398021602a10146010901df00ba008d0052000e00c5ff81ff45ff0dffd5fe9efe6afe3ffe20fe0efe04fef8fddffdb6fd86fd58fd3bfd39fd59fd95fde0fd2cfe73feaffeddfe05ff32ff6bffb0ffffff51009e00d700f600ff00f800e700d400c600bd00b2009b00760048001100daffabff87ff69ff4dff2cff0affecfecdfeaefe88fe4ffefefd9bfd32fdd8fc98fc6dfc4efc2dfcf9fbb2fb65fb1cfbe1fab6fa90fa69fa3efa0cfae0f9c8f9c4f9dbf908fa39fa68fa8cfa9dfa9efa9afa94fa9cfab9fae5fa22fb6efbb6fbf7fb29fc3efc35fc12fcd9fba3fb81fb73fb7efb9afbacfbabfb94fb63fb2cfbf9facafaaffaa6fa9dfa94fa86fa64fa30faf1f9abf973f954f946f94df95ff95cf93ff906f9acf849f8eff7a9f791f7adf7e7f739f88df8bdf8c1f896f840f8e5f7a4f78cf7b5f71bf897f815f978f9a0f998f96ef92ff900f9f4f802f933f97cf9c0f9fef92efa3bfa34fa1bfae6f9adf97df952f93df93cf932f920f9fbf8b1f85cf811f8d3f7b7f7b7f7b2f7a3f77df72df7cff67bf62ef6fff5f3f5f6f50df62ff642f64df648f61cf6e0f5a8f573f560f57af5abf5f4f541f671f692f6a9f6a7f6a7f6b7f6c6f6e7f61bf750f795f7e5f720f856f887f89bf8acf8c8f8e3f810f94bf974f992f99ef982f95bf93cf91af909f907f9f9f8e9f8daf8b6f896f87bf848f80cf8ccf779f737f715f701f708f71af70ef7f0f6c3f67ef645f625f608f6fcf5fbf5e6f5cef5bef5a5f5a0f5b1f5bef5d7f5fbf512f630f65ef684f6b1f6e5f605f729f757f77ef7b8f709f84ff891f8ccf8e5f8f1f8f7f8e7f8ddf8dff8d6f8ddf8fcf81af945f978f991f99ef99ef981f96af966f95ff966f977f96ff958f936f9fbf8c7f8a3f875f850f830f8f8f7c2f799f771f762f769f767f767f769f75af759f773f793f7c6f703f82cf851f879f895f8bdf8f5f81ff947f96cf97bf991f9b9f9e1f916fa52fa74fa89fa96fa8ffa92faa5faaffabbfac6fabafab0fab5fac0fae3fa15fb33fb42fb43fb24fb05fbf3fae0fad5facafaa6fa7afa4ffa1bfaf8f9eaf9d6f9c2f9acf984f95ff946f932f936f950f966f986f9b0f9d6f907fa42fa76faabfadffa02fb2cfb65fb9ffbe3fb29fc56fc71fc80fc81fc91fcbbfcf1fc37fd82fdb6fdd8fdecfde8fde2fddefdd0fdc7fdc1fdb2fda9fdaafda9fdb0fdb9fdb0fd98fd71fd34fdf6fcc5fc9dfc8ffc91fc8ffc88fc78fc54fc2dfc0afceafbd8fbd2fbccfbcefbd4fbd2fbd3fbd9fbdefbeefb0efc37fc71fcb5fcf6fc3afd7dfdb8fdf3fd2efe65fe9efed3fefffe29ff4eff6cff8effbaffedff280066009a00c000d200cc00bb00a5008b0076006400530046003a003300340039003b00380028000300cdff8aff43ff06ffddfecefeddfe00ff2dff58ff72ff74ff5eff31fff5feb7fe81fe5dfe58fe70fea5fef3fe4affa0ffe9ff1c003800440045004b0062008d00d10029018401d80119023a0243023902270220022a023f025d027a02870289028102740271027a028902a302be02cf02d902d702c502af0296027d027302780283029502a2029902800256022202fc01eb01f101180250028602b702d702df02dc02d002be02b802c002d40208035403ad030f046104890489045c040e04c50392037f039a03d30310044d0476047e0476045a042c040204da03b503a603a503aa03c203e003f803170431043d044804460430041904fd03de03d403da03e8030a042d044204580463046504750488049b04b904d404e9040c0538056b05b50501063e0672068d068e0692069806a406ca06f6061b07400753074c0740072307f506cc06a3067e0676067e068c06a706b2069e0679063e06f305b805890561055105430531052c0527051d051f051805ff04e604bf049004750466045d04660469045e045b04560456047604a104cd04fe04160511050605f004dc04ea040d0544059a05f40548069c06d306e606e606c70698067c0672067e06b006e5060e07310739072c0727071e07140715070907ee06d806bd06a606a806ad06af06b406a4068006600637060e06f705da05b8059e057d055d05570556055a05690565054a052905f804c404a6048e047d047d04740463045b044d043c043704290412040404f103e203e903f203fa030b040d0403040104fb03f503fe03fb03ec03dc03be039f039a03a503c403fe033204540469045b0436041404f103dc03e803ff031e044904650472047b04740464045d0454044f045a0464046d04800489048d0499049e04a404b604c104c604cb04be04a1047f044d041304e403ba039f03a103ae03c003d003c0038c033e03d6026a021902e301d201e801080226023a022f020502cc0180013401fd00d700ca00d800ed00fe000801f900d500aa00790051003f003b0043005700660071007f008b009b00b800d600f5001701310146015d01710185019d01b001c201d701e901fd0113022202270223021002f701e001cb01bf01bc01bc01bb01bc01b501aa019e018b01750160014901330120010901ef00d200af008e007300600054004d0040002600fdffc4ff85ff4dff25ff13ff15ff22ff30ff33ff26ff0affe5febffe9dfe86fe7afe7afe83fe92fea5feb3febafeb4fea1fe88fe72fe67fe6dfe83fe9dfeb3febbfeb0fe98fe7cfe65fe5bfe5ffe6bfe7efe8ffe98fe9afe93fe85fe74fe66fe5cfe61fe76fe98fec7fef8fe1eff36ff39ff27ff0ffffbfef5fe08ff30ff5eff8affa3ffa1ff8bff6aff49ff3bff42ff57ff76ff92ff9fffa1ff97ff85ff78ff70ff68ff64ff5dff4cff3bff25ff08ffecfecbfea0fe76fe4cfe25fe11fe0efe11fe16fe0bfee1fda0fd4ffdfdfcc7fcb5fcc0fce6fc10fd28fd2dfd1cfdf5fccffcadfc92fc8bfc94fca9fcd1fc03fd30fd5cfd78fd7dfd79fd6ffd65fd70fd8efdb8fdeffd27fe52fe78fe97feaffecffef2fe11ff32ff4cff58ff62ff68ff69ff72ff7cff81ff88ff8bff85ff7eff72ff56ff37ff10ffe0febcfea6fe9dfeabfec2fed2fedbfed1feadfe7efe4afe15fef5fdeafdedfd05fe20fe2efe2efe17fee6fdaefd77fd46fd30fd31fd40fd62fd85fd9cfdacfdaefd9efd8efd7ffd73fd79fd8bfda0fdbffddcfdedfdfbfd02fefcfdf8fdf4fdecfdecfdf0fdeefdf0fdedfddffdd1fdc1fdacfda3fda1fd9ffda5fda9fda1fd97fd87fd71fd68fd6dfd7ffda7fdd9fd04fe28fe39fe31fe21fe0efefffd04fe1bfe3bfe66fe8ffea9feb8feb7fea4fe8ffe7ffe79fe8bfeb4fee5fe1fff50ff6bff75ff6eff59ff45ff36ff28ff25ff28ff27ff28ff24ff13fffbfed8fea9fe7efe5bfe43fe41fe4bfe53fe53fe41fe13fedafd9ffd6cfd52fd4ffd56fd60fd60fd49fd27fdfefcd5fcb9fcadfca9fcb3fcc6fcddfcfffc28fd4cfd6bfd7dfd7efd7dfd82fd95fdbffdfdfd3ffe7ffeb0feccfedafee2fee4feecfef7fe00ff0aff16ff22ff36ff54ff71ff8fffa4ffa7ff9eff8dff78ff6dff71ff7eff95ffadffbfffcbffd1ffcdffc3ffb0ff8dff61ff2ffffafecffeb5fea6fea4fea8fea5fe9dfe8dfe74fe5afe43fe2cfe1cfe16fe16fe23fe3cfe5bfe7efea2febbfecbfed1fecbfec0feb4fea5fe9bfe97fe99fea3feb7fecffeeafe04ff11ff11ff05ffebfecffebcfeb5fec2fee0fe04ff29ff47ff54ff51ff3fff1efff8fed5feb7feaafeb1fec7fee9fe0eff29ff36ff35ff23ff0bfff3fee1feddfeeafe06ff32ff67ff9affc5ffdfffe6ffdeffcfffbfffb9ffc2ffd6fff2ff11002b003f004c0053005900630070007f008e0098009d0099008f00820079007300730078007c007c00710053002300e3ff99ff50ff13ffeafedbfee4fefafe14ff26ff25ff0fffe5feaffe7afe54fe43fe4ffe72fea2fed5fefbfe0cff0bfffbfee6fed6fed4fee3fe05ff33ff65ff94ffb7ffcbffd1ffd0ffd4ffe7ff0f0048008e00d000030120012801230120012a0145017001a101c901de01d901bd019501690145012e0122011f0120011c0111010001e600c2009a006f004b00390039004d006f008d009a008d0064002b00f4ffccffbdffcaffe8ff09002100260018000100e5ffd3ffd6ffedff1b0057009400ca00f10001010001f700ef00f4000e0136016b01a201cb01e001dd01c4019e0177015501410141014f0166017f018e01900186016e01510139012801220123012501250125011f011c01200129013701480153015a015e015b015301490139012a01230126013f016e01a801e301110224021d020402e501d301dc01fd0134027302a802ce02e102dd02cc02b7029e028802760266025d025d025f0265026a0262024d022902f801c5019a0179016801620160015e0156014601320120010d01ff00f500ed00eb00ec00ef00f9000a0120013a01580174019001a901bb01c901d501dd01e401ec01f101f90104021002240240025e027c0294029d029d0295028a0287029202aa02cf02f8021c0339034a034a033b031c03eb02b00271023702120207020e021e0223020c02d80189012d01de00a7008c008b009500a100ad00b900c600dc00f5000a01150112010301f500f000f8000c01240136013d0138012e012e013b0152016f0185018e018c01840182019301ba01ef012b025d027e028c028702760266025b02560259025e02620264025e0249022802f701b901770138010501e700da00d500d300c700ac008600560029000a00fafff9ff050015002400310039003d0044004b0055006200720083009900ad00bd00ce00da00e200eb00f6000801250147016c019301b301c801d201ce01c301b901b201b201ba01c401c701c201ab01870161013b011c010901fb00ef00e000c600a50082005f00400027001000fcffeaffd7ffc6ffbcffb4ffafffacffa7ffa2ffa2ffa4ffacffbeffd3ffedff090021003800510066007b009200a700bb00cf00dd00ea00f9000401110122013201450157016201650162015401400129011001f900e800d800cc00c300b600a3008800600031000000cfffa6ff88ff71ff5fff4fff3bff29ff1bff0fff08ff07ff03fffefef6feeafee4fee9fef7fe10ff30ff4dff66ff7aff87ff96ffa9ffbdffd2ffe7fff5ff02000f001c003200520075009900b800cc00da00e100e300e600ef00f700000105010201fa00f000df00cd00b8009a00750047000f00d8ffa6ff78ff53ff35ff17fff9fedafeb6fe97fe7efe67fe57fe4cfe45fe47fe52fe65fe84fea9fecdfeecfe02ff0aff0cff08fffffefafefbfefefe08ff16ff26ff3bff51ff63ff74ff80ff86ff88ff86ff80ff81ff88ff96ffb1ffd4fff9ff1d00370043004300380021000500e3ffbcff95ff6dff47ff2bff1aff0fff0bff07fffcfeeffeddfeccfec6fecefee0fefcfe19ff2fff3dff40ff39ff2fff25ff1cff17ff12ff0dff0cff0aff05ff02fffafeebfed4feb3fe8afe61fe3cfe21fe17fe1cfe2ffe4afe66fe7efe92fe9ffea5fea9fea8fea4fe9efe95fe8bfe85fe84fe8bfe9cfeb5fed3fef8fe1aff36ff4eff5dff65ff6aff6dff72ff7fff91ffa6ffbcffcfffddffe7ffe9ffe4ffddffceffb7ff9aff76ff4dff23fff5fec6fe98fe68fe38fe0dfee8fdcafdb5fda5fd98fd8dfd82fd7afd78fd7cfd87fd99fda8fdb3fdb6fdb2fda8fd9efd96fd93fd9afda8fdbffde0fd09fe39fe6cfe99febdfed2fed7fecefebffeb0feabfeb2fec4fedffefefe18ff2aff32ff2eff20ff08ffe5feb8fe82fe45fe03fec2fd86fd52fd28fd06fdecfcd8fcc7fcb8fca8fc95fc81fc69fc4efc32fc16fcfefbedfbeafbf7fb18fc4efc95fce9fc45fda1fdf9fd49fe8dfec5feeffe09ff12ff0dfffffeeefee4fee8fe00ff28ff5aff89ffa8ffb0ff9dff72ff36fff0fea7fe60fe1ffee7fdb9fd97fd80fd72fd66fd54fd37fd0bfdd3fc94fc59fc27fc03fceafbd5fbbdfb9bfb6efb3bfb0afbe4fad3fadafafafa2efb6ffbb5fbf8fb33fc63fc89fca6fcc2fce3fc10fd4ffda0fdfffd63fec2fe10ff44ff5aff52ff32ff01ffc7fe8bfe51fe1efef4fdcefdacfd94fd83fd76fd66fd50fd32fd0cfde6fcc7fcb6fcbafcd1fcf5fc1dfd3dfd4cfd46fd2bfd00fdccfc96fc66fc3ffc26fc1bfc1ffc31fc4ffc70fc8cfc9afc94fc79fc50fc26fc0bfc0bfc2efc71fcc9fc28fd7ffdc6fdf8fd18fe2bfe35fe3afe3afe34fe2bfe1ffe15fe12fe17fe25fe3afe51fe68fe7ffe96feaefec9fee3fef7fe00fffcfeebfed5fec2febcfec7fee1fe03ff21ff33ff36ff30ff2bff36ff59ff97ffe7ff3c008600bc00de00f600130140018301d6012a0270029902a1028f026d024b022f021e0213020802fa01ec01e201e401f3010d0229023e0246024102380236024a027802c2021f038203db031e0440043c041304cc036e030b03b3026c0239021602f901d801b101810151012c011201ff00e900bb006a00faff72ffedfe8cfe59fe5afe83feb5fed9fee0fec9fea1fe76fe5bfe55fe55fe55fe4cfe31fe18fe11fe27fe71feedfe83ff2b00ca004701ae01fd0139027a02b702e60206030403dc029d024e020e02f40102024202a50207035a038803840361032603e402b5029002740268025a0251025c027e02c8023a03bd034a04bd04f104f104b6044404ca034f03db028f025c023d02450262028f02dd0234038e03ec03300451045b044e043804260425043d04560475049e04b104bc04d304d904dc04e804d704b90491043704c40342039002d6012f018d00280025005f00f900e101e502f103d1046d05c405d105b505830541051805fd04e004e80407052d058405fb0580062607c4074108a908e208e908d708ae0877083c08fc07b3075a070607c1068f06a106f5066e071708b40808092909e90841087407670634052a041c033902d001a001cd0171021a03c4034b043d04c703c7020f012eff16fdb8fac6f817f77df576f48af380f2c8f1eaf011f004f075f0aaf126f4fdf6c5f973fc14fea7feddfed9fe59ff1b0109043308550dc3123918671d042212264829822ba52c6f2c3f2b9c29ec273c273e28ee2a8f2fcd358e3c1d43c248764cd34dd14c49496343bf3bd9321e297b1f9816790eb0075f0288fdeff834f4d9ed95e5dddb22d056c33cb7e4ab80a2419c9098a0978399189d5fa240a9b9b0ccb840c130c984d017d7b5dcc3e191e6cbeb07f23af9dc01d40b10167f20a12a2a33533afe3f4443b8446c44ab413c3d6e37fe2f1d287820f1187412430d94083a04d4ff65fa8ef36bebeae148d734cc22c148b645ac8da33b9c03975394d493aa958d99389e10a39ea7e3aaccacc9adf5ade0ad5faed8af85b2a0b632bcdcc250ca7ed2c7dab8e26fea3bf19ff616fb2cfeb7ffd500780191016602d10346057107ca09620b970c080d1d0c560a9507700349fefaf735f086e730de42d48fcac5c102bacab384afcaac61ab17ab12abe6aa87aa91a951a856a795a6bfa655a8efaa51af87b5efbce0c51ed091da04e50fef7bf75afec80369071d0a5d0c060ed70f9c1196122813e5123c110d0f5a0cd8085a059601e5fcb8f79ef110eacde1f1d871cf53c6fdbd62b631b0aeab88a8dea6c9a6cfa76da974ab69ad7daec0ae95aeb5adb0acbeacc3adb3af69b333b8d0bc6bc161c56cc725c800c88ec61dc5c5c4f3c47cc60bca15ceebd225da37e275e987f06bf72dfe1806680f021a9126b6347b4372529560906cc075bf7b587efc7d9e7b27784c74e970476eab6b9b687c64cf5dfb532647c13642231c0ee6f7c8e19acdfabb7fad0fa3419c7e987d972798a799cd9b349e40a1e4a54daca9b46abf30cc71daede9fef9160a371a1b2a5939f7476f555261b26bf673d8798e7d127f6a7e257cab781474c46e0e69d5620b5cc654dd4c2644bd3aae30e825a71a500f080437f996ef63e7c8e04bdcd7d9f9d8ced9f6db94dea6e113e522e8feeaf7ed83f0c3f226f536f702f90bfbeefca8feb400a2023c04e7053407bb07d20739079d057e030a011dfe39fbcff8e0f6bef5bbf5caf6d3f8e5fbc1ffe7031e08170c5a0fd811b713f114d615e6162b18c319ed1b651ed4202e23162525265b268f2574231020721b81156d0e92063cfedef5ebed9fe638e0dada55d68bd278cfe6ccc2ca31c928c8b7c71ec854c947cb22ceded171d602dc82e2c4e9bbf116fa7602ac0a67126619a01fef243b29ba2c772f6831bc3274336833b5328331c42f8d2d0e2b46282225ab21d91d8d19d014c00f740a3205520001fc60f897f594f32ff25ef100f1e4f01af199f117f288f2edf20ff301f31bf370f328f49af5b7f750fa61fd97009e037b0615095b0b990df70f6612f814a5172d1a721c681ef11f13210022d4228f234b241525ba2516261b2681252b243522821f0f1c2418c513fb0e240a5905ac007dfcd2f879f580f2aeefa9ec6de9f6e54ae2c6deaddb2ed99cd70ad755d764d801daf1db21de85e020e305e629e978ecd5ef11f313f6cef839fb75fd92ff8a017e036105020761086309da09f309c40925093908fc062505d1021e00ecfc9bf992f6bff363f1afef3fee02ed00ecc7ea51e9d4e716e62ee467e2a2e0f5de8cdd34dc06db35da9cd95cd998d90fdabbda87db1ddc84dcbfdcb6dcb6dce1dc24ddd0dddede0de08ae137e3d1e4a3e6b0e8bbea13eda5ef0ef26ff4a8f65af8b9f9d0fa62fbb4fbddfba5fb45fbcffa15fa4bf97ff870f738f6d4f4f4f2a2f0dfed7deab7e6cbe2c4de07dbd4d71bd51dd3e1d119d1e9d046d1d3d1bdd208d45bd5ebd6b6d85eda24dc24de17e067e242e55ae8ecebe7efb6f36ef7fafae0fd5e008002ed03dd044005be04a503fc0198fffafc3ffa41f769f4a7f1a9eebbebb6e842e5ade1fcdd01da2fd6bad28fcf07cd44cb1fcabec92bca2ccba4cc76ce63d033d2d5d34fd58cd6a9d7f6d85bdad0db9bdd75dfe9e02ae209e312e3abe20fe2f1e0d1df2cdfc3defbde40e007e24ae43fe716ea81ecf2eefdf09ff2e0f410f87dfc3a038d0c281809266135c8443b53985fc4685a6e7c709c6f7a6c12685e63d65ebf5a39579f53394fa649f0416f37692acc1af8086bf60ae4cdd277c4aab97bb260afaaaf4fb2e0b654bcfbc114c84aceb1d412dc56e4a1ed86f85b048310271dd82961360743414fac5a5a65986edc75457b6a7e007f7e7d157ad2744b6e0767415f5957c24f9a48cf41713b5d35232f9528b921611ab612430b400406fe43f90bf62ef4e6f3e9f491f6fbf8fbfbc9fe81013f043f068e078d089e08d107ca062e051d035f01b7ff23fe40fdb8fc49fc55fc81fc7cfc9afc9dfc38fcb8fb20fb65fae0f9eaf9bffa96fc91ffba03c7085f0e3e14d319a61ea5229325562748287f280d285627702661257424a323c022d621af20df1e431cbc1811144c0eb407820009f9cdf12aeb4ce571e0b1dcfcd960d8ced726d872d988db32de6fe106e5c1e8b7ecc9f0e1f43cf9cbfd84029e07e80c3712a917e61c9f21e4256129bf2b1f2d582d432c322a5027b823d81f031c581809153912e70ffc0d660c0c0bb9094c08d0063a05a6036102860126017d01830211043206cf08920b5f0e1a115c13f714fc154116c815ed14b9132a1299100f0f5f0dc30b4b0ada08ba070e07b506ca063807b6074308d9086909140aef0a0a0c6d0d040fd810e312fa1436179619d61b031efe1f5321f421c5216d20121ef11a1317e312b40e9a0ad0065a030b00ebfcdef9bcf69cf36ef034ed27ea4ee7d3e412e311e2eee1d6e28be4dfe6bae9b7ec9cef67f2ecf42cf756f969fb6cfd64ff3001b602df039304e204d3045f04a903c502af017a0018ff6cfd82fb50f9c6f61bf472f1c5ee47ec11eaf4e70de67fe424e31fe29ee16de189e100e27ee2ede267e3b1e3e0e336e492e402e5a5e539e6afe607e710e7f2e6cce67ce63ee60ee69de507e535e4eee29ae165e047dfbfdedcde59df67e0c4e1f7e23ee48be5a4e6fce7a2e957eb5eed8fef7ef149f3d9f4faf5f5f6d3f764f8d6f815f9e7f86ff8b2f78df630f5aaf3def1efefebedb2eb60e910e7b8e492e2bfe022dfe5dd13dd63dcf7dbeddb0cdc93dcb1dd1adff0e050e3c6e554e8f9ea41ed43ef14f173f2c1f33bf5a2f63bf80afa9cfb12fd54fef3fe2cfff9fe14fed5fc2cfbd6f844f67ff367f09fed4beb39e9cce7e5e602e642e58fe496e3a1e2e2e143e1f0e0f8e020e158e1aae104e273e233e351e49fe51fe7afe8c3e93dea3bea73e9ede72de62ce4dfe1c0dfd8dde6db3bda09d918d8a9d7fcd7bed8e6d98edb2bdd8fde04e039e12ce2a3e3c5e5c0e88fed81f471fdbd082216b724e733d04232503b5b3e63bf67da68fd66e4627d5da1571452264dc048a144f73fd139b531f9265e199f0962f881e699d5b7c699ba36b2b1adb5ac05afc1b302ba37c175c85bcf0bd648dc6fe243e9c4f033f90203b40df918d624a830123c204749512d5ac4617467c06abf6b556a7266a6609c59b9519149da41c93a5a34d42e202ac125a321aa1d5619a514d90fdb0aed05ab0127fe7bfb23fa0efae1fab8fc4affd6015704b1062208bf08c808b3079505e90263ff26fbd4f659f2dced0feafee6b5e49be389e33de4b6e59ce793e985eb4cedcfee2df0acf199f322f68ef915fe7c0395094510f816391dda225327522adf2bcd2b2a2a5c279e235b1f101bdd16eb124f0fd60b6a08e8041301dafc33f810f389edb0e7bee107dcc2d645d2e3ceabccc3cb40ccf6cdd2d0a4d413d9f5ddfee2d1e771ecb5f065f4c1f7d1fa79fd0f00b40267058a084a0c95108c15eb1a2020cf2475287c2ace2a8529c2260023e01eba1ad7168a13ef10ec0e810d990cea0b410b790a3f095807c5049001eefd65fa78f78df500f5f1f512f8fffa55fe7f0126044e06c7078508d608a808cb078c060005230383018100440037015f035906ef09b70d30114414e416fe18c81a631cd41d211f47204c212b22e822c223c224d5251d275928fb28d0288027b1249d20801b9b158e0fb70939045fff1bfb45f704f444f1f9ee51ed27ec3deb7cea94e953e8e6e674e552e410e4ece4f4e628ea2bee89f2faf631fbfafe690291056808dd0ad80c270ea10e4c0e540df10b6b0a16091a086207cd061e06f6042903bf00c1fd7afa40f71bf42ff19aee14eca3e992e7c5e571e408e45ce446e5cee663e896e960ea77eadee901e9f9e7fce64fe6bde539e5cbe442e4bde370e352e397e33ee4f3e49de5ece578e577e418e388e176e042e0eee0aee23ae5fae7c9ea6ced9eef89f130f382f4a9f586f6e1f6d9f673f6c2f52cf5daf4c5f40ff589f5c4f59df5f3f496f3c2f1b0ef70ed4ceb64e98fe7e6e569e4dce27de18ee0f9df05e0e4e045e227e472e6abe8d4eaefecacee42f0d9f130f37df4d3f5e9f6f8f70ef9f0f9e8faf8fbd4fca5fd3bfe36feccfde3fc58fba2f9d9f7fef596f495f3bcf249f2f9f172f1f3f066f0abef1fefc5ee6cee40ee27eee2ed82ed0ded70ecd0eb58eb09ebe6ea08eb69ebe2eb82ec3fedc6ed16ee36eebceda3ec38eb4be9efe6ace47ce24be093de52dd3ddc90db4adb02dbddda04db28db8bdb91dcf7dddfdfa7e2d6e52de903ed21f187f507fb1502f40a3616cc230c332443db52cb60d36b21736676ca75ef71ee6bbd64435d69566750204b8546b641bc3b27341e2a231dd20da2fc7bea37d926ca59be09b751b4beb5d9ba47c2d7cad5d335dcb6e3bfea1cf135f7eefd1f05e70ccb15561f4c29ef33a73e17496353d25cd4646d6bf96ff371a4710e6f2e6ab663425c2454e94b2e443c3d39376832d62e282c0c2a402828264f23da1fd91b73177a137510690ebf0d750ec20f79116513a8144d15ac152e15ee136f120b109c0cb508ee0340fe8af8dff27bed45e956e6aae4aee41ce69ee847ecadf06cf573fa5dffdf03e807570b5a0e4a116a143318da1c36223328532ec7331e38df3a8f3b553a7d373d33142e7d28b722021d7e173612350d7508fa03ceffe0fb24f890f403f166edc1e927e6c0e2c1df58dd9bdb9fda6eda01db70dce0de40e292e6c9eb5df1cff6d7fbddff97024b040305f804dd04eb0434051d0695075209700bb00da80f47114a12491258118f0ff10ce909fc0671049902ba01c1016c0296030d058606fa078c09350bf60cda0ead102d124613ed1328144814a5145d157e16f1174a192e1a6d1ad11957183e1691135110af0c9808fd0339ff99fa6ef648f36cf1d8f084f10df3f6f4f7f6c6f85cfa02fcdbfd1900f30231069609fe0c1c10e2127915ec17721a3c1d1420b622c524b825482574236720981c8918a7143b113f0ea50b6009340726056f03f901cf00030019ffcafdf6fb78f9a4f617f442f26cf1dff160f367f58df74af926fa20fa63f91ff8b4f663f524f4d2f249f162ef0ced76ea05e802e693e4e6e3dee314e45ae48de48ae49ce414e5f7e56ee777e98eeb83ed49ef9af0aff1f4f26df456f6def884fbf3fde0ffa3001a0073feaefb42f8bff43af1faed0deb05e8e7e4b1e12ddec9dae2d763d59cd38ed2aad1e4d029d031cf71ce61ce12cfe7d0e7d383d773db5adfbee2b1e554e8a8eaf5ec39ef2ff1bff29df38df3cbf27cf1dcef7dee82edd3ec8cec5eecccebd8ea68e95fe73ee553e39ae172e0dedf6cdf30df23dfe9ded4de37dfe0df0de1d5e2aee47de62be83fe9dde948ea5aea66ea9feab6eabdeaacea2dea7ce9bde8cde713e7a3e631e6f5e5bae509e52ae41fe3c0e1b8e04de04ee028e1b8e255e416e6d9e729e964eacaeb14ed7eee0df039f1e3f1fcf138f1c2ef01ee23ec6aea1de92be862e7a4e6c1e567e47de216e018dd8fd9e2d52ed26cce08cb24c882c570c329c25ac121c1b0c185c281c3dbc432c69cc7aec94dcc96cf1bd47cd953dfe6e5deecf2f3d5fbe4043b0f5f1b3529fc37f546f954c0606a69476e266f756cdd66625f10579f4eae466a3f8738c1318a2a1c2228185e0c90fe50ef4edf66cffcc032b5deaccca8fba8efacf6b3c7bc55c607d00dd961e18ce96ef14af9bf01690a0613e41b87249e2c8e34303c53434f4ad5505456b05a7b5d205eb65c74595454ba4d6746b13eef36fa2f452acc25f922ed21ef218c22612363230822871fe31b8717831357101f0e2c0d300d5a0d5d0dee0c700b02090f0674026afe72fa3df698f1d8ecd0e76fe253ddc2d8e7d452d23bd1a7d1c5d376d786dcd7e206eabbf1a5f93b011e08150eed12de164a1a8a1d1c2132259729102e0a32c834da35f334fd31512d562791208e199412f30bd5051200cefa29f6e7f124ee0beb56e8f7e508e44ae2a2e034df06de24ddbfdcf1dca8ddd9de8ce094e2ebe4d5e739ebf6ee3df3abf7a6fb2affd00117036003e602b1018400daffadff630014024804e906c9096b0cb50ea4100e1200139613d313cc13b613d5136d14c8151a183e1bd71e72225b25f026fd266f257222a31e8c1a8c1602130010640d2b0b43099c075d068b05f1047304d903d0024a0177ff84fdd6fbf1fa1afb7bfc1bffa002a406da0adb0e8312fd155019861cc71fdf2273255f2773289228f027eb26db25fd2472241f24a923c3224f212d1f741c74194c161113de0f910c2909bd057d02a6ffa0fdb2fcd2fc14fe1200370233049e052f062006a805ed0453040204d803d203d703b4037f0360035c0396030a0467045d04ae032102c4ffe0fcdef933f72df5f9f39bf3d4f376f465f56af67bf7b8f801fa46fb81fc61fdb7fd85fdb2fc71fb2cfa09f93ff801f80ff82cf82bf8a7f77cf6d3f4c5f299f0a6eefdec98eb5deaffe867e7abe5e3e36ae2a0e18ce12de268e3d0e422e653e73ce8fae8d6e9d1eaf5eb54eda9eed2efe9f0d9f1cdf220f4d0f5daf735fa75fc3afe3cff29ff05fe0bfc8bf910f7fcf47bf3b1f25bf223f2f4f18ef1e6f055f0e3efa4efceef13f037f044f0f3ef56efdfeea9eee8eedbef3bf1ccf260f4a0f588f62df79cf72df8eaf8c3f9b9fa8dfbf9fb04fca9fb0afb7efa3ffa78fa2cfb2efc47fd15fe68fe4cfe9efda3fcbefbcbfafef981f9dcf838f8cdf746f708f75bf7c9f77cf85df9c5f9dff9a0f9c2f8d0f7f1f611f6b4f5b4f5b8f5eaf5e1f555f587f45af3f5f1baf0a7efeeee8dee36eeeeed62ed60ec55eb14eab8e8e9e733e75ae6dde524e5ebe3efe2f8e1e3e05ae02ae0f2df01e032e030e03ee0aae057e165e24ee4d2e68ae9f1ece3f0f2f40cfaa1006e0854127e1ef22b643ae848cc5544608d67116b416b9c68f063465e0c58df51024cf745d53f4e3984319f28671e4112e704c4f611e853da8dce59c5e9bf60be55c086c5b7ccefd4a4ddc2e53ced77f41dfbbb01e30812105f17df1edf25692cac327638103ea74306490a4e6052b655b2570e58fe5675547050a04b2446fe3f083a8e349a2ff62bcd29cb28ec28b129542a5a2a682973278324fa20941d681aa917d11538146e12aa101d0e9a0aea06b00214fef0f9b8f542f116edade809e4d3dff8dbdad805d763d63cd79fd940dd4ce292e8b2efc4f74600a408b310d117a81d6d220726be281b2b372d502f72313d337634a33441334e30ae2b9725bf1e76172b107309390381fd82f80af426f016ede0ea8ee906e911e97ee9e9e936ea8ceacbea30eb12ec25ed59eebbefcaf06ff1e9f116f22bf2a6f285f3b1f43ff6f2f748f91bfa70fa17fa4ff9bdf878f8aff8d5f9a2fbbefd66004b0323064809970ccc0f0413e8150e187319031ade1976191a192019ad19941aaa1b841ca91c001c611ac5178d14ea10030d290957057901a2fdcff925f6e8f23ff065ee66ed0ded4aede0ed8fee6def8af0f7f1f4f392f6c8f983fd77017e0583095b0d2011dd146818c11ba81ebc20f4211d220221f61e181c7a18b114fd10650d3f0a91071505dc02d900ddfe05fd64fbd6f963f80ff7b3f54ef40ff305f25df165f113f240f3ddf47af6b0f77ff8ccf89af842f8d6f754f7d7f628f62df5faf367f2a0f0edee39edceebe5ea3deaf0e902eafee9fce908eacfe9a2e9bbe9dde95cea5ceb6decaded20ef59f07af1abf2a5f378f412f50ef567f41df30ef18beee2eb25e9a6e682e46ce26fe07bde3fdce9d9b5d789d5b2d36cd266d1afd04cd0d3cf65cf42cf35cf8ccf92d0edd1a7d3cbd5c8d79ed967dbcedc16de79dfa9e0d7e1f9e293e3dae3e2e370e313e308e30fe38de36ee422e5e1e590e6c5e6f0e622e715e733e76fe761e750e71ae762e686e586e434e3fde1efe0e0df21df9dde11deb1dd6cdd1cdd12dd58ddcadd99dea6df9ce08fe175e21fe3d4e3cde4ece567e74ce943eb49ed54ef0af177f2a3f33cf461f423f447f31ef2e0f06bef24ee32ed4becb6eb72eb1debf6eaebea97ea44eadde90fe946e88ae7a2e610e6e6e5e4e56fe687e7d9e899eaaaeca6ee8ff030f237f3b1f39ef3faf2faf1bff059efdced56ecd7ea5be9f0e7b4e67fe53ae4f4e268e16cdf35ddbcda03d87cd569d3d3d108d131d110d293d3b2d50dd880da26ddc6df4fe210e5d8e77eea71edaef036f4cff8dcfe710609107f1b0a280f3585413b4c7d54b459a05b955afe568f51254b4e44aa3d9037d231642ceb26b42085190f11ff06bbfbaaef4be3c5d7f0cd7ac644c26ac1a0c399c84bcfcdd69cdedde569eca8f262f8dafda3035409ce0e6914bb19ae1eb823af288a2d9e32af377f3c27415f45bf482f4b774c3d4c764a64473f43603e76390f356431c92e6f2d052d452d012eb12ed72e5a2e022d902a4e278f23471fd21a97164312da0da40937059b005bfc3ef857f42ff15deeafeb7be94ee700e508e334e1a1dfefde15df57e041e39ee772eddff43afd1106210f8717c71ec2241229c02b372da62d672df02c6c2ce42b552b9f2a8229c4276d258022fa1e2e1b55176e13c90f9c0cca098107de05a904dd039e03ca0343042805610681076b081809160950081d074705d302440059fd09faf9f60bf445f157ef2bee8cedceed77eef0ee65ef9aef70ef72efc6ef89f038f2e0f4a6f8ecfd9204750c7715e01e022863304737443c5c3f88400140433ea53b7e3838351c325c2f142d362b7b297827d1244a21e51cf317fb127b0ed60a5108ef067c06d406d00711097c0a130c740d800e600fb40f600fce0ed20d6b0c1c0bbc092908cf06930577040c0454044e054d070c0a3a0dca103e1436179919221be71b331c241c2c1c901c431d831e3e201a221824ef252827d427d027f2269125bd236321d21efd1bcd1889151f128c0e1f0bcd078d04a601fbfe71fc3dfa5af8c1f6a8f5fbf481f41bf48ef3aef2a6f1c1f03ef077f0a1f194f311f6dcf886fbb5fd4eff34005c00efff1bff06fee5fcf2fb5afb23fb51fbddfb79fcf2fc51fd65fd34fd0bfdd1fc7cfc47fcfbfb8afb43fbf9fa94fa43faadf992f820f72ef5cbf25af0e7ed8eeb6fe94fe71fe5d3e23fe0aadd55db4ed9ffd789d7bcd7bad85fda53dca6de21e171e3b6e5cee791e951eb1aede3eefdf060f3e2f595f83bfb85fd64ff9700fc00bf00e1ff89fe12fd8dfb05faadf869f70cf6b0f449f3b9f135f0d2ee71ed2cec08ebcce995e884e779e6ade550e533e575e529e603e70de850e982eab5ebfbec1fee44ef6ff063f136f2c7f2d4f296f20bf225f165f0dcef6aef64ef9eefbdeffdef43f068f0dcf09df188f2dff360f5aaf6dbf7c1f822f956f982f9a3f905fac7fab3fba6fc73fdbdfd3cfde7fbc8f9faf6e2f3dbf003ee8eeb85e99ce7c6e513e44ee29de04fdf2ede1ddd3ddc34dbb9d90cd83fd64ed4aad2a5d12ad168d180d223d44ad616d93ddcc0dfe5e363e820ed5ef2cef747fd2d0388097d10aa184522492da739aa464653615eb066526be86b7468b661b8586f4e04443c3a4b315e293722431b2d147d0cd7034cfae5eff7e44cda7ad050c8c9c248c019c158c542cc23d542df47e989f2edfae0019907ef0cd21167163e1bec1f0024be27e62a422d562f55312d3335357d37a2398a3b253d123e2c3eb13da33c083b5139d0378136bb35d4358e36ce37a5398a3bef3cc43da33d0e3c42396a356730b22aaf24281e371700102208b4ff2af799ee7ee685dfbcd946d552d276d079cf5ecfcdcfccd095d208d553d8b1dce7e111e850ef3ef7c8ffde08cc11281ab821cd270d2c9c2e612f7a2e6a2c972937269822f51e311b2017d412470e6909a40450007bfc89f9aaf782f615f666f6f0f6b0f7e6f843fabefb9bfd97ff660114037104230520056b04d8025f0033fd5bf9d7f4f4efdceaa0e5ade057dcb4d828d6e2d4abd484d55ad7c0d9a0dc03e0b9e3d5e77eec9cf128f708fdfe02e4087a0e8313f217981b4a1e242030216e212a219a20c31fcb1ebf1d751cd31ad018471627138a0f800b2407bf028ffec0faa0f764f503f48cf3f5f3eef443f6d9f76bf9cffa16fc46fd5dfe7fffd60061021204f105e007a409320b7d0c670d070e6e0e980ea30e960e490ec70d0c0df30b980a2709b20765067605f904ec043f05ea05c00692075d080b097509ac099a090e091e08c106eb04f302fc0012ff7ffd2ffcecfacaf99bf836f7d7f57cf421f303f20bf128f07cefe5ee78ee6eeeacee4bef6bf0bdf130f3c9f43cf690f7dcf8eaf9d7faa7fb20fc6bfc9bfc85fc65fc53fc14fccdfb7ffbebfa3dfa7df981f87df774f62df5d4f36ef2caf023ef92ede2eb3aeaaae8f1e631e596e3fee194e08edfb5de0ade9edd27dda3dc37dcbbdb4edb1fdbfadaeada05db07db09db2ddb41db70dbc4dbeddb0fdc2ddcffdbe0db06dc3ddcf0dc3bdeb1df84e1a5e39ae59de7b0e973eb28edcaeef5efeaf0b0f108f252f29ef2b4f2c8f2b0f209f2f7f05bef12ed87eae0e719e598e25de031de4edcb2da36d92dd8bbd7bfd770d8e0d9c8db2ede16e12ae459e798ea8bed1bf03ff2b3f38ff4f5f4caf44ff4b1f3c3f2bff1bcf07bef44ee30edf7ebe5ea05eaf7e817e888e7f6e6d6e652e701e82ee9e1ea8fec66ee66f01bf2b5f33cf553f628f7bcf7c1f76ff7d5f6c7f58ef44af3e6f1a5f0a8efd5ee43eeeaed8ded0ced56ec54eb10eac1e893e798e6fce5bee596e579e562e50ce590e442e4fde3bae3b2e39ee326e374e28de14ee011df2ede8bdd4fddb6dd6dde5ddfbae029e286e32ee5efe6ade808eb2aee34f2fef7ebfffb096816cb243334b4430a52ee5d7666ec6a346bc467516117594850ab47024063393b33212d4826d81dbf13f707c6fa3bed2de06cd424cbcac4a9c124c2c1c5fccb70d4dfdd7ce7f6f056f97300e306610c2b111316c31afc1e16238426df28a12acd2b802c842d1b2f2931e0330537e9393a3ccf3d573ee23dfd3c153c783b9f3bbd3c883eb84014431e457046fd46a4463445de42c93fd43b3a374332ca2cff263221141b9814e90d9a06b7fedcf620ef14e8aae2ecdef9dc08dd52de53e0e9e250e57ce7f2e988eca2efe8f3ebf888feea044b0b4f1119171e1c21205b237c25632660266825802301211a1ede1a7c172f14fe10dc0d0b0bbf08f10601064d06b707570a3e0edf12c917b01cdd20ce238225e125e924062391208a1d131a6e167112030e67098c044affe6f962f49eeef6e89ce3afdec0da27d801d78ed7a6d9eedc25e1dce5e5ea60f037f6b0fc2c04610c2b156e1e3b27df2e203548391f3b303ba239bd3642335f2f0b2b972602221e1d1e181e13120e160941048cff06fbe3f67df343f1b5f057f253f66dfc3b04f90c96155e1dd4237a286a2b1e2db12d692dba2c712b4f298826f6228d1ee0193d15cf100d0d080a9107b70559045803e2021703230436063d09240da6113716a81ac51e2222ec244e27ef28e7294f2a9c29b827d924cf20e91bcf16c411280d56092906720301018afe09fc97f962f7c7f5f3f4eff4dbf581f79bf931fc17ff120241057f08710bfd0def0ffa102b11ac109a0f370eb90c300b9609d007c70562038d0074fd46fa24f76df462f2f8f04ff067f0e1f0a7f1c1f2dcf3fcf460f6def76bf939fb0cfda7fe1f004701ec012502dd01ec0051fffafce6f93df631f216ee3beac4e6dde37fe160df75ddaadbd3d93bd838d7d6d66ad727d9b8dbfcded3e2c7e6b5eaa8ee71f218f6a5f9e2fcbaff06028a03520458048f033b026300f5fd2efb0cf87cf4dbf04eede2e906e7dbe443e382e282e2ece2e0e34ae5d0e69de8c9ea0ced7fef2ff2b4f4e6f6b3f8caf92afa0cfa8df9e9f862f8fef7b1f74cf773f613f52bf3bcf02beec6eb95e9e2e7aee6aae5f0e487e435e443e4dde4cae537e728e940eb95ed29f0aef240f5cef7faf9c6fb05fd68fd23fd44fcc6fa2af99df70ef6daf4e5f3cef2b2f166f099ee9aec94ea87e8e8e6ebe56be57fe507e697e61ae784e7aae7b0e7d4e70ee867e8fae89ee914ea64ea88ea43eaa6e9e8e8cce735e666e43ee28ddfc6dc2adaabd7bcd5a4d41bd42cd4e6d4d7d5f1d66cd802dab3dbd5dd20e06ce212e513e88feb4bf0d0f679ffb70a6d18f42760384a4844560c618c676169d26679609957a94dcb430d3bfd33652edc29a525c220961ab512fb08e4fd08f239e6aadb39d3a7cdb3cb53cd30d2c1d9bce212ec0ff5a5fca0028b07400b1f0e0e11cd132c16a818de1a831c251ec41f582171230b26ec28422cce2f153304366e38f6398d3a663aa53977385137aa368a3609374b38e1395b3b943c073d503c943ac337e933932f052b5e260422f61de719c6154611ff0b06067aff75f896f161ebf9e5c1e1d7ded5dca0db22dbf7da33db14dc71dd75df52e2a8e55fe98dedbff1cff5ebf9b5fde9009f038e058406c4067406bf050d059504560441043304e5031103bc01050004fe24fcecfa84fa2ffb24fd0a008f036f07fd0ace0dc70f9b104110050fe50cf90988069b024afed1f955f5f6f0c8ecc2e8dee401e126dd7bd934d6a6d33cd221d268d305d697d9bfdd37e2a6e6f6ea40ef90f31df80dfd4202ac070f0de711f215ef18861ad11a021a2b18b115f21201101f0d820a0e08db05090471020301c2ff89fe49fd17fc0dfb57fa2bfab8fa10fc14fe99005e03f5051408a2096f0a8d0a4f0ad1093209bf086b0804089e071a073d062e050e04d402b301e1005a00360096007101b3027704a6060409810bf80d1a10cd111513d3130f140014a51302133a122a11b30fe00d920bd108de05ca02bcffecfc3bfaa4f73bf5cef276f074eeb6ec6bebd1eaa4ead1ea5bebd7eb3cecc5ec51ed0dee3fefb4f05cf225f4a9f5d9f6b3f702f8f8f7b5f718f767f6b4f5bef4d0f3f2f2daf1d7f0faeff4ee21ee9fed1bede3ec0eed21ed43ed85ed7aed5eed6eed61ed63ed9bedb0eda0ed7eed10ed69eca9ebb9eab3e995e83ee7b9e5f8e3ede1d2dfb1dd8cdbaad911d8b3d6c9d549d517d560d507d6d6d6edd728d953daaadb1cdd81de20e0f1e1b2e39ae59be762e90ceb91eca7ed79ee19ef5aef76ef81ef4def12efdfee7dee34ee16eed7ede0ed12ee18ee45ee68ee49ee0deec6ed44edc4ec70ec21ecf8eb10ec2eec58ec94ecb7ecd0ece8ecf3ec16ed58ed9dedf9ed55ee7cee7aee59ee06eeb0ed7eed57ed53ed7aed84ed5eed16ed7deca6ebdeea31ead5e913ead1ea03ec99ed38efc0f022f22bf306f4cbf467f515f6bcf611f745f727f77cf6baf5d7f4a8f3b3f2d5f1aff0b0efb9ee7fed8fecf4eb69eb50eb9debeceb56ecc8ec04ed16ed17ed15ed21ed5eedf2edb7ee9cefa3f04ef165f11af123f0a1ee4bed1cec19ebafea81ea0aea50e911e823e6e5e3aae1aadf3ede89dd76dde6ddb1de8fdf56e024e1f5e1cfe228e450e685e980eec5f57fffe30baa1a072beb3bd24b5c595c63c368926933664f5f6d56f24ccd43f73bce35d6309c2c5c280a23431cd313cb0902ff40f474eadae2f7dd38dc02deb9e2d7e9eff296fcf305bb0ec815d41a7b1e6c20ef201e21ea205b202320fe1fa11f791f7a1f921f3520802147238a252128972aa72c602eb72fa4309f31f53287349f367639a03cfd3f9343d4465949184bba4bf64a0049034608426c3d8f387733502e50293a24f91eae1909140c0e18080f0238fc33f7e7f276ef43edceebe7eac5eadcea32eb48ecc9ede1ef09f39af658fa6bfefd01be0401076508f1082e09090997083808ea07b707b407ef077a082f090e0a220b010cac0c620dc60d0a0ebe0eb40f15114913e615b818ae1b2e1efe1fe820be208f1f621d6f1ae616f012b10e760a3f061d025afee2faadf7e8f46cf23ff08eee52edcbec1bed29ee31f006f343f6fbf9cffd4f01bd04e5079b0a740d59101313131602195d1b5f1db51ef31e751e3e1d371be418891643146f123811a810d0109211ca123f14a615e116cf175518be185719501a1e1c181f1d230228712d9332a33626398a399e37d933ac2e9f289422ff1c0218e2138310940d160bea08fe06780549047a0334035603fb0364057d076f0a610ef812ff17251dab214025b327a0284028f526bd24eb21c31e201b1c17ca12140e4509b4049e0078fd83fbbdfa36fbaffccdfe5e01fd03620698087b0af60b3a0d2c0ead0ee70ec80e260e510d370c930a8e080f06ea0240ff27fbbbf64ef227ee8aeabde7d3e5cce487e4b2e42ce5e7e5b9e6b4e700e98fea6beca2ee08f17ef3e8f50bf8d1f935fb0efc57fc27fc81fb87fa5df90af8adf652f5eaf389f234f1dbefa3ee94ed8feca7ebdaeaf6e91de96de8d5e78ee7b7e721e8d2e8b8e985ea38ebc9eb0cec36ec65ec7deca6ecdfeceaece7ecd7ec96ec65ec56ec47ec6fecbbeceaec1fed45ed24ed02ede7ecbbecccec13ed57edc8ed4bee97eee6ee3aef5bef87efcdeff6ef2ef077f095f0b0f0d5f0cdf0c2f0d0f0c7f0caf0f6f01bf151f1adf1eff11ef242f216f2abf115f119f0e3ee9eed1cec92ea38e9dee7b3e6e2e522e597e460e42ce421e45ce491e4e4e464e5c5e537e6bfe60be75de7c9e705e852e8b4e8d5e8f9e820e9ffe8dfe8bfe85de80ee8d7e772e741e74de758e7bde782e852e95cea8feb8dec74ed43eeb1eedfeee4ee9aee21ee9aedeeec20ec40eb36eae6e85ae79de59fe37ce17cdf9ddddfdb95dabfd91cd9d1d8dcd8ddd8ead825d94bd971d9d2d93ddabfda99db97dcb2dd31dfefe0f4e2b7e55fe914ee50f43efcd6050d11761d6f2a2e379e42e24b445221558454e950d74a5a43963b2f34c62da22861249620be1c1e185e12720b860340fb5df3a6ecf8e7cfe57ae60feaf9ef9ef75300d90860108316751a261c2d1c8f1acd17ed141512770fac0d840ccd0bc10b1c0cb70ce10d750f45117b13f1157e18311bfb1dd520cd23f126592af22d9d315e35e238c53bf23d223f0b3fd33d863b28381734892f982a93259520981bbe16f211150d4b08790389fec3f938f5f1f04fed64ea20e8c4e636e622e69de678e74ae83be94dea24ebf6ebf8ecdcedadee93ef3af08bf0a5f05ef0b5efe6ee0eee49edbbec70ec62ec85ecd7ec4eedd1ed76ee4def39f05cf1d7f290f4a4f635f91afc50ffd00247068609590c630e7f0f970f920e9e0ce5099006020370fff6fbd2f8f5f545f3dff0aaee97ecdeea82e994e850e8b7e8cbe9a6eb23ee2ef1bcf47ff845fce0fff802720543074f08d208f408b7085d08020887071507b1062e06af053b05c20466042604f90309046204fc04ec052c079d082b0aae0b0e0d460e3d0f0510bf1061110112ae123e139e13c1137713bb12a21133109c0e110dad0b8f0acb09580935095909c1096f0a500b5f0c9a0ddc0e1210471170128f13bf14f9152c174d183519be19c9192a19dd17f8158913b710bb0db10abc07ff0474021e0006fe1bfc5afacbf85ff71af611f53af495f32bf3f1f2e1f208f35bf3ccf34ff4c5f41ff55cf571f569f55af549f537f525f504f5d5f4a1f462f41af4dbf3adf398f397f3a2f3b7f3d3f3eff3fff3f5f3cff397f348f3e8f28cf241f20cf2f4f1f3f1fef10bf20cf2fbf1dff1bcf19af182f178f178f175f161f139f101f1bdf06bf023f0eaefabef6def22efb5ee1cee60ed88eca4ebcbea08ea6be9fee8b3e88de88ee8afe8fee886e933ea04ebfbebf2ece2edd5eebbefa1f0a7f1c8f20df47df5e8f639f863f93efacffa38fb79fbacfbeefb2ffc73fcb9fce0fce6fcd2fc8bfc28fcc0fb3ffbb5fa2dfa8bf9e6f852f8bef740f7e2f688f647f62cf619f628f673f6d4f658f711f8d0f895f965fa15fbabfb32fc7dfc8ffc74fc06fc5bfb96faa5f9a1f8a7f792f66ff549f4fbf2a7f173f04def6deef6edc1ede8ed6dee09efccefb2f073f126f2cdf220f34cf363f328f3ddf2acf260f238f25cf28cf2ecf287f3fff355f482f42cf463f34af2d3f04aef02ee04ed87eca6ec31ed05eef8eeb6ef0ff0e8ef37ef0eee7eecc4ea0be954e7e1e5d3e4fae37ce362e34be346e351e317e3c3e279e201e2aae1afe1cce145e25de3cae4c8e6b3e970ed3cf26ff8e8ffab08b6128a1dbf28d033c83def45bd4b844e2d4e1e4bc145f43ec737eb30f82a4726a522c31f2d1d571afd16f6123f0e43095e040f001efde2fba8fcd0ffde04480baf12cd19b51f38246a260f26f8231320c91a84157610ec0b010987073c07a0081e0b2b0e09121f16031a0c1edb214225ad28f32b112f6032bc3520399b3cce3f8d42ac44b5459c456844ee416e3e3f3a83358c30b12b1427e7224c1f461cdb19ee174b16de147913e1111710210ef50bc809cd0702069904af031403c702d202da02d8020003cf025202db01e8007fff12fe3ffc17fa2cf845f673f43df37af21df273f244f35ef4d2f562f7e1f853faacfbe9fc13fe3aff6d00a601f902840443064408980a230dc00f341234147815af15cb14ea121310af0c3609cd05e002c60053ff9efea9fef9fe74ff0b005a00710073003f0024006100ec000802b603b8050908650a730c2d0e510fbd0fb40f2d0f3c0e420d400c300b4e0a8309b208f7074a07a4062b06eb05f805630621072a087209dd0a510cb10ddf0ecd0f6c10bc10d110bd109e109110ac10f6106211dc11491275124d12cf11f610e10fbf0eab0dda0c7d0c910c190d190e680fe5107112dc130415e7158816e5161f174f177a17a717c617c2178a170f1745162d15d01329124610380efd0ba1094207ee04bd02c30004ff8efd61fc6ffbc3fa68fa43fa48fa77faacfad2fae7facffa88fa23fa8ff9d2f811f847f77cf6cff52bf58af4fff368f3b4f201f238f15cf09feff7ee79ee53ee66eea7ee2fefcfef7ef055f128f2f2f2bef352f4abf4d8f4b9f471f427f4ccf392f389f380f38ef3aaf39af383f369f329f3f4f2c3f265f204f28ef1d5f013f04bef5eee8bedccecf3eb28eb66ea82e9b4e80fe87fe738e73ae74ee785e7d9e710e84ee8aee80ce986e92deac0ea45ebc8eb10ec34ec5bec5bec52ec60ec54ec49ec5cec5fec7aecc9ec18ed86ed19ee8fee06ef7eefe3ef65f0e0f01bf14df179f16cf173f19bf1b6f105f285f2f6f287f32df4aff43cf5c5f512f647f658f61af6c5f569f5f8f4adf495f48ff4aef4e2f4f8f4fcf4e6f490f410f466f372f256f134f007ef0fee7fed3bed4fedb1ed02ee27ee16ee96edcdecf7eb12eb64ea27ea35eaaeea99ebadecf7ed6befb9f0f1f101f3a1f3fbf313f4c2f357f3eaf253f2ddf189f11af1c3f078f0fdef81ef03ef5beebeed30ed98ec1fecc4eb70eb3eeb1eebfdeae7eac8ea9bea6cea25eacfe977e900e981e812e89ee745e725e71ee73de78be7dae72ce88fe8e6e840e9bee94deaffeaf7eb21ed95ee88f0fbf213f60afacefe5c04b60a84117f18691faf25e82ad42e013156311030522d90297c257321dc1d111bf81867172d16d9142c130311430e200bdf07d30486024b015e01ff02ef05ca09460e9e123516da180f1aad1918185915b411df0d170ab00650040c03f6024f04c606ff09dc0dd1117c15d518951bad1d5c1f9c2088216e22472329243e255a2663275028ce28af28f02766261f245c213b1efb1aed172d15e1122911f50f440f0b0f0e0f300f480f0e0f780e880d290c970a06096c070106da04b903b202cc01c400c1fff0fe20fe7afd28fde4fcb4fcabfc7cfc28fcccfb3cfb93fa06fa8df94df96ef9cbf958fa02fb88fbd7fbedfbc3fb7afb34fbfdfaecfa05fb3cfb99fb26fcebfcfbfd5fff0901d0028704f705e3063107e7060406ac0418036301bdff62fe62fdd4fccefc2cfdc9fd8afe2fff95ffc2ffb4ff89ff75ff98ff0c00de00ff015c03d8044b06a107ba087309c0099909f208e8079f063405da03bb02df014e010501e100ce00c100a70085006e0069007e00b7000d017001d5012e027202940294027e0258022c02190227025302aa0219038303e5032a043c042c04ff03b20366032403ec02d602ed022d03a4034f041b05f705cd068f073508c5085309e909860a300bd30b560cb50cda0cbc0c6b0cda0b070b030ab9082a077805a003b701ebff36fe9ffc44fb08faeef817f86bf7eaf6aff68df669f650f617f6abf531f59cf4eef350f3c2f23ff2e4f1a6f176f15cf143f119f1e2f094f031f0d3ef86ef5cef6aefa9ef1df0bdf070f13cf21df3fbf3e8f4ddf5b2f675f71df883f8c6f8f3f8f6f803f92bf950f995f9f1f924fa3efa31fabef90cf92df8fef6c0f592f45bf352f284f1c2f02bf0bbef38efc5ee66eef0ed8fed4ded04edd7ecc7ecb2ecb6ecd6ecfbec47edb6ed26eea9ee28ef74efa5efbaefacefb0efd9ef20f0aaf06df145f23ff341f41ff5eff5a3f61bf785f7e8f731f893f816f994f92afacafa3afb95fbd9fbe1fbe6fbf8fbeefbf6fb0bfceefbbefb7ffbfafa5dfabaf9ebf822f87af7d5f666f642f63ef675f6e2f64af7bcf738f896f8f4f85cf9b2f90afa5ffa8cfaa3faa3fa77fa43fa0cfabcf96df920f9baf85af810f8c4f792f77cf757f72ff703f7aff654f610f6d3f5caf50df671f6fcf6a5f726f883f8bdf8b0f883f84df8fcf7bbf791f757f729f7fff6aff65ef613f6b5f574f553f533f52cf528f5fdf4b9f442f480f390f270f12df000eff6ed2eedd4ecd7ec3aedffede6eee1efdff09df11cf26ef270f24cf236f221f238f29ff232f3f6f3eaf4dbf5c7f6b9f79ef891f9b3fa02fc99fd8dffd8018a04a107ff0a940e2d1281156918ac1a161cb81c9a1cc51b7f1aee181f174d158413b8110e10850e0a0dc80bbb0ad40947090e091c09a7099b0ae00ba20db60ff6118a142b17a319101c1b1e8c1f98200321b9202220301ff41def1c191c781b621b991bf01b861c001d341d541d301dd81ca41c791c701cc61c391dca1d9b1e5d1f1c20ff20b9215422f522462353234b23ef225422bb21f4201520571f821e981dba1c9f1b391aa918b5166e141a12ab0f560d720bee09e50885088908e808b309970a890bae0cb50da20ea60f7d102911e5116e12b912fc12ec127912d411bf103a0f8a0d930b72097c07a005f503b802c5011b01df00e3002601c3018e028603c1040a065807b908f109ed0abc0b2d0c320ceb0b450b410a1609c5075606f904b50385029401e80072004f007500c1003d01e3019c028603aa04fd058d073f09ec0a8b0cf00d020fda0f6710a710c210a2103610a50fd90ed60dd60cd70bdd0a150a6409b9083408ba074507f806c0069106810677066c0677068906a806e8062f077707c607f80708080608dd0794074107d3064d06c3052e0598041f04c60394039803c60313047c04f2046b05e7056806f60699075d084909550a6e0b8c0c8c0d4e0ece0efa0ebd0e280e3a0de70b500a820885068a04b3020a01b9ffc4fe09fe82fd0ffd7efcd2fb09fb1dfa3af975f8d2f76df736f70ff7f7f6c9f66ef6fcf56ef5c7f42ef49bf309f388f205f27cf103f18ff02df0f3efd1efd4ef0ef06ef009f1e8f1f3f22cf482f5c1f6e6f7e6f8a2f942fad7fa51fbcbfb43fc87fc9dfc80fc10fc6bfba4faacf99ff88cf75bf628f502f4dcf2d2f1f4f02cf086efffee79eef8ed7fedfaec7fec1fecd4ebbdebeeeb56ec05edf4edf3eef1efd8f078f1d0f1eaf1b7f156f1e3f05df0ecefaeef9defd5ef5df009f1d1f19cf232f397f3d1f3d5f3d0f3e2f302f450f4d3f465f516f6e6f6aaf770f830f9b3f9f7f9f7f98ef9def80df81ff746f6a4f51ff5bdf47af41ff4a9f326f37af2bdf116f175f0e9ef8fef49ef1fef2fef5fefbcef63f02cf110f21af317f4fcf4e2f5a6f651f705f8a2f826f9a6f9f4f90efa10fad9f97ef927f9b5f83bf8d6f75af7d6f667f6e1f55cf5f5f486f427f4f4f3bcf393f385f356f313f3caf248f2abf111f154f09befffee57eec1ed4bedc4ec4aece5eb64ebe4ea70ead9e947e9d0e851e8f4e7c8e79de78ce79ae799e7b2e7f7e74be8d3e890e94dea11ebcdeb4deca9ece9ecfdec0fed2bed3fed69ed9fedc2edebed0cee06eef7edd1ed79ed19edadec2beccdeb96eb7eebbbeb3fecf3ecfbed36ef7ef0eaf150f386f4a3f57ff605f759f76ef74ef738f728f729f767f7b8f707f860f891f898f89ef89cf8b0f810f9a8f97dfa96fbbefcecfd2aff5b009501ef025604d6056a07e808570aa30bb20c9e0d620ef30e7b0ff70f5610c01026116e11b811f111fc11fd11e4119e1159111311c710ad10c61008119a1165124a13571467155c164c171f18c6186719ed194b1aac1af61a201b521b6e1b591b2f1bc41a021a1519f017a0166a1547143e137a12d8114c11f910c110a610d4102b11a7115b121013b5135a14c614fd141b15f3148d140c143d132612e810570f860da90bb309d50752061e054e04f403d003cc03df03d803bf03b503ae03c40308045504a404ea04ff04ec04bf046a040804ab034103d9027e021f02c70180013201dc007e00030075ffe7fe63fe03fedffdf7fd47fec4fe50ffd6ff46009200bd00cb00be00a10073002d00d9ff77ff0affa9fe5dfe26fe0dfe06fef9fde2fdb1fd64fd10fdc5fc97fca0fce2fc56fdf7fda7fe51ffebff58009700ad0094006200360016001a005300a90010017901bd01d601cc01a20178016f018f01e70177022303dc038b0410056505840566052205c70460040d04d703b803be03e003090440047c04a304b604a6045404c6030103080201010f0038ff93fe1dfeb3fd4cfdd8fc43fc9efb01fb6ffa06fad2f9c3f9dff921fa6dfaccfa3afb9cfbfffb5ffca2fcd6fcfafcf5fcd8fca3fc43fccefb4dfbbafa37fad3f989f973f98ff9caf92dfaaafa27fbaffb33fca2fc0cfd69fdacfdeafd18fe2bfe35fe31fe12fef5fdd8fdb5fda6fda6fda6fdb4fdc3fdbefdb2fd94fd54fd05fda5fc2efcbafb50fbedfaaafa8afa82fa9ffad6fa10fb50fb84fb96fb91fb70fb30fbecfaa9fa66fa30fafef9bdf975f920f9c0f870f83df828f83ef874f8b3f8faf83ef97bf9c1f917fa76fadffa43fb8dfbb9fbc7fbb5fb95fb70fb41fb0cfbcbfa72fa0afa9cf92ff9d3f892f864f845f832f81df806f8f8f7ecf7e7f7f1f7fbf704f814f825f83df870f8b6f814f98ef912fa97fa1dfb8efbe6fb27fc43fc3afc1afcdbfb87fb32fbd0fa66fafcf97bf9e2f836f868f786f6a5f5c5f400f470f310f3edf20ef356f3bff33cf4a9f403f548f569f57ef599f5b4f5e5f531f680f6d5f622f749f74df72ef7e1f682f61ff6b8f563f520f5daf49af454f4f9f39bf33af3d4f282f241f20ff204f21ff261f2e1f290f35cf443f51ff6d6f670f7dcf727f875f8c4f822f9a6f936facefa79fb19fcb4fc58fde6fd65fedefe2eff63ff91ffa6ffc4ff0a006500f200b9018c0276036c043d05fe05b8064c07e8079c084a09160aff0ad90bc60cc50daf0eb20fc810c511cc12c71382142615a315d215ed15ea15ab1573154015ff1400154015a1155b1647172a182b19211ae11ab01b791c231df51dcf1e8a1f66203921e0219b223d23a02300242b240224d2237a23f12291223622d221ae21972174218c21a621ae21e4210722fe210422d7216b210b218d20f81fa51f681f401f6b1f9a1fb21fd91fbc1f4c1fca1e021e0a1d321c4b1b5e1aa419d418eb171c172b1629155e149d13fc12b01272123d122912e7117511fe104e10810fce0e060e3c0d960cd90b150b750ac7092709bc084c08e10791071e079a062c06af0545051305eb04da04ee04f004f20408050c05120527051905ef04b3044004b8033c03c00269024c024402590285029d02a902ac028a0256021502b3014401cf004900cbff65ff0fffe4feecfe17ff72ffefff7300f7006b01b501dd01e201c301970163012a01fb00d300af00990089007d007a0076006b005c0041001700e5ffa1ff4efff4fe90fe2ffee8fdbffdc7fd0bfe7afe0cffafff3e00b000010128013c0154017301af010c027902f4027403de03350476048d0482045804fa037703d20202021f013a004bff6dfea9fdeffc50fccefb55fbf5fab3fa74fa43fa19fad2f977f907f96bf8bff713f75df6bef545f5e1f4acf4b1f4d4f428f5a7f520f695f6f7f614f700f7c5f650f6cef55bf5e5f491f469f448f43ff44df441f430f421f4f1f3caf3c4f3c8f3fbf365f4d1f448f5bbf5ecf5ecf5c4f54ff5bcf425f471f3d0f25bf2f0f1b8f1bbf1c0f1d5f1eff1caf17ef11cf18af00af0c9efb3eff9efa1f065f14df23ff3edf364f4a4f479f40ff481f3b4f2eaf148f1b7f06cf077f09cf0ecf054f187f192f177f108f179f0ebef44efbbee67ee1beefeed18ee36ee7ceef4ee68eff5ef9df025f1acf139f29ef200f36df3aff3e2f30af4eef3b5f377f314f3c8f2b2f2abf2d4f22ef375f3b8f3f5f3f0f3cef39ff340f3e0f29df257f23bf260f298f2fff296f31af497f407f52cf521f5f4f485f408f4a3f344f320f352f3aaf339f4eef478f5d3f5f0f596f5e9f40af4f0f2e2f110f169f01df034f076f0edf085f1fef163f2b5f2caf2caf2c8f2aaf296f299f28af281f27df24df209f2b1f123f183f0deef1def6aeed2ed36edb7ec53ece8eb94eb56eb14ebefeae7eae1eaf9ea2ceb63ebc1eb47ece1eca8ed8bee63ef36f0e6f055f19bf1b6f1a9f1a2f1aaf1c3f10ef27cf2fbf295f327f499f4f1f41af513f502f5f0f4f9f44bf5e3f5c6f6f5f745f99dfaf5fb26fd34fe32ff1300ec00d101ac0289037004470522060e07f307e808e909d10aa80b5d0ccc0c0f0d280d0e0df00cdd0cc60cd40c020d320d850ded0d510edb0e850f3c1034115f12a4132515bb1631189719ba1a701be51b081cdc1bb11b861b591b631b7a1b781b7a1b481bc91a341a72199018e41765171f175817e417aa18c619ec1af31bf61cb41d1d1e661e5e1e0b1eaa1d121d541cb11b061b601af51988190f19a61807182c17471630150314071316124511bd103b10bc0f590fd10e2e0e9b0dec0c3d0cbf0b440be10ab60a850a550a3a0af50992092b099308e50746079006e1055505c0043604c8034503c3025302cc014c01e7007f00330018000c00250064009900c200cd008700faff2eff1dfefffc02fc37fbccfacffa1efbadfb52fcd0fc16fd11fdb2fc1bfc69fbb6fa32faf3f9fdf957faeefaa0fb55fce7fc33fd2ffdc9fc06fcfbfabef972f83ff73cf67ff511f5e3f4ecf419f552f599f5e9f53ef6a5f614f778f7c8f7e9f7c7f771f7f1f662f6fdf5ddf512f6aef68ff784f866f9ecf9dcf924f9a7f76df5b3f2aeefb9ec4eeac1e863e875e9e5eb7aefdff376f8a7fcf6ffe70147023401e3fecafb8ef8acf59bf3b8f201f354f46bf6c4f8e5fa76fc17fdabfc51fb2ff9a3f62af422f2eef0e1f005f246f46df7fdfa72fe5001150375036a021100c6fc18f98af59cf2baf00cf08ff01ff265f4fbf68bf9b5fb37fdf9fdf1fd32fdf3fb6cfad3f86cf75ef6baf58cf5c4f537f6cbf65bf7bef7f4f701f8ecf7e0f700f855f8fcf8f3f917fb58fc95fd9efe67ffe4fffbffbcff34ff5afe4efd2dfcfcfae6f90af961f801f8e5f7e3f7f4f70af801f8ecf7dcf7c5f7cbf7f8f730f87df8d3f807f921f91ff9e2f881f805f857f796f6d0f5f5f42ef48cf3fdf29ef272f251f24cf25bf25bf26af28df2b1f2f8f268f3e3f382f43bf5ecf5a7f664f701f894f814f962f998f9b3f9a1f986f96bf949f945f963f991f9e6f955fac0fa38fbaefb0afc65fcb6fcedfc22fd4cfd5afd64fd64fd52fd4ffd5afd70fdacfdfffd56febafe10ff42ff5fff59ff35ff11fff0feddfef0fe21ff67ffc7ff27007800bc00e000e400da00be00a00096009e00c400150181010a02ae025303f5038d040305590591059c058b0564051d05c8046404e3035603bf0217027e01ff009b0071007e00b10011018701f0015702a802d502fa0214031c0332034a035a037f03ae03e0033704a7042405c6056f0603079207fc07300852085a08490856087a08af081e09ac09430a010bc30b740c3a0df70d9d0e550f011093103811d1115112e5126a13cf133c148c14b014da14ee14e514fa140d1512153a155715551567156515481550155f157415cd154316c9168f175d181719e719911afe1a641b951b8c1b911b7d1b551b611b761b911bf31b631cd41c771d061e691ecf1ef51ed11ea91e521edd1da11d7a1d761ddc1d6c1e161f0320d7207a21122252223a220d229821ef205f20b31ff71e6f1edb1d431de61c821c211cf71bbb1b6d1b3c1bdc1a571ae6194b199e181e188e170117ab164816eb15c2158c155c155e1548152a152515ec1491143c14ab1301136d12b9110c1191101010a80f760f340ff40ec50e600ede0d570d9b0cd70b300b7f0af0099d095209320948095c098809c709db09d309a609200964088107600639051d04f302e601f600070040ffa3fe1afec9fda1fd7efd6efd53fd0bfdaefc31fc8cfbe8fa44fa99f90df990f819f8c3f777f72ff700f7d3f6a7f697f691f698f6c4f6f6f629f765f784f78bf78df776f75cf755f744f732f71ef7e0f682f610f67af5e4f46cf4fef3b4f391f367f342f31df3d5f287f23df2dff18bf143f1e2f083f023f0a8ef39efe1ee8eee6fee86eebaee2eefd5ef8bf067f155f22af3fff3bff449f5bcf50ff624f623f604f6b1f55bf505f5a5f473f46df47ff4c6f428f579f5cef50ef620f62ef636f62df641f66ff6a1f6fcf672f7e4f76cf8f1f849f985f98ef946f9d4f83cf87bf7caf635f6b2f569f54ef53ef54bf55df54bf528f5eaf477f4f9f37df3fbf2a4f284f284f2bef229f396f316f49ef406f56cf5d4f524f67ff6eff64ff7bcf732f883f8c0f8e6f8cbf88bf837f8b2f728f7b0f629f6b6f561f5f9f497f445f4d8f378f33df308f303f33ef380f3d8f339f453f431f4d3f305f3faf1d9f08def57ee5ded79ecdaeb8beb50eb47eb6eeb7deb8beb92eb4eebe4ea64eaaae9fce884e827e825e88fe824e9fce904ebe8ebbfec81edf3ed45ee89ee92ee9beeb5eeb2eec9ee02ef25ef62efb4efdeef0ef042f04bf05ff085f08ff0aff0dcf0def0e2f0e2f0b3f092f085f067f06df08df093f0a8f0bdf0a5f093f081f04bf023f000f0bcef88ef5cef1aeff6eee5eec6eec5eed1eecaeedeee03ef24ef71efdaef46f0d9f07af10df2b6f25ff3f3f396f433f5b8f546f6c7f62ef79cf7fef74cf8a5f8f7f83af98cf9d8f917fa60fa9afac0fae7fafbfa00fb13fb29fb4bfb93fbeffb61fcf3fc8bfd27feccfe63ffefff7b00f5006601d8013a029502ef0235037203ab03d503030440048604eb0473050e06c7068e074a080209a909320ab30a2e0ba00b240cb60c4b0df90db40e760f57104f1155127613941491156916f616231704179416e21521155a14a1131d13c51292129512b012cf120013241335134e1360137413af1301146a14fb148d150b167816a91694165616de154115ae141b1496133a13e8129a1262121e12cf118e114111ef10b310751042103c1050108a1003118f112112b7121b1342134113ff1292122212a0111e11b7104f10ed0fa70f580f040fb30e380e940dd70cec0bef0a100a4709ad0856081308d907a3074207c4064706c105560523050a050f052d0530051805eb048c0415049f031e03ad0263022902120224023b02580277026d024202fb018501fb007300e4ff69ff0effbffe8bfe77fe6afe75fe98febafee5fe12ff27ff2fff29ff03ffd0fe93fe3bfedcfd74fdf3fc6bfcd8fb2bfb74faaef9d0f8f3f721f75ff6d3f57ef55af56df59cf5cbf5f9f515f620f634f654f683f6cef61bf756f77cf776f744f7fef6a4f648f604f6d2f5b7f5bff5d9f505f647f685f6bdf6edf6fcf6f0f6d5f6a0f667f638f608f6e3f5cef5b6f5a6f5a2f59af59af5a2f59af58df579f550f52af513f504f511f538f55ef587f5a5f5a7f5a2f5a0f5a3f5c6f506f64af692f6c0f6b8f688f635f6cdf580f563f580f5ebf595f65ff745f829f9f2f9a5fa35fb96fbd9fbf8fbf2fbe4fbd3fbcafbe4fb1efc6efcd6fc37fd78fd94fd77fd1dfd9afcf2fb31fb74fabef918f995f832f8f3f7e3f7f7f729f879f8d1f828f97cf9bef9eef913fa27fa30fa34fa30fa2ffa3dfa61faaafa25fbccfb9cfc82fd60fe1effa5ffe8ffeaffb6ff5efffafe9cfe50fe21fe0cfe0ffe29fe4ffe7cfeaefed9fefefe1fff34ff46ff59ff6aff83ffa8ffd6ff14006400ba0016016c01a701be01a7015701d90038007dffc0fe12fe74fdf9fca2fc67fc4dfc4bfc50fc59fc59fc3efc10fccffb7dfb30fbf0fabffaaafaacfabafad9fa03fb31fb6bfbadfbeefb34fc77fcb0fceafc24fd63fdaffd05fe5bfeacfee8fe03ff02ffe6febcfe98fe84fe88fea7fed8fe12ff47ff6cff77ff64ff2fffd9fe66fedefd4ffdc2fc46fce5fb9bfb67fb40fb13fbddfa9cfa4efa00fac0f98df973f976f98af9b8f902fa5cfacffa57fbd9fb51fcb0fcdbfcdffcc9fc97fc71fc67fc6bfc8bfcbdfcdbfcf4fc09fd10fd33fd86fdfefdb6fe9fff8b007c015a02fc028003e70325046804b504f6044d05b20508067506f60674071b08e208a4097e0a530bf80b8b0cfa0c2a0d520d6d0d6b0d820da80dc20dfe0d480e800ed50e320f7c0fe40f5610b4103011b01114128f1209136c13f3138d142715fa15e716cd17d118c619821a2e1ba21bc51bcf1ba71b431be51a791afb19ae197c1956197319a619d419201a581a621a6b1a4e1a021ac0196c190419c2188918541858186c188118ba18de18d718c3187118db1732175b1663158814b413f4127b122812f7110612201234125612571234121412e011a811981195119f11d011ff1126125c127e128e12a112941266122b12c9114d11d8105910de0f750ffb0e690ec00de80cf00bf80a040a300992081408af075707ea066306ca051a056804c8033603bc025c020302b5016c011f01d10082002a00ceff6dff03ff98fe2cfebefd56fdf2fc94fc45fc04fcd5fbbcfbacfb9ffb8efb6afb35fbfcfac4faa6fab4fae5fa37fb99fbe0fbfcfbddfb75fbdafa28fa6af9c7f84cf8edf7aef780f743f7f9f699f615f680f5e6f43ff4a9f32cf3bcf270f24bf23af250f289f2cff22df39af3f7f34df493f4b2f4c1f4c6f4b5f4acf4aff4a5f49cf488f449f4f5f393f319f3b3f272f24af253f282f2aef2dcf2fdf2eef2caf29af252f21af202f2f9f11df272f2d7f25ef3fdf38af40ef57ff5b4f5c1f5adf564f50cf5bbf462f423f407f4ebf3dff3e0f3c2f39bf370f328f3e4f2b6f285f26bf271f26ff278f290f292f29bf2bcf2dcf21cf38ef30ff4b0f472f51ef6baf642f784f794f785f739f7d9f688f62bf6e8f5d4f5c5f5cff5f9f50cf616f61df6ebf596f52ef590f4e1f344f39bf210f2b8f166f12bf10ff1dcf0a9f08bf05df045f059f069f089f0baf0c0f0aef095f04af0f9efc0ef79ef45ef34ef13effaeef9eee2eed6eee6eee2eee3eeeeeeceee9eee74ee30ee03ee12ee40eeb4ee76ef4af033f122f2cef244f389f376f33ef300f3acf270f25df248f243f249f226f2f2f1b7f157f1f9f0acf04df0f5efa4ef30efb8ee47eec9ed6ded47ed41ed7aededed6eee0aefb3ef3ff0c0f031f173f19ff1b6f1a2f185f169f145f140f165f1a6f11bf2b9f25ff312f4b9f434f58ff5c3f5c9f5c6f5c3f5c9f5f6f547f6b0f637f7c7f74df8d0f844f9a5f905fa5efaaefa04fb56fba5fb04fc6efcebfc88fd33fee5fe95ff26009000d800f6000301180137017701da014602b502140344034c033103f302b90299029602cd023b03c3036a041705a9052e069906df061f0759078407bf07030842089b0804097209050ab10a620b330c060dc00d760e0c0f6e0fc10ff70f0c102f1055107610ba1008115011b71123128612091391130d149d141b156f15b815d415b81596155b150815d314a6147a147d149114ab14f8145215ac1528169a16ec1640176d17681762173a17f016b51667160016b1155515ed14a914681425140b14ed13be13a413751330130813e012c112df1211135213be1319144f147c146b142014d0136413f512be129e129812c312e012db12c7127212e5115311a110e80f560fc20e330ec00d3a0da50c210c8a0bf10a780afd098d0949090c09e808fc0826097409fa09870a1c0bbe0b370c890cc20cbd0c920c5f0c100cc50b970b670b440b310b000bb90a5f0ad60937099b08f3076307fd06aa067d06770673067b06860670064506020693051805a1043004ed03e20300045104bb0410054c054f0502057d04c103d602e601f40003002fff6cfeb4fd1cfd98fc25fcd9fba2fb7afb6efb61fb48fb31fb03fbc2fa88fa4bfa16fa02faf9f9f9f908fa02fae1f9b4f964f906f9b9f874f84bf851f863f883f8aff8bef8b8f8aaf87ef84ef830f810f8fef702f8faf7f0f7e9f7c7f79ef77df748f715f7ecf6abf660f611f69ef520f5a8f422f4b1f368f32ef31af331f34cf377f3aff3cdf3e0f3eff3dbf3c3f3b6f3a0f3a5f3d1f30bf464f4d9f43df594f5d8f5e0f5c3f58ef533f5d8f493f455f43af44bf469f4a5f401f55af5c0f534f691f6e6f635f75bf76ef778f765f753f757f75ef783f7cff71ef879f8dcf81bf943f95df950f93af936f92bf931f94ef956f94af928f9cbf845f8b2f704f765f6f5f5a2f580f597f5bcf5f1f538f666f688f6adf6b7f6bdf6d3f6ddf6f0f620f749f780f7d0f713f856f8a3f8cdf8e5f8f5f8dbf8b2f894f86af856f86ff893f8d3f82ef971f9a0f9bcf99bf959f909f997f828f8d1f775f72ef701f7c4f68cf65bf609f6b1f55bf5ecf487f43df4f6f3d8f3e5f3f9f325f459f467f462f445f4faf3aff373f33ff33ff374f3c0f335f4b7f41cf570f59af583f54ff5fff494f445f416f407f43df4a1f41bf5b5f547f6baf61ff75df772f784f783f776f780f78bf799f7c6f7f4f723f86bf8a6f8d7f811f92df935f942f934f924f92ff938f958f9a5f9f8f962faebfa63fbdcfb5cfcb5fc06fd5bfd8cfdc1fd05fe30fe6afebdfefdfe5affdbff59000301db01b102aa03b904a00582064e07d1073f089708b908ef083b097f09fc09a30a440b130cf20cae0d810e550f0410d210ac1169124b133114ed14bf1582160d17a7172e188018e6183b195c198f19ad1998199a1990196319661973197819c119201a791a0b1b9c1b0a1c941c021d401d9b1de61d181e801eed1e4c1fde1f5f20b72020215d2162217621662135212a211321ec20f720f920ed2012212a213221632179216f21782154210321c1205920d71f791f0a1f911e3f1ed81d5d1dfb1c761cd61b491b981acd1915193b184f177d169615ad14f0132e137a12f91177110211b6105d10ff0fb40f470fc60e4f0ebb0d280dbb0c560c130c0c0c150c360c760c9d0caf0cb20c780c110c900bd90a090a3e0964089c07f8065b06d6056605e6045f04d20325037402ca011c0185000f00a5ff59ff28fffafedbfec5fea0fe7afe48fef6fd93fd1afd7ffcddfb32fb7bfad4f935f99af814f895f716f7a7f63bf6d0f57bf530f5f3f4d5f4c5f4c2f4d7f4eef406f52df551f579f5b7f5f9f542f6a0f6f1f634f76df779f75cf722f7b6f62bf69cf5fdf469f4f9f399f356f338f314f3ebf2bbf25af2d9f14af19ef0f9ef7cef14efdceeddeee9ee06ef30ef33ef1feffeeeb0ee56ee06eea6ed58ed2cedfdece4ece9ece0ece1ecf4ecebece7eceeecd9eccaecccecb7ecb2ecc9ecd6ecfdec47ed85edd4ed36ee76eeb7eefeee25ef59efa8efe8ef41f0aff0f9f036f161f144f10bf1c8f05ff00cf0e4efc3efceef02f01df039f04cf01ff0dfef9aef2fefdceeb1ee8cee9beee1ee27ef8eef0df069f0c6f022f14ef178f1a9f1b8f1d8f10ef22df261f2aaf2d9f218f367f39cf3dff332f467f4a3f4e6f401f51df53cf534f532f53af524f51cf527f51ef52ff560f589f5d4f53cf691f6eff64cf773f787f785f74bf708f7c9f676f641f631f625f63df673f694f6b7f6cff6aff678f62ff6bbf54df5f5f49ff473f473f475f48ff4b3f4b0f49cf472f414f4aaf341f3c8f26ef23ef21bf221f248f261f27ef293f27ff262f246f21bf209f219f231f267f2b1f2e6f215f336f32af30ef3e9f2a8f26ff244f211f2f2f1e2f1c7f1b3f1a0f175f147f116f1cff08df052f00ff0dfefbfef9def91ef93ef8fef98efa3ef9cef99ef92ef80ef81ef98efc2ef19f095f021f1c3f15ef2d7f236f36ef37df384f389f39af3d7f339f4b9f461f512f6bbf65ff7e4f749f8a1f8e1f819f962f9b0f90efa87fa04fb86fb16fc9afc21fdb9fd50fefafebeff840055013202fb02c10389043c05f405b90671073408fe08af095f0a0b0b980b2a0cc00c400dcb0d5a0ec80e340f920fc40ff80f2b104e1099100a11881140121b13ed13d814bc1573162c17d7175f180519ba19681a461b341c0c1dfb1dd91e851f3720ce203721b32121226c22d2222a235c23a823e523022445248424b1240b256325a32508265c268c26d62605270c272c272f270b270127d92688265026f62574250c258724e1236123ca221c229621f9204320b31f0a1f4c1ebb1d171d671ce41b4a1b9e1a181a7919cf185a18e017721748171c17f016ed16c41678163616bd151f159914f1134513ca124312c41174110b1195103510a40ff70e570e8c0db50c000c360b750ae1093e09a4083008a7072107ba063706b3054405b3041a048f03e1022f029201dd003400aeff23ffb3fe70fe2dfe03fefbfde2fdcefdc6fda0fd79fd5efd2dfd09fdfafce1fcdbfceafceffc03fd26fd38fd4efd63fd56fd3cfd13fdc1fc65fc02fc8cfb23fbcafa74fa3dfa1ffa0bfa12fa2bfa41fa63fa83fa92faa2faa9fa9ffa9cfa97fa8cfa8ffa95fa98faa8fab6fabcfac7fac6fab6faa1fa79fa3ffa04fabef974f93bf909f9e5f8dff8e8f804f939f974f9b2f9f5f926fa45fa59fa52fa3dfa2afa10fa01fa09fa17fa34fa64fa8dfab5fae0faf5fa01fb07fbf3fad4fab1fa7bfa48fa23fa01faf5f905fa17fa30fa49fa3dfa14fad0f95ff9dff866f8ecf792f764f746f747f75ef765f768f765f743f71df7fff6d5f6bdf6bdf6b9f6c5f6e1f6faf626f759f779f79ef7cff7f0f71bf84ef86bf884f89bf892f884f878f85ef84ef855f85af86df892f8a9f8bff8d8f8daf8d3f8cdf8aef886f865f832f802f8e6f7c8f7b8f7c6f7d0f7def7f9f7fbf7eaf7daf7aff777f74ef720f7fdf6faf6f7f6f9f613f719f713f71bf70ff7fcf609f718f736f77ef7c3f706f85af890f8abf8cdf8d1f8cbf8e8f806f935f997f9f8f95ffae5fa4efb9dfbeffb10fc10fc12fcecfbb9fba0fb71fb49fb4cfb3cfb2bfb35fb1cfbf5fad9fa92fa3efafaf996f936f9f9f8abf86ef858f82df809f8f5f7bbf782f75ef721f7fbf6fbf6edf6f5f616f716f712f707f7c7f680f638f6d7f597f57bf562f582f5cdf50bf66ef6c9f6eff61af71cf7e5f6b2f671f616f6dff5c6f5b2f5caf5f9f52cf67ef6cef611f75cf78bf798f79ff782f74ef72ff714f711f74ef7b3f748f814f9e9f9c3fa97fb37fcb7fc1dfd4efd76fdadfde5fd46fed7fe79ff42002001ed01c50294033a04e1047905ed056d06e4064607c5074808c1086609170ac60aa40b850c570d3e0e090fac0f5710da103711a71100124b12c3123713ad135814fb149b1565161517b2176418ea184e19be19fd19251a6b1a931ac11a251b7c1be01b761cf11c611de11d241e491e731e651e4d1e561e461e471e7d1e9d1eca1e161f361f4c1f6c1f531f2d1f141fce1e891e601e151ed51daf1d631d171dd91c6a1cf71b911b071b881a201a9a192019bc183218a91728177416ba15071526144f138f12b311f3105510a00f020f7b0ecd0d260d860cb60bed0a330a56099408f107340795060e066405ce0442048d03e8024e028d01e200460087ffe4fe58feb4fd31fdc0fc35fcc4fb5bfbc9fa45fac0f913f97df8f2f74ff7cff663f6ecf596f549f5e3f491f438f4c0f360f309f3abf279f261f24ff260f26df263f25ff23ff200f2c7f182f137f10ef1eef0d3f0d2f0cdf0c8f0d0f0c7f0b4f0adf096f07bf06ef053f039f02ff01ef018f02af036f04ff081f0a4f0c7f0eff0f7f0f6f0fbf0ecf0ecf008f121f155f1a6f1e7f12cf27af2a3f2bef2daf2d9f2def2f8f205f32cf35ff37ff3acf3d0f3c8f3b2f394f34bf307f3dbf29ff27ef288f288f299f2bbf2b7f2aaf2a2f270f23cf21af2e1f1b9f1aff194f185f18df177f162f159f130f108f1f1f0b9f082f05af011f0c6ef88ef30efdfeea6ee5cee21ee03eed4edb1eda2ed74ed42ed19edd1ec8eec60ec24ecfeebfdebf5eb01ec28ec3bec53ec71ec74ec73ec79ec6cec62ec66ec57ec58ec6cec6fec8becc8ecf8ec3fed99edd4ed0fee47ee52ee56ee5dee4aee4dee6cee83eebdee18ef67efc9ef30f070f0aff0e7f0faf018f147f167f1a3f1f6f13df296f2f3f234f380f3d5f316f46cf4ccf415f561f5a6f5c0f5ccf5c8f5a8f597f598f59ef5caf516f65ff6b5f60af73ff769f782f77bf777f77df77df793f7bff7eef72cf874f8aef8e9f824f94af96ff99bf9b9f9dff90ffa36fa61fa96fac3faf8fa34fb63fb93fbc7fbebfb0cfc28fc2cfc28fc20fc07fceafbcefbabfb91fb83fb73fb73fb83fb94fbaefbc8fbd2fbd8fbd6fbc3fbadfb97fb82fb80fb8dfba5fbcdfbf5fb0ffc1ffc18fcf7fbc8fb89fb46fb0cfbd8fab1fa9efa8ffa84fa80fa77fa72fa7afa83fa9afac4faf3fa31fb80fbcffb2cfc96fcfefc77fdfcfd79fefdfe82fff1ff5f00ce002c01940108027b020803a3033304cd046205d00537069506d6062a079007f70789083709da09920a430bc90b540cd20c2a0d9c0d1b0e880e1d0fc10f4c10f3109f113012e612a813561435152016e816ca179b183219db19751ae61a841b311cd21cb21d9c1e621f43200621862117228d22d5224e23cc233224d3246f25dc256426ca26f9264d279427c2273328a72802298f29fc29272a5e2a632a2e2a232a0f2aef291e2a532a782acc2af72ae62ae22aa52a302adf297329f528b6286b280b28db278d271527b72637269d253025a324ff238323e02220228521c620fb1f5f1fa91ef11d6b1dca1c201c981be41a1c1a6f199618b317f5161b1643158f14b813d9120b120e110610120ff90dea0c020c050b160a4509550863077c067005670473036a027601a100c1fff6fe3ffe71fdadfcf5fb2afb73fad4f932f9aaf836f8b9f747f7cff63af6a6f50cf567f4dbf367f304f3cbf2a9f290f287f271f245f20ff2bef15cf103f1aff071f05ef061f082f0c5f006f145f17ef196f19af193f16ff14cf132f10ef1fcf001f100f110f130f145f167f191f1a8f1caf1f2f105f221f240f247f259f272f27af294f2bff2e4f225f37df3ccf329f488f4cdf414f556f57ef5b7f5fff53bf68ef6f4f64ef7b8f72af888f8eff857f9a7f9f9f944fa6bfa89fa9afa86fa6efa58fa32fa20fa28fa2ffa4cfa7afa95faa9faaffa89fa50fa0cfaacf955f913f9d1f8acf8a7f89af892f88bf866f837f805f8b9f76bf72af7dcf698f664f61df6d7f59ef556f51df5fff4e1f4d9f4f0f4fff40df518f5fbf4c6f487f428f4d0f398f36df36cf39df3d2f311f451f464f457f431f4d9f374f318f3b2f264f237f206f2e7f1d8f1b4f196f183f15bf13ef132f116f102f1f2f0c1f08bf054f003f0c7efaaef90ef9fefd4ef03f03cf072f07af073f063f035f018f018f018f03df07ef0aef0e6f01df12df140f15bf160f17cf1b1f1d9f111f24ef267f27cf28ff283f288f2a7f2c3f204f369f3c1f323f483f4b5f4daf4f7f4f3f4f9f416f529f552f58cf5aef5d1f5f2f5f2f5f5f504f605f618f640f658f671f68bf68bf68af694f697f6b5f6f9f647f7b1f72ff896f8eff833f946f93ef92af900f9e0f8d9f8def8fdf836f96ff9acf9e7f908fa1ffa2ffa2bfa25fa25fa23fa2bfa42fa5ffa8cfac4fafdfa3ffb82fbbbfbf1fb1efc39fc48fc45fc31fc13fce6fbb0fb7dfb49fb24fb18fb1afb34fb68fba0fbe1fb25fc52fc72fc88fc8bfc98fcbbfcecfc4efde4fd92fe66ff4d001e01e50194020f037b03dd032904900413059a054b061807dd07b9089a095b0a230be50b820c270dc90d4c0ee40e850f1410c61086113012f512ba135a140715a7151c16a0161f17811703188818f1187819f719501abc1a1a1b551bb11b101c611ce01c621dc81d451ea31eca1ef51eff1ee91e001f231f521fcb1f5920e32092211f227822cf22f322ea22fc22fe22f82225234b2363239423992372235123fc2283221d229521fa207a20dc1f2f1f9d1eef1d391da61cfa1b491bb21af51923195c1866176216771578148913cc120c126211db1038108c0fe20e040e160d2f0c2b0b360a68099808e9075c07c3063706b3050a055d04aa03d202f7011c0126003aff59fe6efd9dfcdffb20fb7bfadef931f98bf8d8f708f738f65ff578f4abf3ebf238f2abf12df1b9f05ff001f0a0ef4feff2ee93ee47eef2ed9bed53edfbeca1ec53ecf6eb9deb5aeb11ebd9eac0eaa5ea9feab6eac4eaddea02eb0aeb0deb0cebe9eac6eaadea8aea86eaabead8ea2deba1eb08ec77ece3ec22ed59ed87ed98edbdedfded40eeb1ee49efdeef8ff04bf1e7f185f21cf38df302f476f4c8f420f574f5a4f5d8f50ef62bf65ef6a7f6edf654f7d1f73bf8abf80ff942f964f977f965f960f971f981f9b4f904fa49fa96fadefafdfa11fb1efb0cfb03fb08fb01fb07fb1dfb1dfb22fb2cfb1ffb14fb12fbfbfae7fad9faaffa83fa5cfa1cfae0f9b5f97ef951f938f90bf9d8f8a4f849f8ddf770f7eaf66df610f6b8f57cf563f541f51df5fbf4b2f456f4f9f382f30cf3b3f259f210f2e0f19ff15bf120f1cef07ef046f00cf0e9efe7efe0efe0efe5efcaefa3ef7eef45ef1eef1fef30ef6aefd0ef36f0a6f014f15cf18ff1b0f1adf1a6f1a6f19df1a9f1cff1f6f135f286f2ccf218f360f38bf3aff3c7f3c4f3caf3daf3e9f319f463f4b0f414f579f5c6f50af638f644f64ff65bf668f69bf6eef653f7ddf770f8f4f871f9d4f911fa44fa69fa85fab8fafbfa46fbaafb10fc68fcbffc02fd2cfd52fd6dfd7ffd9bfdb7fdcdfdecfd03fe10fe23fe33fe44fe67fe95fec8fe09ff46ff77ff9fffb4ffb5ffb1ffa5ff97ff96ff99ffa1ffb3ffc4ffd3ffe5fff6ff080021003a0053006a00760077006e0058003f002c00200025003a0056007800930099008c006b003300faffc7ff9eff90ff9bffb1ffd9ff04002300440062007a00a400de001f017701da0130028b02de021f036b03c3031d049b042d05b8055206dd063f079607d807fb0732087c08cc084b09e309720a160baf0b1e0c920cfa0c430da70d150e6f0ee90e630fbb0f28109110e0105a11e81170122e13f7139d145315eb153f169616d916f9164e17c0173918fe18dd19a81a961b6a1cfc1c931d051e3f1e971eea1e251f991f142079201121a2211222ac22332391230b2464248324af24b0247a2463243a240024072415241c245b2483247e2485245024dc237123dd223022b4213321b52076202c20d81faa1f5d1ff81eac1e3a1eaf1d3d1da21cf21b5a1ba11ae3195019b1182118c4175717e6168216e71525155514461323121411f40ff30e280e600db10c1a0c590b830a990972083a070606c0049b039f02ac01e0002e006dffb8fe03fe32fd6afca6fbd1fa12fa59f997f8ecf746f799f607f67df5f1f481f413f49cf335f3c2f23df2c3f139f1a5f028f0a5ef27efc7ee65ee09eec7ed7eed3aed0cedd1ec96ec67ec1deccaeb7ceb12ebabea5dea0eeadfe9dfe9e8e910ea52ea81eaafeadbeadfeadceae0eaceead5eaffea2eeb86eb03ec7bec06ed98ed06ee70eed1ee0bef47ef87efafefe9ef34f072f0c9f035f196f10bf28bf2f2f25ef3c4f303f43ff476f48ff4b3f4e4f408f543f58ef5ccf519f66bf6a5f6e5f625f74af777f7aaf7c9f7f5f72cf856f88ef8d5f812f95ef9b9f906fa5dfab9fafafa38fb70fb8afb9efbb3fbb2fbb6fbc3fbc2fbc7fbd5fbd1fbd1fbd7fbcbfbc2fbc0fbacfb99fb88fb60fb2ffbfafaacfa5bfa14fac9f993f97ef974f97ef997f99af989f961f90af999f826f8adf74ef71ff70df724f75ef793f7c1f7e2f7d9f7b6f788f745f70af7e5f6c8f6c4f6d7f6e8f6fef617f71df720f725f71af710f70af7f5f6ddf6c5f69bf673f651f62cf615f60ef607f60af614f611f60df609f6f9f5eff5edf5eaf5f4f508f616f62df649f65bf677f69cf6c1f6f4f631f765f798f7c1f7d2f7d9f7daf7d3f7dff701f832f87bf8cdf80df93cf94bf92ff9fcf8bff882f865f870f89df8f1f857f9b2f9fbf923fa1cfafcf9cef9a1f991f9a9f9e7f94ffacffa4efbc6fb22fc55fc6efc6efc5efc56fc61fc82fcc2fc19fd7dfdecfd55feacfef8fe31ff56ff77ff94ffb1ffdcff120051009c00e7002c0169019201a601af01aa01a001a001a901c001e5010d023502570267026e02730275028c02c1020d037603f3036b04dd0438056f059605b605d3050e066e06e5067d072408b3082f098709aa09b909bd09ba09d9091c0a700ae50a610bbe0b0b0c340c2a0c170c010ce60bf30b220c5b0cb60c140d530d8e0dae0da40da10d9f0d970dba0df90d400eb00e2c0f960f12108010cd1027117811b51117128612f61295134114e01492152b169116ed161f172117301739173e177a17ca1718188618db18f9180219cd185b18f0177e171717fa16051728177a17b517bb17a5174717ac1616167915f614c314b914d01414153f153a151915af1412147513ce124112f911d211cd11f111fa11de11a61126117810c10ff30e350ea80d2d0dd20c9b0c540c000c9c0b010b470a7c098e08a607d70611066f05f20478040a049a0305035f02a801d4000b0056ffaefe33fed8fd83fd41fdf6fc89fc0dfc76fbc5fa21fa8af903f9aef875f847f82cf8fcf7a1f72ef78ef6cdf517f567f4d4f37ff349f329f322f300f3b8f256f2bff108f15cf0b2ef2aefe3eebfeec3eef1ee10ef1eef1befdeee7bee0fee8ded1dede0ecc2ecdbec30ed8aedeeed4bee6cee61ee38eedced7ded3eed14ed29ed85edf8ed8dee2def9aefe1efffefd7ef97ef5eef20ef0def31ef67efbdef22f05ef080f084f04af003f0c3ef7eef62ef77ef9defe3ef38f06ef09bf0b6f0a8f09ff0abf0bcf0fdf06ff1eff18cf234f3baf333f495f4c9f4f7f429f550f591f5edf547f6b5f62cf788f7e0f72ef856f875f88cf885f87df877f85ef852f855f851f85ff87cf88cf8a0f8b2f8a7f896f883f85ef844f83bf832f83ef85df873f890f8b1f8bef8cef8e5f8f4f812f942f96ff9a8f9e7f911fa32fa47fa3dfa2bfa19fafbf9eaf9e9f9e5f9e9f9f2f9e5f9d0f9b6f983f94ff91ef9dbf898f855f8f8f795f732f7c3f662f61bf6e2f5c7f5c6f5bef5b4f59cf559f5fdf494f41af4b3f374f359f375f3c4f329f49ff414f567f59ef5baf5aff59af58cf583f595f5c5f506f663f6cdf62bf786f7d4f702f81ff82df824f81bf816f811f81ef838f852f879f8a2f8bef8dcf8f4f801f916f931f94bf973f9a0f9c6f9edf90afa14fa1cfa1cfa18fa28fa4afa7efacffa31fb99fb05fc5efc9dfccbfcddfcddfce2fcedfc0efd51fdaafd16fe91fefefe5bffa6ffd2ffecff0500170039007300b30002015c01a601e8012102410262028a02b102f0024803a2030a047604c7040f05490568059005c70506066f06fd06980750080c09ab09410aba0a030b430b790ba00be50b420ca60c320dcb0d500edc0e4e0f890fb40fbc0f970f7e0f660f490f5f0f910fc90f2c109310dc102a11571151114b113011fe10f61004111b116f11da114012c6123d138c13e51324143e147414a714ce1423158015d1154616b016fb165b17a317ca170818391852188b18b618c418e918f118cf18bc188e1840181218da1796177f176117321727170617c4169c165d160716d915aa157c1589159e15b415fc153b166616ac16d416dc16f516ef16cf16cb16bc16a616bd16d316e7161f173f173e1740171217b5165a16da154a15dc146d140914d513a0136913471303139c122d128b11c9100c10390f690ec60d2f0db40c6c0c2a0cf20bcc0b890b2e0bcf0a460aa90916097808ea078807370708070807100726074807500746072d07e9068c062306a1051c05a3042904c403790333030003d50297024e02ea015a01ae00e7ff05ff29fe59fd9bfc09fc9bfb47fb15fbecfab9fa84fa38fad1f961f9e4f860f8eef785f727f7e4f6acf680f66cf65ef658f666f670f676f680f670f64af61cf6d5f588f546f508f5e3f4e2f4ebf407f536f552f563f56af552f52bf503f5c9f496f472f446f423f410f4f0f3dbf3d6f3cbf3cff3e9f3fdf31af43df445f443f439f410f4e8f3d0f3bbf3caf306f454f4bff43bf5a3f5fef54cf672f685f691f686f681f68bf68ef6a2f6c3f6daf6fcf628f745f767f78cf79af7a0f79bf775f745f711f7c9f690f674f665f67cf6b8f6fbf651f7abf7e5f70ff829f820f814f811f80cf822f855f88bf8d5f82bf96ff9b0f9f1f91cfa46fa72fa8efaa9fac3fac3fabefab5fa96fa79fa6cfa5cfa59fa68fa6dfa71fa6dfa46fa0afabef954f9eaf88df82df8e5f7b7f788f761f73ff709f7d2f69ff65ff631f619f601f6fcf509f609f60ef619f615f618f625f629f638f64ff655f65cf665f65af651f652f64cf655f66ff680f699f6b1f6aaf694f66ef628f6e1f5a4f56af551f55cf573f5a1f5d6f5f2f5fef5f2f5bdf57af531f5ddf4a1f482f473f48df4c5f40af568f5cdf524f67df6c9f6f7f61ef73af744f75df784f7b5f70bf87af8f4f884f916fa92fa03fb59fb8afba9fbb5fbaefbaffbb7fbc4fbe7fb15fc44fc7efcb3fcdefc0dfd38fd5bfd85fdadfdccfde8fdf7fdfbfd00fe01fe09fe29fe5cfea7fe0eff80fff7ff6f00d400260165018c01a801c701e70118026102b50219038603ec034d04a504ed0432057105a705e0051906460672069806b306cf06eb06060731076707a207f10747089708ea082d0957097409730954092d09fb08c808ad08a508b508ee0839098709df091f0a390a3a0a100abf096a091209c408a508ab08d3082a098a09e0092d0a530a490a270ae5098f0948090709d008b808aa089e08a308a108950895088f088208860885087f0885087f086a0859083e081e08130810081b084a088508c1080d094c0973099309990989097a095f09400934092a09230936094a095b0977098b09900995098709680948091809dd08ab08730836080908db07ac0787075f0735071007e406b6068f0660062e060006ca058c054f050a05c5048a0452042a0417040d0411042004280427041b04f703c60388033c03f302af027002430222020602f701ea01d201b30183013b01e5007900f7ff73ffe5fe51feccfd50fddffc87fc3bfcf9fbc6fb8afb42fbf5fa8efa13fa99f914f992f82af8cef78af76bf758f756f76bf776f778f779f759f724f7e8f68ff62df6daf583f53bf515f5f7f4eef401f50bf513f51ff50bf5e5f4b9f471f423f4e4f39df367f34df332f329f335f336f340f355f356f358f361f351f33ef32df302f3daf2bdf293f27cf27df279f28cf2b4f2ccf2ecf215f328f33ff35af35ff36af37cf377f379f384f37ef387f3a1f3b3f3dcf31df455f49bf4e9f41cf549f569f564f559f54cf52cf520f52af535f55af597f5ccf50df655f689f6bff6f1f604f712f71af701f7e7f6d0f6adf69df6a6f6b4f6e3f62cf771f7c4f716f849f86ff882f870f856f83df81af810f823f83df873f8c1f808f956f9a5f9dbf90bfa36fa45fa4bfa4bfa32fa17fa01fae1f9d4f9e3f9fef936fa89fadefa38fb8cfbc1fbe0fbeafbcefba6fb7efb50fb36fb39fb4bfb79fbbbfbf8fb38fc6efc85fc89fc80fc5cfc30fc02fccafb9cfb7afb58fb46fb47fb4afb57fb69fb6dfb6bfb62fb43fb20fbfffad9fabffab2faa6faa2faa3fa9afa8ffa83fa72fa6afa72fa87fab2faf0fa35fb7dfbbbfbe2fbf6fbf6fbe7fbdafbd9fbf1fb28fc7bfce5fc60fdd9fd45fea1fee3fe0eff26ff2cff2aff29ff27ff2fff45ff63ff90ffcdff0e0052009600ca00f10007010201ec00cc00a1007d00680062007900ac00ee004701ac0108026002ad02e3020e032c03370347035c036f039a03da0323048b0405057d05fc057006c306070732073a07450751075a078307c20706086708d1082d099109ee09340a820aca0afe0a420b830bac0be00b0d0c210c400c5f0c700c9e0cd90c100d670dc50d120e6e0ebb0ee40e0f0f260f1a0f1c0f1a0f0b0f210f460f710fcd0f37109c1022119b11ed113f126e1267125d123b120112eb11e311e2111f127312c7124213b4130014501479146f1467144214fc13d513b11388139513b513dc133a149e14f2145e15a915bc15c21594152c15cc145f14ec13b813a413a913ef133e148114d514ff14f114dc149c143414e01385132813fd12de12c712e112fa120b133b135913571362134c130f13d71281121612cc11821143113b1140114b1173118611781168113011d7108b103610e40fbb0f9c0f830f870f790f540f310fed0e900e400ee50d8d0d540d1d0dec0cce0ca00c640c2d0cdb0b750b160ba50a2f0ac8095909f208a90866083408230815080c080a08ee07bb0776070d078f0616069a053305f304cd04cc04ec040f0532054b0541051705d0046604ec036e03ec027d022602df01b401a30199019c019c01870162011d01ab001f0078ffbafe06fe5ffdcefc6afc25fcf8fbe5fbd2fbacfb7afb28fbb2fa2ffa9bf900f97af802f89df75df72ff711f70af702f7f9f6fbf6f0f6ddf6cdf6aef686f660f62af6eff5bef584f550f531f512f501f506f508f510f524f520f50ff5f6f4b7f466f412f4a7f343f3fdf2c2f2acf2c3f2e1f212f354f377f386f384f354f315f3d8f288f24bf231f21ef228f252f276f2a7f2e5f209f32ef359f369f37af392f38ef38ef396f38bf38ff3aaf3c3f3fcf353f4a3f403f56bf5adf5ddf5fbf5e8f5cbf5a9f573f553f551f54ff570f5b0f5e5f529f674f69ff6c3f6daf6cbf6b5f69cf66bf64af643f63bf657f695f6d2f61ff774f7a7f7c8f7d4f7b1f782f74ef709f7dbf6cdf6c5f6d9f605f725f745f760f75ef756f74cf72ff71cf714f7fff6f4f6f1f6dff6d3f6d3f6cdf6d6f6f1f607f728f74af753f74ff73df70bf7d4f6a6f678f666f679f69cf6d5f61df752f777f787f76df73ef70af7caf69bf68ff695f6b7f6f6f634f770f7a3f7b4f7acf792f75bf71bf7e4f6b0f692f694f6a6f6cdf606f737f75ff77bf778f760f73af702f7cdf6a8f68ef691f6b4f6e9f633f789f7d6f71ef858f876f884f888f87df877f87ef88ff8baf800f953f9b9f926fa86fadcfa20fb42fb50fb4ffb41fb38fb3efb51fb7dfbbffb09fc5bfcaafce6fc13fd2cfd2ffd27fd1afd0bfd07fd12fd2bfd58fd92fdd2fd1afe61fea2feddfe0bff2eff4eff68ff83ffa9ffdaff1d007500d5003a01a101f8013f0275029402a802bd02d302f7022f037103bf030f044e047c0497049504860473045f045b0467047e04a104c704e104f504fb04f004e504da04cd04cc04d104d604e204eb04ee04f604fc0404051a05360555057f05a405bc05d005d605d005ce05cd05d305f005170644067d06ad06cd06e306e306cb06ae0686065a0639061e06080603060006fe0508060b060506fd05e505b70580053805e804a20465043f043d0451047804af04dc04f204ef04c20472041404aa0348030403de02dd02ff022b0358037e03830367033403e5028a023202e0019f0177015d0155015e01640169016c015d0143011c01e400a60064001c00ddffabff82ff6dff66ff63ff67ff65ff52ff36ff0affd1fe9afe65fe35fe18fe07fef9fdf5fdedfddbfdc3fd9efd6dfd3efd0cfddbfcb6fc95fc76fc64fc4efc33fc1bfcf7fbcafb9dfb60fb1bfbd9fa91fa4dfa1dfaf6f9e1f9e7f9f2f9fff90efa05fae7f9bcf974f922f9daf892f85df84cf84bf85ff88cf8b0f8ccf8e4f8daf8b7f88cf843f8f3f7aff766f72bf70ff7fcf6fff620f73df761f78bf797f78cf76ff727f7ccf66ef603f6abf579f559f55ef587f5aef5dbf505f608f6f6f5d2f58bf541f5fff4b8f489f477f46bf479f4a0f4c2f4f3f42af54bf568f57df56df552f531f5f9f4ccf4b1f497f49bf4bdf4ddf407f533f53cf533f51bf5e2f4a9f47ef455f448f458f466f47df496f492f482f46bf441f422f41bf41df43cf474f4a7f4dcf409f513f50ef501f5e1f4cff4d4f4e1f40bf54bf584f5c3f500f624f647f66af67ff69ef6c7f6e5f607f729f738f74af760f770f792f7caf706f853f8a8f8e8f81bf93cf938f925f90ff9f2f8e9f8f8f813f947f98ef9ccf90afa45fa6efa90faaefabffad2fae8faf5fa08fb21fb38fb5efb96fbd8fb2efc91fcf2fc4cfd90fdaffdb3fd9bfd6ffd4bfd3cfd47fd7cfdd2fd38fea4fefdfe34ff4cff41ff1efffcfee6fee4fe06ff42ff91ffecff3e008400be00e300fd0017012e014b0172019901c601f701220252028702b902f3022f035e038903a803ae03ad03a903a303b603e00318046c04cb0417055a05820583057a056a0552055a058105b90515067e06da063a078907b407dc07fc070b082a0855087d08bd0803093f098c09da091a0a6f0ac80a150b6e0bbe0bf20b240c430c460c570c6b0c7c0cb10cf60c380d8f0dde0d120e480e670e660e6d0e690e520e510e4d0e3f0e4b0e570e5e0e860eb20ed70e140f4a0f670f8a0f920f790f6d0f590f3d0f4b0f690f920fe40f36107510bc10e810ed10f410e810ca10c810c510bb10d110e210e010f110f510e910f6100011fe1016111f110e110711e710ad1088105f103610351039103b105a106710571050103010f70fd50fae0f860f830f7e0f6f0f780f6e0f4d0f400f290f090f0e0f170f1d0f3d0f4b0f410f420f290ffa0ee70ed30ec00ed40ee60eeb0eff0ef80ed00eb00e7d0e3f0e250e0f0efb0d060e050eeb0dd60da70d5b0d200de10ca40c910c870c7d0c8f0c930c7f0c730c530c1f0c040ce80bcb0bd10bd50bcf0bdc0bda0bca0bcf0bd10bd40bfb0b210c3d0c640c6e0c540c360cff0bbd0b9c0b8a0b8d0bbb0bed0b140c3b0c3a0c0e0cd80b880b2f0bf30ac60aac0ab60ac10ac20ac40aa90a750a440a0b0ad609be09ab099e09a009900969093d09fe08b6087f0851083608390840084808530846082208f907c0077e0746070b07d606aa0674063c060706c505840552052005f404d204a5046e042904c9035d03ed0276021002c401870164015501440137012101f700c400890042000400c8ff82ff43fffffeaefe62fe16fecffda1fd84fd70fd6dfd60fd3bfd01fd9efc14fc7dfbd7fa38fabdf95ef923f912f909f900f9f4f8c5f878f818f896f707f783f6fdf584f52af5d9f49cf47cf45af442f440f434f426f421f405f4ddf3b9f380f346f322f3fcf2eaf2fef218f341f380f3aef3d5f3fbf302f4fdf3fbf3def3bcf3a6f37af34ff332f309f3edf2ecf2e5f2eef20cf314f31af31df3f7f2c5f293f246f207f2e5f1c0f1b8f1d1f1e1f101f22af233f23ff250f243f240f24df247f252f269f268f26ff27ef274f279f291f29cf2bef2f1f211f336f35af35df35ff360f347f339f338f328f325f32cf323f321f323f313f30ef317f317f327f344f352f364f371f364f353f341f321f313f321f33bf37bf3daf33cf4aef422f57bf5cdf512f639f660f68cf6aef6e4f62cf773f7d1f73ff8a4f813f981f9d4f91dfa52fa5bfa50fa34fafef9d1f9b2f996f998f9b2f9d0f9f9f91bfa21fa17faf6f9b2f968f922f9ddf8b1f8a3f8a6f8c2f8e8f805f91df929f91ef909f9f1f8d5f8c4f8c1f8c8f8def801f926f955f98af9b8f9e3f909fa22fa31fa32fa26fa1dfa1bfa1efa37fa6afaa9faf5fa43fb7ffba6fbaefb8efb56fb11fbc6fa93fa82fa91faccfa2afb93fb00fc62fca5fcd0fce2fcddfcd7fcd9fce6fc10fd53fda4fd09fe7cfef0fe67ffdaff3e009600d900010113010e01f300cf00ac00900088009500b400e6001e014f0172017b0166013601f0009c004a000200cdffb1ffadffbbffd8fffcff23004a006e008a009f00ab00b000ae00a700a400aa00bd00e2001b016101b20107025902a402e40217034003610377038c039e03a703a803a30394037e036703510349034e035c0374038e039c03970378033b03e80287022202cd0195017b018301a501d601100244026a0284028e02860276025f02420225020902f301ea01ed01fd011e024b027b02aa02ca02d102c0028f023f02dd0172010801b0006f00490043004f0064007c008b00890076004c001200d2ff8dff48ff0cffe0fec7fec8fee1fe0dff4bff91ffd3ff0c003100410042003500220018001d0032005b009400d7001a0156018801ad01c301ce01d001ca01be01ad019601770149011001d000890042000200c7ff90ff5fff2bfff1feb1fe67fe16fec7fd77fd2dfdedfcb1fc7dfc52fc2afc07fcf3fbedfbf6fb15fc3ffc70fca4fccafcdffce2fccffcaefc8dfc70fc63fc74fc9cfcdafc2cfd82fdd3fd15fe3cfe4bfe46fe2cfe05fedffdb8fd9afd8efd8ffda2fdc8fdf8fd2ffe66fe8bfe9cfe96fe6cfe2afedefd89fd43fd1bfd0cfd20fd54fd90fdd1fd0afe25fe2cfe1ffef7fdccfda8fd88fd7bfd7ffd87fd97fdaafdadfdaafda0fd85fd65fd41fd12fde4fcb5fc7afc3efc05fcc8fb90fb62fb35fb11fbeffac4fa96fa67fa2ffafdf9d7f9bdf9b8f9c6f9def9fef91ffa35fa40fa40fa34fa2bfa2cfa34fa4efa7dfabafa06fb59fba8fbfbfb49fc89fcc3fcf4fc15fd2efd3dfd3cfd3cfd3efd41fd58fd86fdc2fd13fe6cfeb4fee9fefefee1fe9efe3dfec5fd58fd04fdccfcc5fcebfc2dfd83fdd9fd19fe3ffe43fe1efedffd91fd39fdeefcbdfca9fcbafcecfc38fd96fdf9fd55fea3fed9fef3fef2fed9feb3fe88fe61fe4bfe4afe5cfe81feb3feeafe23ff58ff83ffa6ffc1ffd0ffd4ffd1ffbfffa1ff7bff4eff26ff0eff09ff22ff5cffadff0d007400ca00040123011e01fc00cd009e0081008600ab00f3005f01d8015602d2023b039103d303fb03150425042b04300438043f04500469048304a804d5040305380568058805a305ab059705770548050805cd0494045f04450440044b047904bc0406056205ba05fd05360654064e063e0622060006f7050806340691061107a2074c08f4088109f609410a570a4e0a290aed09bf09a2099a09c0090a0a6a0ae50a620bc70b160c380c1e0cda0b6e0be00a570adb0978094d094e096b09ad09f309200a3c0a2f0af509aa094909df0893085d083d084d087308a008e008150936095809660963096f0978097e099709ab09b309c309c009a90998097a095409420932092509350949095a0977098309770965093909f208af0866082208fc07e907ec0715084a088008c408f908140923091809f408cd089d086c085308450846086c089f08d80826097009ab09de09f209e509c40982092709cf0871081c08eb07ce07c407da07f207ff070608e807a6074c07d0064206c1054605e104a804870480049704b004c604e004e404d704c804a904870471045c045404630473048604a804c204d304e804f50403051805280538054e05570553054a052c05fc04c9048b0449041204e503c903c303c603ce03d903d303b8038c034703f10297023b02e701a70177015b015701600175019601b301ca01db01dc01d201bf019f017c015c013c0125011e012201380160018f01c401f701170223021702e801a0014801e30082003000edffc6ffb9ffbfffd5fff1ff01000100eaffb1ff61fffdfe90fe2bfed7fd9bfd7ffd84fd9efdc9fdfbfd28fe4bfe59fe51fe37fe0ffeddfdacfd82fd65fd59fd5afd65fd79fd8dfd9ffdaafda8fd99fd80fd58fd27fdf6fcc0fc8dfc62fc3bfc18fcfcfbdcfbbcfb9afb6dfb3efb12fbe4fabbfa9dfa83fa6efa61fa4ffa3bfa26fa0afaeaf9d0f9b8f9acf9b5f9cbf9f3f92ffa71fab4faf8fa30fb59fb76fb7ffb7afb72fb66fb62fb6cfb85fbb1fbf0fb36fc7efcc6fcfdfc20fd2dfd20fd01fdd4fc9cfc6cfc49fc34fc37fc54fc80fcb9fcfbfc31fd5afd6ffd67fd48fd16fdcffc86fc46fc0cfcebfbedfb06fc3afc83fcc9fc05fd31fd35fd19fde6fc95fc39fce5fb97fb64fb57fb63fb8cfbcefb0ffc44fc6cfc71fc55fc22fcd4fb7bfb2cfbe5fab3faa3faadfad0fa0bfb4dfb8ffbcefbf8fb0dfc10fcfcfbdefbc5fbb1fbaefbc2fbe6fb19fc5bfc9afcd4fc09fd2cfd41fd50fd4efd47fd45fd40fd3ffd46fd46fd48fd4bfd41fd37fd34fd2afd27fd30fd33fd39fd40fd36fd22fd08fdd8fca1fc6afc26fcecfbc6fba3fb91fb98fba2fbb4fbc9fbc8fbb9fb9cfb64fb1efbd7fa8bfa4cfa26fa0ffa12fa32fa58fa83faaffac8fad0fac8faaafa83fa5cfa33fa15fa0afa08fa17fa39fa60fa8efac2faeffa1afb40fb57fb65fb68fb5bfb4cfb3ffb2ffb2ffb43fb65fb9dfbe8fb33fc82fccafcf7fc12fd18fd00fde1fcbffc99fc84fc86fc93fcb8fcedfc22fd5cfd94fdb6fdcffdd9fdcefdbcfda4fd82fd69fd59fd4efd55fd69fd84fdadfddffd10fe45fe76fe9bfebafec8fec4feb5fe9cfe79fe58fe3dfe30fe3bfe5cfe92fedffe36ff88ffcaffedffedffcaff86ff30ffdcfe97fe70fe74fea2fef4fe63ffdbff4a00a200d600e200ca0094004d000700ccffa8ffa8ffc9ff06005d00c3002a018c01de01120228021c02f201b40167011b01e400c800ca00f10036018b01e4013002650277025c021902b9014101c3004e00eeffabff8cff90ffafffdeff110040005d005b003e000400b3ff54fff6fea6fe70fe58fe62fe8dfed0fe22ff78ffc5ff06003600510058004e0037001a00fbffdfffd0ffd2ffe7ff16005d00b40014017201c101f7010502eb01b0015b01fe00aa006d0053005e008600c40007013e015c0156012c01e6008b002900d1ff8fff67ff59ff60ff76ff92ffa8ffb1ffb1ffa6ff92ff7dff6bff5fff59ff59ff5aff57ff4dff38ff19fff2fec6fe9dfe81fe73fe77fe8efeb2fedafefcfe0dff05ffe5feadfe65fe1cfedefdb4fdaafdbdfdedfd33fe80fec9fe06ff2cff3aff36ff23ff0bfff7feebfeecfefafe10ff33ff5fff91ffcdff110057009e00e100150136013a012001f400b70073003c001b0014002d005f009e00e00014012b012401f4009f003500c0ff48ffdffe90fe5efe4dfe58fe78fea8fedafe00ff18ff1dff0affe0fea6fe62fe1efee4fdbafda6fdacfdcbfd00fe46fe90fed8fe17ff46ff60ff62ff4cff22ffecfeaffe77fe4efe3dfe49fe74feb7fe0fff6fffc8ff0f00380040002800f3ffadff69ff30ff0bff07ff20ff54ff9ffff4ff48009600d100f50006010201e900c4009600630035001000f7fff9ff16004b009500ed0043018b01b501b80194014901df006a00f8ff96ff51ff34ff3cff61ff97ffd2ff050020001900f2ffb2ff5dfffefea2fe55fe1ffe02fe00fe1afe48fe85fecbfe11ff50ff86ffaaffc1ffcbffc6ffb8ffa8ff97ff8aff87ff8effa6ffd2ff0f005f00c10029018f01e9012b024e024e022802e8019d0152011a01060119015801be013902b70224036c0382036403110399020c027c010001a60077007a00a800f5005601b9010b0241024f023102ec01890111019a003300ebffd2ffe6ff23008300f8006c01d101170233022602f00199013701d10073003300180021005300ab001b01990113027c02cb02f202e902bf0278021a02bf017901510158019001ef016a02ed026103bf03f303f303cc0387032b03cf028102480232023f026802ac0201035c03ba030b044304690473045b042d04ee03a3035f032803030301031c034d039603e0031a04450450043304fe03b30359030403b8027c025f025d027002a102df021e0362039a03b803c403b6038e035c032103e702c302b002af02ca02f3021f034f0377039003a103a5039e039a0394038d038e038e038a038a03880386039103a303bf03ea03190444046d0485048604780457042704f703c8039f0387037b0375037c0386038d039b03a703ae03bb03c203be03b903a803870362033a031103f702e902eb020b03370366039c03c803df03e503d103a4036c032703dc02a0026d02490241024c0267029602c602f4021d03300327030a03d20289024002fa01c601b201b601d4010d024c028a02c202e502ef02e802cb029c0265022702eb01bd01990188019401b501e80130027d02c002f5020d030203d7028e023402de0192015d014e015c017f01b201e40104020f02fe01d5019d0159011301d5009a0066003f001f000700feff02001500370063009500c900f00008010e01fd00da00af0080005a0047004b006a00a100e50031017a01b701de01ec01dc01b40177012d01df009c006f005d0068008e00c300fd002d01460143012201e40091003600ddff8fff51ff24ff07fff8feedfee5fee0fed9fed4fed2fed2fed3fecdfebafe98fe68fe2afeeafdb3fd8ffd89fda1fdd6fd20fe72febefef2fe06fff8fecefe8dfe44fe01fed1fdbcfdc5fde6fd1cfe5afe99fed1fefafe11ff17ff0ffffcfee5feccfeb7feacfeacfebafed3fef3fe1aff44ff6bff8dffa8ffb8ffc0ffc2ffbcffb5ffa9ff98ff88ff77ff67ff5fff5fff6aff83ffa6ffccfff2ff0a000e00ffffd7ff9bff57ff15ffe1fec2feb9fec7fee6fe08ff21ff2eff29ff0fffe5feb6fe8cfe6ffe61fe61fe6efe83fe9afeadfebdfec7fecdfed2fed4fed6fed9fedcfeddfedffee0fee2fee4fee5fee9fef0fef4fef7fefafefbfefbfefefe01ff0dff22ff3aff54ff6dff7dff85ff83ff76ff66ff59ff4dff48ff4cff55ff63ff70ff76ff79ff79ff70ff67ff63ff5dff59ff58ff55ff53ff4fff47ff41ff42ff46ff51ff64ff78ff8aff99ff9cff92ff7fff62ff3eff18fff0fecafeacfe90fe7bfe6ffe63fe5bfe59fe54fe50fe4bfe3efe29fe0bfee1fdb5fd8dfd68fd55fd59fd6dfd92fdc0fde6fd02fe0efe03fee5fdb9fd84fd57fd3afd27fd28fd3dfd5bfd7efd9ffdb6fdc6fdd0fdd0fdcefdd1fdd5fddffdeefdfdfd0ffe24fe36fe46fe57fe64fe72fe81fe8afe91fe98fe9afe99fe95fe89fe78fe62fe42fe1ffefefdddfdc3fdb9fdb9fdc5fddcfdf4fd08fe13fe0afef2fdcefda0fd74fd55fd42fd43fd5afd7cfda4fdcdfde9fdf6fdf3fddafdb9fd96fd6ffd51fd42fd3bfd41fd54fd68fd82fda1fdbbfdd4fdeffd00fe0ffe1afe1bfe19fe1afe18fe1bfe28fe35fe47fe5ffe6ffe79fe7dfe71fe5dfe44fe1efef5fdcffda5fd82fd6bfd55fd47fd44fd44fd4afd55fd5afd5dfd5cfd50fd3efd29fd0efdfbfcf3fcf3fcfefc14fd28fd3cfd46fd3dfd25fd03fdd6fcaafc86fc69fc60fc6bfc7dfc97fcb6fccbfcd9fce1fcdbfcd1fcc9fcc0fcc2fcd0fce0fcf8fc17fd2ffd41fd50fd4ffd44fd33fd18fdfcfce4fcc8fcb2fca6fc97fc8cfc89fc82fc7bfc7afc75fc70fc74fc77fc81fc94fca4fcb5fcc6fcc9fcc5fcbefcabfc98fc8cfc83fc85fc94fca2fcb2fcc1fcc0fcb4fc99fc6afc39fc0cfce3fbccfbcffbe5fb0ffc46fc79fcacfcd2fcdefcdafccafcaafc88fc6efc5afc58fc69fc84fcacfcdafc01fd21fd35fd34fd27fd12fdeffccdfcb3fca1fc9cfcabfcc6fceefc1dfd46fd6dfd8efd9efda3fda4fd9dfd94fd8ffd8afd8dfd97fda3fdb5fdccfdddfdeefd01fe0efe1bfe28fe31fe3bfe46fe4cfe53fe5cfe64fe72fe84fe97feb1fed3fef3fe13ff34ff54ff71ff85ff90ff98ff9aff91ff86ff7dff74ff6fff6eff71ff7bff89ff95ffa2ffadffb1ffaeffa2ff8cff73ff59ff3eff28ff1eff1eff2bff40ff5bff7aff97ffadffbeffc6ffc2ffb8ffabff9fff97ff98ffa2ffb6ffd3fff9ff24004d0070008e00a300ae00b000ac00a700a500a800b300c600df00020129014a01680181018e0191018c017e01710165015c015b015f01640170017d0185018c0190018e018b0185017e017c017c017e018a019701a301b201c001c701d001d301d101d301d401d301db01e801f90111022602370247024e02490241023502290228022e023b02550274029502b902d202e002e802e202d102c002ad029e029b02a102ac02c202d702e802fb0208030b030903fe02ec02e102d502c802c802d202de02f5020f0325033c034a034e0355035303460340033a033203340339033b034303470345034803470342034a03570365037f039903ac03c403d403d603d603d003c303bf03be03c003d403ec03030421043a0445044a04400427040c04ec03c803b103a503a303b803d703fc032c0454046e04810482046e04550433040d04f403e203d803e403f8030f042c043d043d04390429040a04e903c603a3038f038203780380039103a403c503e503ff031d0433043b043f043a042a041d040e04fd03f803fb0302041504270432043f04440439042e041f040a04fa03ed03e003e003e703ed03fa0305040904120418041504160416041104110412040a040404f903e603d603c103a2038c0379036503600365036c0380039503a003a903a7039503810368034d0341033e0342035c037e039e03bf03d403d603cd03b3038b036603450328031e031d03220332033e033e033b0330031d030c03fa02e902e602e902ef02000312031e032b0330032b03240319030b03070307030b031a032c033e0351035a03560349032f030c03e802c402a30295029802ab02ce02f7021e0341035303500340031f03f302ca02a6028c0286029102a702c902ec02070319031a030503e302b10276023f021002eb01dc01e101f501190243026b028c029e029d02900276025102300219020b020d021a022f024b02620270027602700260024d02340219020202ec01d801cd01c301b801b401b301b501b901c001cc01de01eb01f201f501ef01df01ca01af0194017c0169015c01570156015c01650169016901660158013f011f01fa00d700b700a100970098009f00ae00c000cd00d400d300c800b3009700760057003b00230010000000f4ffecffe3ffd8ffceffc7ffbeffb5ffaeffa5ff98ff87ff74ff63ff52ff43ff3dff3eff46ff54ff65ff75ff82ff87ff87ff81ff75ff66ff58ff4cff43ff3fff3eff3dff3fff40ff3eff3cff37ff32ff30ff2cff28ff25ff21ff18ff0dff00fff3fee7fedafed0fecdfecbfec9fecbfecefecefecbfec3feb7fea9fe95fe7cfe66fe52fe41fe3afe38fe3bfe44fe4efe55fe58fe51fe41fe2ffe18fe01feeffde1fddcfde3fdebfdf1fdfafdfcfdf6fdecfddbfdc8fdbafdaffdaafdaffdb6fdbffdccfdcffdccfdc6fdb9fda7fd98fd8afd84fd88fd90fda0fdb4fdc1fdccfdd6fdd2fdc2fdaffd98fd82fd70fd5ffd5afd62fd6dfd7dfd91fd9cfd9efd98fd84fd68fd48fd24fd06fdf3fce6fce4fceefcf8fc05fd10fd10fd06fdf7fcdcfcbefca2fc87fc74fc6cfc67fc67fc6dfc6ffc71fc74fc70fc6bfc68fc5dfc54fc51fc4dfc4bfc4cfc4cfc4dfc50fc4bfc46fc44fc3cfc34fc2ffc27fc20fc1efc19fc16fc17fc13fc0efc0cfc03fcf9fbf4fbe9fbe3fbe5fbe6fbebfbf5fbfbfb02fc0bfc09fc04fc00fcf4fbe8fbdefbd0fbc6fbc2fbb8fbaffbadfba7fba3fba5fba3fba2fba5fb9ffb99fb93fb85fb79fb75fb6cfb68fb6bfb6ffb7dfb90fb9afba5fbb1fbb2fbaffba9fb99fb8afb80fb75fb6ffb70fb6efb74fb80fb88fb93fba1fba6fbaafbb1fbb0fbaffbb0fbadfbadfbb2fbb5fbc0fbd1fbdefbeffb04fc11fc19fc1dfc1bfc19fc14fc09fc01fcfefbf9fbf8fbfefb02fc0bfc1bfc28fc37fc49fc57fc65fc73fc7afc82fc8bfc8afc88fc8cfc8ffc96fca3fcb0fcc2fcdafcecfcfafc04fd03fdfffcf7fce3fccdfcbdfcabfc9ffc9dfc9efca9fcbdfcd2fce9fc00fd0efd17fd1bfd12fd04fdf7fce7fcdcfcddfce6fcfafc1bfd3efd64fd88fd9efdaafdadfda1fd8dfd79fd66fd59fd57fd5ffd74fd95fdb9fddffd07fe28fe41fe53fe58fe57fe53fe4cfe49fe4ffe5cfe72fe8efeadfecffeeffe03ff0cff0eff08fffcfeeefee2fedafed8fedefeeafef9fe08ff15ff23ff2fff38ff3fff4bff5cff70ff84ff99ffacffbcffc4ffc7ffc6ffc1ffbeffbdffbcffc1ffcbffd4ffddffe6ffe9ffe7ffe0ffd3ffc3ffb5ffa9ffa3ffa6ffafffc1ffdbfff8ff1600330049005900610060005d005a00570059006200710083009900ab00b900c200c400bf00b800b100af00b500c500dc00fa001a01380154016701710175017401740178017b017f018c019e01b001c101cc01d201d001c301af019a0180016701580150014f015c0174019201b301cf01e601f601f601ea01dd01cd01c001be01c501d501f0010e0228023e02470246023f022c021302fd01ea01db01d701d801db01e401ec01f301fb01fe01fd01ff01fe01fd01020207020b0215021c021f0221021d02160211020902000201020602100225023d0253026a0276027702710260024b023b023102330249026a029402c502f20217032f03330329031603f702d502bf02b302b302c302dc02fb021c033803490350034b033c0325030803ee02dd02d002cb02d602ec02040320033b035203610363035c0355034b033b0330032a0325032503250321031f0319030f030803ff02f802f602f402ef02f102ee02e102d402c102a90297028a0284028d029d02b502d702f5020a031b031f0315030503ea02c902ad029502870289029602b002d8020203270349035c035c034e0333031003f002d502c602cd02e10201032b03550377038f0391037f03620338030703d902b2029602880284028a029a02ab02b902c602ce02cf02c902b802a00288026e02540241023702340238024302520263026f02740275026d025d0246022b020d02f201dd01ce01c801c901d301e401fa010f0226023502390237022a021202f801de01c701bb01b601b801c401d501e401f001f301ee01e401d301bf01b001a3019b019e01a401ad01ba01c201c701cf01d201d101d301d101cd01cd01c901c201bc01b101a7019e0193018a018801850185018801890189018d0191019401970197019901990192018b0185017a017001680162015d01590154014f0148013c012e01210111010101f600ed00e500df00db00d800d500d200cd00ca00cb00ce00d200d300d300d600d500cf00c800c000b400a7009b009100890081007b007a007a007e00860090009d00ac00b700bc00ba00af009c008700710060005b00610072008e00aa00c300d500d900cb00af00870056002400f7ffd7ffcbffd0ffe4ff020025004900630068005e0047002200f5ffc7ff9eff82ff78ff7dff94ffb5ffd9fffaff110016000900ecffc4ff97ff6aff43ff2bff1eff1dff28ff36ff44ff53ff5eff62ff62ff60ff59ff52ff4aff40ff35ff2aff20ff17ff0fff0dff14ff21ff32ff4aff62ff73ff7cff7bff6dff52ff2eff09ffe7fec8feb3feaefeb4fec3fedcfefbfe1bff36ff46ff4aff3eff22fffdfed7feb3fe95fe87fe88fe99feb4fed3fef1fe08ff11ff0cfff6fed0fea4fe77fe4efe32fe28fe2afe38fe50fe6cfe88fea2feb6fec5fed0fed7fedafed9fed3fecdfec7febdfeb6feb5feb6febafec5fed1fedafee1fee3fedffed4febffea4fe8afe6dfe50fe39fe29fe22fe27fe37fe50fe70fe8ffeacfec2fecbfec9febcfea2fe7ffe60fe44fe31fe2efe39fe51fe72fe91fea9feb7feb6fea8fe91fe73fe5afe4dfe47fe4efe65fe83fea8feccfee8fe01ff14ff18ff18ff12ff04fff9fef2fee8fee5fee7fee4fee4fee5fee1feddfed7fecbfec3febdfeb7feb9febffec5fed4fee3feeffefcfe02ff00fffffefcfef6fef7fe00ff0cff1eff31ff3dff44ff46ff3dff2fff1eff0cfffefef3feeafee7fee6fee6fee9feecfeeffef4fefafefefe05ff0bff0eff13ff16ff12ff0cff08ff01fffbfef8fef7fefdfe09ff14ff20ff2cff30ff32ff31ff2bff27ff24ff1aff10ff08ff00ff00ff02ff07ff1bff38ff53ff6fff87ff94ff9aff96ff85ff72ff5cff45ff38ff31ff30ff3dff51ff68ff84ff9dffadffb6ffb6ffa9ff95ff78ff57ff39ff1fff0cff0bff1bff39ff65ff99ffcafff2ff0a000d00faffd5ffa8ff7aff53ff3dff3cff4cff6bff94ffbcffdcfff1fff6ffeeffd9ffb8ff92ff6fff53ff40ff36ff38ff42ff54ff6cff85ff9bffafffc0ffc8ffcaffc8ffbcffa6ff8fff7aff66ff58ff52ff54ff5dff6dff82ff9cffb7ffd2ffe7fff5fff9ffeeffd7ffb8ff96ff77ff64ff60ff72ff9cffd2ff0d00470073008d008d00740048001400ddffb2ff9aff97ffacffd5ff07003a00680085008e008400680046002100ffffe4ffd6ffd3ffdcffefff070020003600470050004c003f002b001300fcffe9ffdcffd8ffdfffebfffaff0600100018001b001d00220026002b00320038003b003a003200260018000700f8fff1fff1fff9ff08001b002e003b0040003f00360028001a000e0009000b00100015001d00230028002f00340037003900390035002c001f0012000500fafff3fff1fff3fffbff0700110019001f00240024002300230027002f0037003e00440046003f00310020000900f3ffe8ffe4ffe7fff4ff02000f00180016000b00fbffe5ffcfffbdffaeffa5ffa4ffaaffb7ffc9ffdefff7ff0c00190020001f001000f7ffdbffbbff9fff89ff7bff78ff81ff92ffa6ffb9ffcaffd1ffc9ffb7ffa1ff88ff70ff60ff56ff53ff56ff5aff5eff63ff69ff70ff78ff82ff8eff96ff96ff8fff7eff61ff3fff1dfffefee7fedffee3fef4fe0fff2dff47ff61ff73ff78ff71ff61ff4bff34ff1dff0bff01ff01ff0dff23ff3fff60ff85ffa6ffbfffcdffc9ffb2ff8dff5cff29fffffee3fedafeeafe09ff32ff5dff7eff97ffa4ff9cff86ff6bff4aff2aff13ff01fffcfe06ff19ff35ff58ff7aff98ffadffb4ffafff9aff78ff55ff33ff12fffefef8fefbfe0cff29ff45ff5dff6cff71ff6eff63ff55ff4eff4dff51ff5bff6aff77ff7fff7eff79ff76ff74ff74ff7cff88ff94ffa2ffadffb0ffabffa0ff8fff7aff68ff5bff59ff60ff70ff89ffaaffcdffedff08001c0028002d0029001e0012000600fdfffafffeff0d00260042005b0071007b0077006900510034001e000f000c001a0031004d0069007e008c00940094009300960099009f00aa00b500bc00bf00bb00b000a100910083007b007c0086009500a500b100b700b700b300a8009a008f008a008d009500a100b200c200ce00da00e300e800ea00e600de00d600ca00bc00b400b100b200b900c300cf00db00e000df00dd00d600d000d300da00e600fb0010011f012b0130012b0123011501060100010501120125013b014f015b015c0152013f0124010901f600ee00ef00fb000c011e01320143014a014c014b0144013c01310124011a0112010c010e0115011d012a013a0144014a014a0143013701280117010d0106010101070113011e012801300132012f0127011c01160116011a0124012f0135013b013b0135012f012a01260128012b0131013a014301490150015301510150014d01470143013b012f0125011f011b011e0122012c013d014e015c01670166015c014d0136011b010801fb00f600fd000b011f013601430149014a01400132012601160107010001fa00f700fc0002010a0118012901390147014e0151014f014501330120010e01fc00f400f500f900050113011d0125012801200116010e010101f700f100e800df00db00d300cc00c800c400c400c700cd00d600db00d900d600cc00b800a50093007d006f006a006a0070007a00850092009b00a000a1009d009400870077006500530045003c003600360040004f005d00690070006f006600520037001e000a00fdfffbff040016002c003f004d00540051004600360028001c0012000f00120016001a001d001e001c00140009000300fffffafffaff0000060011001d002200230021001b0013000700fbfff3ffefffeffff3fff9ff000009000c000700fbffe6ffcaffaeff96ff86ff82ff89ff9dffb7ffd1ffe6fff2fff0ffe4ffd0ffbaffa7ff97ff91ff97ffa4ffb4ffc6ffd1ffd3ffcdffbdffa9ff97ff84ff75ff6fff71ff77ff82ff8eff98ff9effa0ff9fff9bff97ff94ff93ff93ff96ffa0ffaaffb3ffbfffc8ffc9ffc7ffbeffabff9bff90ff88ff85ff8bff96ffa5ffb5ffc2ffc9ffcaffc4ffb9ffacffa2ff9eff9dffa3ffb3ffc4ffd2ffe2ffebffe8ffe4ffdaffcbffbdffb0ffa5ff9eff9aff98ff9aff9cff9dffa1ffa3ffa0ff9dff99ff94ff8eff88ff85ff84ff84ff89ff92ff9affa1ffa7ffa9ffa7ffa1ff99ff93ff8fff8cff8bff90ff99ffa1ffa5ffa6ffa2ff9cff95ff8aff7eff77ff78ff7dff84ff8fff9cffa9ffb4ffb9ffbcffbaffb4ffadffa3ff99ff94ff94ff98ffa1ffb0ffbeffcbffd7ffdaffd7ffceffbdffa9ff9aff8dff83ff85ff8fff9dffafffc4ffd5ffe1ffe2ffddffd6ffccffc2ffbbffb9ffbdffc5ffceffd6ffdeffe1ffdeffdbffd6ffcfffc9ffc5ffc1ffc1ffc3ffc3ffc4ffc6ffc5ffc2ffc0ffbbffb8ffbaffc0ffc9ffd6ffe5fff5ff04000d000d000400f6ffe3ffceffbaffabffa5ffa9ffb4ffc6ffdaffebfff5fff8fff0ffe0ffccffb5ffa1ff95ff92ff9cffb1ffc9ffe5ff0300190025002a0021000f00faffe3ffcdffc0ffbaffbaffc2ffd0ffe2fff3ffffff05000500fffff5ffe8ffdaffd0ffcaffc8ffceffd8ffe3fff1fffdff020003000100fbfff1ffe6ffdcffd2ffc5ffbdffb9ffb5ffb2ffb1ffafffacffacffaeffafffafffaeffadffabffa6ffa0ff9bff97ff93ff90ff8cff8bff8aff85ff80ff7eff76ff6bff63ff5aff50ff48ff41ff3cff3bff39ff35ff37ff37ff34ff30ff2dff2cff2bff2bff2dff30ff32ff36ff3aff3bff39ff36ff30ff28ff20ff17ff10ff0dff0cff0fff15ff19ff1eff22ff1eff1aff17ff0eff04fffefef9fef5fef5fef8fefbfefbfefcfefdfefbfef5feeefee8fee1fed9fed4fed2fed0fecafec5fec3fec0febbfeb9febbfebbfebbfebefec2fec3fec3fec2fec1febcfeb3feabfea8fea3fea0fea2fea6feaefeb8febdfebffec1febcfeb4feadfea4fe9dfe97fe92fe91fe96fe9bfea2feabfeb4febcfec1febffebefebcfeb6feb0feacfea7fea7feaafeabfeb1febafec3fecefed7fedefee4fee8fee5fedffedafed4fecdfec7fec5fecbfed7fee4fef2fe03ff13ff1eff21ff1dff17ff10ff05fffafef5fef5fefbfe07ff12ff1eff2cff34ff35ff32ff28ff1cff11ff07ff01ff03ff0bff18ff29ff37ff44ff4eff4fff4cff48ff40ff3cff3aff39ff42ff52ff5eff6cff78ff7dff7eff78ff6dff61ff55ff4eff4fff55ff5fff70ff83ff93ffa0ffa9ffabffa9ffa2ff9aff96ff95ff9affa3ffafffc1ffd6ffe6ffeffff5fff7fff2ffebffe2ffdaffd8ffd9ffdaffe0ffecfff6ff01000b00110016001c00210026002d00370042004900500056005500510051004e00470049004d005100590064006f00780079007500710069005c0053004c004b005500640078009300ad00c000d100d900d700cd00be00ad009f00950090009400a200b600ca00dd00ef00fb00fe00fa00f300e700d700cb00c600c800d000e000f4000c012401390147014f0151014b01420139012e0123011f01210125012f013f015001610171017c018401850181017d0176016e016d017001740182019401a401b801c801d101d901da01d101c901c101b801b201af01b001ba01c501d001e001ea01ee01f101ee01e801e501e001db01de01e301e901f60102020b02140218021902180214020f020c020a020b02110216021d0227022b022e02320231022c022b0227022202240228022a023002360238023e02420241024402460242024302440244024702480247024b024d024a024f025202510259025d025b02600263025f025f025c025302530253024e02520255025702600267026b02740275026f026f026c0261025c02580253025302530254025c026002620268026a02680266025f0255024d024202380233022c0227022a02300236023f02440247024b0247023e02330221020d02ff01f301e901ea01ef01f9010c021a0223022a02260217020602f101da01c601b601b001b701c001cf01e401f401fe010302fb01ea01d701be01a30191018601810189019701a701b801c101c101c201b901a50191017c0168015c015501520158015e0164016b016c0166015c014d013b012e0122011601120111011201170118011801190114010c010401fc00f400ed00e600e200df00d900d300cb00be00b400aa009a008c0083007a0073006f006b0066006000580051004b00420037002f00290024001f001a0016000f000300f8ffecffdcffcbffbeffb2ffa8ffa4ffa3ff9eff97ff91ff8bff82ff76ff6bff5fff55ff4eff4fff54ff59ff60ff65ff69ff69ff63ff57ff48ff37ff27ff1aff0dff04ff01ff01ff04ff05ff04ff00fffafef0fee4fed6fecafec0feb8feb4feb3feb3feb7febcfebdfebcfebefebbfeb3feaafe9efe91fe86fe79fe69fe5dfe52fe46fe3afe32fe2cfe28fe24fe23fe23fe20fe1cfe15fe0dfe05fefdfdf2fde7fde1fddffddffde3fde8fdecfdf0fdf0fdecfde6fddafdc9fdbbfdacfd9ffd97fd91fd91fd97fd9dfda3fdacfdb1fdb2fdb3fdadfda7fda1fd9afd95fd95fd91fd91fd97fd9afd9dfda2fda1fda2fda6fda2fd9afd95fd8cfd83fd7dfd72fd6bfd69fd65fd65fd69fd69fd6dfd76fd78fd79fd79fd73fd6cfd67fd5ffd58fd56fd56fd5bfd64fd6bfd74fd7cfd7dfd7bfd79fd70fd63fd5afd51fd4dfd4efd4cfd50fd5bfd60fd60fd63fd60fd57fd4ffd47fd3ffd3cfd3afd3ffd47fd4cfd53fd5afd58fd54fd50fd47fd3dfd34fd2cfd2bfd2efd2ffd34fd3afd3bfd3cfd3bfd32fd2afd26fd1ffd19fd18fd1bfd22fd2bfd34fd3ffd48fd4cfd4ffd4ffd4cfd4cfd4cfd49fd4afd4efd4ffd51fd52fd50fd52fd55fd52fd51fd54fd50fd4ffd53fd51fd4ffd50fd4efd4efd4ffd4efd53fd5cfd63fd6cfd76fd7afd80fd82fd7afd75fd71fd65fd5dfd5afd57fd5cfd62fd67fd71fd78fd77fd78fd75fd68fd5ffd59fd52fd51fd56fd5cfd68fd79fd84fd8dfd93fd92fd8cfd84fd7bfd72fd6dfd6dfd73fd7efd89fd94fd9ffda7fda8fda6fda1fd98fd93fd8efd8bfd92fd9cfdaafdbdfdcbfdd2fdd9fdd8fdd0fdc9fdc0fdb9fdb9fdbafdc0fdd0fdddfdeafdf9fdfffd01fe02fefafdf0fdeafde3fde2fde9fdf1fd01fe14fe1ffe29fe2ffe2cfe27fe20fe16fe10fe0ffe11fe1bfe27fe34fe46fe54fe5bfe60fe64fe62fe5efe5cfe5dfe64fe6dfe79fe88fe95fe9efea5fea8fea3fe9afe92fe8afe87fe8afe8efe97fea5feb0feb8fec2fec7fec4febffebafeb5feb3feb3feb8fec7fed7fee7fef7fe03ff07ff06fffdfeeefee2fed6feccfecafeccfed4fee3fef4fe02ff0fff16ff18ff18ff14ff0fff0bff0aff11ff1dff2cff41ff57ff69ff79ff84ff86ff84ff81ff7aff71ff6cff6eff72ff78ff83ff90ff9cffa5ffadffb2ffb2ffafffadffabffaeffb7ffc1ffcdffdbffebfff7fffeff02000200fffff9fff2ffebffe7ffe8ffeaffeffff6fffbfffdfffdfff8fff0ffe8ffe0ffdaffdaffe1ffedfffdff0c001e002f003900400042003c0033002c00250025002b0034004200530063007000780076006f00640055004a00430043004c005d0073008e00a900bc00c800cc00c900c000b600ac00a500a700b100c100d600eb00ff000f01160114010a01fb00ec00e100d800d800e300f30005011d01340144014d014d0147013f01360131013301390148015f0177019001a401b001b801b601ac01a4019b01920192019a01a601bc01d301e401f501000201020002fa01ee01ec01ef01f401020216022a0243025b02690276027b02770274026e02650266026b026f027e0290029c02aa02b502b802bc02bb02b602b702ba02b902c202d102df02f4020803160329033c03460353035d0362036d037803810391039d03a203ae03bc03c203ca03d403da03e503ee03f403ff0308040a0416042204280437044704530465047704830493049e04a404ac04b004af04b304b404b504bd04c004c304d004d704d504da04dd04db04de04e004e004eb04f8040305190530053f0556056a0574057f0588058905900598059b05a805b805c205d505e605ed05f905010601060406050602060b0615061c063006440655067006830689069806a1069e06a406a606a006a906b406b906c706d306d606e106e606e006e206dd06d106d206d306d106df06eb06f306080717071a07240728072007230724071f07280733073a074d075e076607740779077207710769075a075a075b07580769077d0789079e07ad07b007b707b207a10799078d077b077a077e0781079407a407a907ba07c007b007a407920775076307530743074807510754076707770778077c0776076107500739071c070f070607ff060b0717071e073107380730072e0722070a07ff06f106e006e406ea06ec06fd0608070a0712070e07fc06f306e006c506bb06b106a606ab06ad06ab06b106a906950687067006520641062f061e061f0620061f0629062a06200617060306e305c705a6058405730567055f0567056d056e056d056005460528050205d704b5049904860485048c049704ad04be04c104be04ac04890464043a041104f703e703e003eb03fe030c04170416040404e803bf038a0358032a030403f302f002f70209031b03250328031b03fa02cd029a0267023b0217020302ff0103020c0217021b021302fe01d801a80174013f011001ec00d500ce00d100d900e200e500de00cc00ae0086005c0034001000f4ffe2ffdcffdeffddffddffd9ffccffb5ff96ff6eff45ff1efff8fedbfec7feb6feabfea1fe90fe7dfe66fe44fe1dfef7fdd1fdadfd90fd76fd62fd54fd43fd31fd20fd04fde2fcbefc95fc6bfc4afc2bfc11fc00fcf0fbe3fbd6fbbffba4fb88fb5efb33fb0bfbe1fabffaa9fa94fa87fa86fa7cfa73fa6cfa53fa33fa15faebf9c2f9a5f986f971f96af95ff95bf95df950f940f92ef907f9dbf8b5f883f855f834f811f8f8f7eef7ddf7d0f7c8f7aff795f77df752f729f70df7e7f6c7f6b7f69ef68cf687f678f668f65cf63df61ff609f6e1f5baf5a0f578f557f545f524f509f5fdf4dff4c4f4bbf4a2f48ff48bf476f467f466f451f43df437f41ef407f4fff3e5f3d1f3d0f3bef3b2f3b3f39ff38cf383f35ff33bf321f3f2f2cdf2baf29af28cf293f28af28df29ef292f287f285f264f246f234f20bf2f0f1edf1dbf1d8f1ecf1eaf1ecf1f6f1dff1c5f1b2f17ff151f135f10bf1f4f0f9f0f0f0f9f017f11cf124f135f125f112f106f1ddf0c1f0bdf0a8f0a5f0bcf0c2f0d5f0f4f0f2f0eff0eef0caf0a8f094f066f047f041f02df02ff049f050f061f07af074f06ff06ff04df034f02bf00ef005f015f013f021f03ff042f04bf05df04bf038f02ff00ef0f7eff6efe4efe4effbef01f013f033f033f036f042f033f02af030f023f025f03bf041f057f07cf085f095f0aef0a6f0a2f0abf09af096f0a6f0a5f0b4f0d8f0e6f0fbf01bf11ef123f131f122f11cf126f11ef128f148f154f16df195f1a4f1b8f1d0f1caf1caf1d1f1c3f1c5f1dbf1e1f1f7f11ff236f256f27df288f293f2a4f29ef29ff2acf2a9f2b3f2d0f2e3f203f32ff347f365f389f394f3a0f3b3f3b2f3baf3d1f3dbf3f6f322f43ef464f495f4b0f4cff4f4f4fef40df525f529f535f550f55ef579f5a3f5bef5e3f510f628f643f664f672f685f69df6a9f6c1f6e3f6f9f61cf74af76cf797f7c6f7e4f707f82bf83df855f872f882f89cf8bdf8d6f8fcf826f942f968f994f9b4f9d7f9fcf916fa38fa5dfa78fa9afac1fae2fa0cfb38fb5cfb85fbaffbd2fbfbfb24fc45fc6bfc91fcaefccffcf0fc0afd29fd48fd67fd8efdb5fdd8fd04fe32fe5afe85feaefed2fef6fe13ff2dff4dff6aff88ffb0ffdaff06003a0067009200c200e700060125013d01550171018b01ac01d801030236026e02a202d7020a033003540374038a03a503c103da0300042d0456048d04c904fb04310563058705ad05cc05db05f4050f06240649067806a506e206210755078f07c007dd07fd0715081a082b0840084e0871089f08cb080a0948097709af09d909e909020a120a100a220a3d0a560a890ac10af10a350b750b9d0bcb0be60be80bf50bfa0bf30b0c0c2a0c440c7f0cbc0cec0c2d0d5d0d720d920da30d9c0dab0db70dbd0de60d130e3a0e800ec00eea0e1e0f410f480f580f590f4b0f5a0f690f720f9e0fce0ff30f2f105f107a10a310b610ae10bb10c010b610cd10e510f7102d1160118311be11e811f31110121b120a1212121212031218122e123c126c129612ac12db12fa12fb120c130b13f412fb12fa12ee120c1328133c1373139e13b113d813ea13df13e613d813b713b513ae13a113bf13db13eb131b143c1440145714551438142f141714f413f913fc13f9131f14411452147b148f1485148c147a144b143b14241402140a141414141437144e144e1464146214421437141b14ee13e513d713c013d213de13dd13fa130414f413f913e813c013b4139a137513781371135f1370137313611369135e133c1334131b13f212e812d412b412b612ab12931299128f126e12671252122c1222120d12ec11e911d911bb11ba11a81184117b1165113d1132111c11f810f010dd10ba10b3109f1079106c1052102a101d100310e00fdd0fcc0fad0faa0f970f720f650f470f1d0f0d0fef0eca0ec30eb00e930e920e830e620e540e330e010ee40dba0d850d6d0d500d320d310d290d170d180d060de10cc70c9a0c600c380c080cd80bc80bb70ba60bb00baf0ba10b9b0b7c0b480b1a0bd50a870a540a230af609ec09e809e609f809f809e409d309a80964092609dd08920862083c0823082b0835083b084b0843082208f807b4075d071007c0067b0656063b0630063e064b06500653063c060d06d40587053105e804a40472045d045504580467046f04680456042b04ee03a90356030303c1028902620255025302570261026202520236020502c3017b012f01e800b000850069006100630069006d00660050002d00f6ffb0ff63ff16ffd4fe9efe76fe65fe64fe68fe70fe74fe68fe4cfe1cfedafd90fd40fdf0fcb0fc80fc63fc5dfc62fc6dfc7afc77fc63fc3efc01fcb4fb65fb14fbcffaa0fa7efa73fa7efa87fa91fa99fa88fa62fa2efae2f98ff943f9f9f8c2f8a5f894f896f8a7f8adf8adf8a8f883f84ff818f8cff788f751f71df7fcf6f4f6ecf6eef6faf6f0f6dcf6c4f691f654f61ef6daf59df579f553f53af536f527f51bf516f5f9f4d9f4bff48bf459f437f405f4def3cdf3aff39af394f377f35df34cf31ef3f1f2d3f29ef273f25af22ff20ff204f2e1f1c4f1b6f18ff16bf156f128f1fff0eaf0c1f0a6f0a1f086f073f071f053f036f021f0eeefc1efa4ef6def41ef2fef0beff5eef7eee1eed4eed6eeb5ee95ee80ee49ee17eefaedc6eda7eda8ed95ed91eda8eda0ed9ceda2ed7eed5aed40ed02edcfecb6ec88ec72ec7eec74ec7bec9aec92ec8aec8dec63ec3aec22eceaebc3ebbbeb9feb9cebb6ebb3ebbcebd6ebc9ebbbebb7eb8ceb69eb5aeb31eb1eeb27eb19eb1deb39eb34eb37eb47eb2feb1eeb1feb00ebf2eafdeaeaeae9ea00ebf4eaf0ea00ebebeaddeae3eac7eabceacdeac4eaceeaf2eaf5ea02eb1eeb0feb05eb0aebe9ead6eae0ead4eae1ea0aeb17eb38eb69eb6feb77eb86eb64eb47eb3beb10ebfdea0feb12eb33eb75eb9debd2eb0eec19ec22ec2eec0aeceeebe7ebc9ebc6ebe9ebffeb30ec7beca4ecd2ec02ed00edf7ecefecbeec9aec94ec7eec87ecb7ecd9ec12ed64ed93edc0edf0edf3edf1edf5edd7edcbedd8edd3edeaed20ee41ee73eeb2eecbeee4eeffeef3eeefeef5eedeeedbeef1eef5ee10ef41ef5aef84efbdefd6eff8ef25f033f04bf070f07bf093f0b8f0c2f0d6f0f6f0fdf011f131f13af154f182f19bf1bef1eaf1fdf118f237f23cf249f261f265f27cf2a8f2caf201f34af380f3bff302f424f442f45df457f457f462f461f474f49df4bff4f7f43df570f5aaf5e3f5fcf513f62af62bf637f64ff661f68cf6caf602f74af798f7cff704f834f849f85cf86ff876f88af8a6f8c2f8f1f829f958f990f9c7f9edf913fa33fa47fa62fa81faa0fad3fa0dfb43fb86fbc4fbf2fb1ffc42fc53fc64fc74fc85fca6fcd1fc02fd44fd8dfdcffd10fe41fe5efe6ffe71fe69fe69fe75fe91fec8fe14ff6fffd7ff37008900c700e300e300d200ae00880077007d00a600f4005c01d8015702c0020f033b0338031503e102a4027c0277029602e8026503f4038f041c057e05b705b90583053605dc04850459045f0494040805a4054706ea066c07b707d307b40761070707af0668065f068f06ed0685073308d7086f09d109ed09d9098f091a09ae0855081c0829087008e0088409310ac40a410b8b0b8f0b6c0b210bbb0a6b0a370a250a5a0abe0a3b0bda0b700cdb0c2d0d470d230de90c920c2c0cef0bd10bd20b180c810cf50c840dff0d4e0e8a0e950e6c0e420e080ec90db90dc30de00d340e960eef0e570fa10fc20fd90fc80f920f6d0f460f200f2a0f480f6f0fc00f11104d109510c010c610d110c710a810a410a1109b10bf10e81006113f116a117811921196117e117a116f115b116d1181118e11bf11e411f2111712281219121d121412f91100120412ff11231240124c12731289127f12831274124d1240122c121212221234123f1270129712a912d012df12cf12cd12b512871278126112431250125c1260128912a512a912c012bf129f129512771247123a122b1218122f12471258128d12b312bf12de12e312c312b41292125a12421224120012081210120f1231124512421257125412321225120812d811cc11be11ac11c611e011f11120123f1246125c1254122d121612ea11aa118b1167113e113e1140113f115e1170116c117c11751150113f111d11ec10de10cd10b910cd10e410f2101a1136113a11461134110211dc10a11055102910fd0fd00fcf0fd30fd40ff40f0710061011100110d60fbb0f8b0f4c0f2f0f150fff0e130f290f390f630f790f730f730f520f0e0fd40e880e320efd0dcc0da40dab0db70dc10de70dfe0dfa0df70dd60d970d600d1b0dcf0ca50c860c710c870ca20cb80cdd0cee0cde0cc60c8d0c330cdd0b7e0b1f0be50abd0aa70abc0ada0af50a1a0b230b0c0be90aa40a460af1099809480921090f0912093a0960097c099909930964092409c6085708f6079b0754073b073707470772079607a907b30799075e071407b3064c06fa05b6058b0585059005a905d005e605e605d605a70560051105b90463042404f603dd03df03eb03fc030e041104ff03e003aa0363031b03d202910261023e02290221021e021b0217020502e901c30192015b012501f100c2009b007e006b005c004c003d0028000a00e8ffbdff8cff5aff23ffedfebffe91fe65fe45fe25fe07fef0fdd3fdb3fd96fd72fd4afd27fdfefcd5fcb4fc90fc6bfc4cfc2afc07fce9fbc1fb98fb72fb42fb11fbe6fab3fa83fa5cfa30fa08fae7f9bef995f976f94df924f903f9dbf8b7f89df87bf85cf846f825f804f8ecf7c6f79af773f73ff70cf7e3f6aef67ff65ef635f614f602f6e2f5c3f5aff58cf567f54bf51cf5f0f4d1f4a4f47ef46cf450f43cf43af428f418f412f4f1f3ccf3aef374f33bf311f3d7f2a7f290f271f263f26cf265f265f270f25bf241f22cf2f4f1bbf195f15df134f129f118f118f131f136f140f151f13cf11df101f1c2f080f051f016f0f0efecefe4eff2ef1cf030f047f062f054f03df027f0edefb5ef8fef58ef39ef3def38ef4aef75ef85ef9aefb4efa1ef88ef73ef38ef06efebeebeeeaaeebaeebeeedaee0def23ef3fef5fef51ef40ef31effbeecceeb3ee88ee75ee80ee7dee92eebbeec7eedaeef4eee4eed4eecdeea3ee85ee7cee61ee5eee76ee7cee95eec1eecfeee1eef8eee8eeddeedceebbeea6eea4ee8dee87ee98ee93ee9ceeb5eeb3eebaeed0eec8eecbeedeeed6eedceef5eef6ee00ef18ef15ef1aef2def27ef2def44ef46ef56ef76ef7fef91efabefa8efabefb6efa4ef9befa1ef95ef9defbcefcfeff5ef2bf04bf073f0a0f0a8f0b1f0bdf0acf0a3f0abf0a1f0adf0d2f0ebf015f152f176f19ff1cbf1d1f1d4f1d9f1bff1b0f1b4f1a7f1b2f1dcf1fdf132f27af2acf2e1f218f32af338f344f32ef31ef31ff311f31af341f362f398f3e2f317f44ef484f495f49ef4a4f489f473f46cf45af462f487f4aaf4e4f431f56cf5abf5e6f5fcf509f610f6f9f5eaf5e6f5daf5e5f50cf632f66df6b6f6f0f62bf761f775f782f786f771f762f75cf751f75df77ff7a3f7dbf71ef854f88ff8c4f8dcf8f2f801f9f8f8f5f8f8f8f5f807f92bf94bf97ff9bdf9edf923fa53fa6afa7dfa8afa84fa83fa88fa85fa94fab1facefafbfa30fb5bfb8bfbb6fbd1fbebfbfefb04fc11fc22fc31fc4cfc6ffc90fcb9fce4fc08fd2cfd4afd5efd74fd86fd95fda8fdbffdd7fdf7fd17fe35fe56fe72fe89fea2feb8feccfee7fe05ff28ff50ff78ffa0ffcaffecff07001f002f003a004700550068008600aa00d6000801370165019001ab01bd01c901cd01d101d801e201f9011e0248027c02b802ee022003490362037103760370036d036f0373038703ab03d6030c0447047e04b104d904ef04fd04fc04f004e704e104de04ee040c0533056905a205d7050b06300642064d064a063b06310626062206330650067406a906e20613074407660774077c0775075f07530749073f074d0765078007af07e1070708310850085b08660865085608520850084c085d0878089208bc08e70806092c09480951095c0960095409530952094b095809690976099609b709cc09ec09060a100a230a300a2f0a3b0a460a490a5c0a6f0a7a0a960aaf0abc0ad50ae90aef0a010b0e0b0f0b1e0b2c0b2f0b410b4f0b500b610b6d0b6e0b7f0b8e0b940bb00bca0bda0bfc0b190c250c3f0c4c0c470c4f0c4d0c3d0c440c4c0c4e0c6b0c890c9d0cc60ce60cef0c030d070df40cf10ce70cd00cd90ce70cf00c190d450d650d980dbb0dc30dd40dd30db70dac0d9b0d810d870d920d9a0dc20dea0d030e2d0e4a0e4e0e5c0e590e410e3d0e330e200e2b0e390e400e640e850e960ebb0ed20ed20ee00ee10ecf0ed00ec60eb10eb80ebb0eb40ec90edb0ee00efd0e110f150f2d0f370f2e0f3a0f390f270f2c0f270f160f1f0f220f1c0f310f3d0f3d0f550f600f570f630f5f0f480f460f3a0f1f0f200f1a0f0d0f200f2d0f2f0f4d0f620f640f780f7b0f690f670f550f320f270f150ffa0eff0e010ffc0e170f2b0f300f480f500f410f400f2c0f050ff30edb0ebb0ebc0ebe0ebf0edf0efa0e070f260f320f250f200f050fd50eb70e910e680e600e5b0e590e780e930ea40ec50ed20ec70ec20ea60e780e5b0e350e0c0e040eff0dfc0d190e300e3b0e560e5b0e490e3c0e190ee40dc10d950d660d570d4c0d410d550d650d6a0d7e0d820d710d680d4c0d1d0d000dda0cac0c9b0c890c730c780c790c6f0c750c6f0c580c4e0c340c0b0cf20bd10ba50b900b790b5c0b540b480b350b350b2d0b180b110bff0ae00ace0aaf0a820a640a3f0a110af609d609b409a70997098309810976096109570940091c09ff08d508a4088108590831081e080808f307ef07e107ce07c207a4077a0757072407eb06bd0689065a063e0621060a060506fb05ee05ea05d705b9059e0573053f051105d804a10478044c04290416040104ef03e703d403bb03a103760341030b03ca028c0257022402fe01eb01dd01db01e001de01d801c801a30171013101e100930049000200ceffabff95ff90ff91ff8eff8cff7aff53ff22ffdffe8efe41fef5fdb1fd86fd68fd59fd60fd67fd6bfd70fd5efd37fd06fdbcfc65fc12fcbafb6cfb38fb0dfbf5faf6faf5faf6fafcfaecfacbfaa2fa5ffa10fac7f975f92bf9fbf8d1f8b9f8baf8b7f8b9f8c0f8aef88df866f820f8cff782f728f7daf6a5f673f656f654f64ef651f65cf64cf634f618f6ddf59bf55ef511f5d0f4a7f479f460f45ef450f449f44cf431f411f4f1f3b3f376f343f3fef2c8f2aaf280f268f267f253f248f247f22af20ff2fbf1ccf1a1f183f150f129f114f1eaf0c9f0bbf095f076f067f03ff01ff010f0e9efccefc2ef9eef81ef75ef4def29ef15efe7eec2eeb2ee8cee74ee73ee5dee51ee58ee41ee2cee23eef7edcdedb2ed7bed50ed3eed19ed09ed15ed0ded10ed27ed1eed16ed17edf1ecccecb7ec83ec5eec53ec34ec2cec41ec3eec48ec65ec5cec55ec57ec2fec0becf7ebc2eb9deb96eb79eb72eb8aeb86eb93ebb3ebacebaaebb4eb91eb74eb68eb38eb15eb0eebeeeae3eaf4eae7eaeaea07ebfeeaffea12ebfceaedeaf1eaceeab7eab7ea95ea87ea94ea84ea88eaa8eaa8eab6ead8ead4ead7eae6eacbeab8eab6ea8fea7aea80ea6eea74ea9aeaa7eac7eafbea0beb20eb3deb2deb20eb1febfaeae6eaedeadfeaecea1beb33eb60eb9febb7ebd4ebf5ebe7ebdbebdaebb5eba3ebaceba2ebb8ebedeb0cec41ec88eca8ecccecf3ececece8ecedeccfecc2eccfecc9ecdfec12ed2fed60eda0edbceddcedffedf8edf4edf9ede0edd9edeaedeaed06ee3dee61ee96eed9eefcee21ef48ef49ef4def59ef49ef48ef5eef65ef83efb9efddef11f052f076f09df0c9f0d6f0eaf008f110f127f153f172f1a3f1e4f113f24df28ef2b4f2e0f210f327f347f371f38bf3b3f3e7f30ef442f47ef4a8f4daf411f533f55ef58ff5b2f5dff516f640f674f6aff6dbf60bf73ef75ef784f7aff7caf7eff71cf841f870f8a5f8cef8fdf82df94bf96df98ff9a3f9bdf9dff9fbf924fa58fa86fabffafcfa2dfb5ffb8dfbaafbc7fbe2fbf4fb0dfc2bfc4afc76fcaafcddfc17fd50fd7ffdadfdd5fdf0fd0bfe25fe3dfe5ffe89feb6fef1fe31ff71ffb4fff0ff2300510073008e00a900c100dd0003012f016401a001dd011a0254028302ac02d002e80200031d03390360039003c203fc0339046c049d04c704e104f8040c0519052d05490567059405c705f4052806560674069006a306a706b006bd06c606e206080730076807a107cf070008280839084c085808570866087b088e08ba08ef0820096209a109ce09010a2a0a3c0a580a700a7d0aa10acb0af00a2f0b720bab0bf60b390c670ca10cd00cea0c130d380d4f0d7e0dad0dd10d0f0e4c0e790ebb0ef70e1e0f580f8a0fa40fd20ff80f0b103210521060108610a710b510dc10fd100c1132114f115711741187118211921199118a11941199118d119e11ab11a811c011d111cd11e011e711d411d811cf11b211b011a81190119911a2119b11b511c811c511dc11e811da11e211dd11c311c911ca11bc11d511ed11f711241249125912811298129312a612a81293129f12a6129f12c212e412f7122e135a136d139a13b213ab13bd13be13a813b613bf13bc13e2130414151448146a146e148b1490147414731461143b143a14341423143c144d144d146c1479146a147214621438142b141214e813e713e213d213eb13fa13f5130c140f14f613f813e513bb13b413a5138c13a013b013b413de13fd13041424142d141b1424141e14061417142914331469149d14c2140615361548156e157815651570156d155e157e15a115bd15051645166f16b016d416d016db16c9169b168b167516561668167e168a16bc16df16e316f416e216a71678163016d1159515571516150415f414da14df14cf14a0147d143914d31380131a13a61257120812ba119711711140112c110511c51096104e10f00fac0f5b0f010fcd0e980e610e500e390e180e150e020edf0dd20db40d850d6f0d4c0d200d130dfe0ce30ce90ce90ce10cf60c010d010d160d1b0d120d1b0d130dfd0cfb0cef0cdb0ce20ce30ce00cf70c050d0a0d220d270d1b0d1b0d080de30cca0ca40c780c610c420c220c1a0c050cea0be00bc70b9f0b820b500b110be10aa30a600a310af809bf099e09730944092709fe08ce08a908750838080708ca07880757071c07e206be0695066c065806410629061d060706ee05de05c205a0058a056b054c053c052b0520052505280530053f0548054d0553054b053d0530051705fe04eb04d604c704c004ba04bc04c004bb04b604ad049804790450041b04e403aa036b033203fb02c5029702670233020202c7017c012f01d5006c00040094ff1fffb4fe4cfee7fd91fd3dfde8fc9ffc4efcf5fb9efb3cfbcefa64faf3f982f91cf9b6f858f80ff8c8f789f75bf729f7f4f6c8f691f654f61df6d9f597f565f52ef502f5eef4dbf4d6f4e6f4f0f4fbf411f517f518f51cf50cf5fcf4f7f4e6f4e1f4f1f4fbf413f53ff55ff583f5aff5c2f5cef5dbf5cef5bef5b5f59af589f58af57df57cf58cf588f588f591f57df564f551f520f5ecf4c4f485f44bf423f4e8f3b2f38ff357f323f300f3c7f28ef262f21ff2def1abf160f116f1dbf089f03df006f0bdef7def58ef24effceeebeec6eea7ee97ee6cee41ee23eeededbceda3ed7ced69ed73ed71ed82edabedbdedd3edf3edefedeaedeeedd1edbeedc1edb1edbbede4edfced29ee6bee8deeb3eee1eee1eedeeee4eec2eea8eea6ee88ee80ee98ee94eea0eec2eebaeeb2eeb2ee7fee46ee18eebded68ed2cedd2ec8dec69ec27ecf7ebe1eba4eb6beb40ebe4ea86ea38eac0e953e901e994e83de80be8bde785e76ae72ce7f9e6d8e689e641e60de6b5e56ce541e5fee4d6e4d2e4b7e4b6e4d4e4d3e4e2e407e507e515e537e538e54be578e589e5b1e5f4e51ae656e6a9e6dbe61fe779e7ade7f2e74de881e8c6e81de94ce989e9d9e901ea38ea83eaaaeae5ea37eb66eba6ebf7eb1dec50ec8eec97eca2ecb8eca0ec94ec9bec7fec79ec90ec87ec90ecafeca7eca3eca7ec7aec4dec27ecd7eb94eb69eb23ebf6eae9eac7eabaeac6eab2eaa4ea9cea69ea39ea12eacbe993e973e942e92ee93de93fe95ae98ee9a7e9cce9fae901ea0bea20ea18ea20ea3fea4dea79eac6ea04eb5bebc8eb1aec77ecdbec18ed5beda7edcfed06ee53ee8aeed9ee44ef98ef03f07ef0d8f03af19ff1d9f117f25bf279f2a0f2d7f2f2f220f35ef382f3b5f3f2f310f435f45ff467f477f48af482f488f495f487f489f495f48af489f490f47ff478f479f468f463f463f451f44df44ef43bf433f430f41df416f41af418f426f444f461f48ef4c8f4fbf436f573f5a0f5d0f502f629f659f692f6ccf61bf778f7d7f748f8bff82bf99af903fa57faa9faf8fa37fb80fbd5fb2bfc94fc09fd7efd01fe85fef8fe66ffc5ff0a004a008100a600d100030133017001b401f40139027702a102c202d202cd02c102aa028c02770265025502540257025a025f025a024a0231020a02d901a5016b0132010101d500b000940079006500510036001d000100dfffc3ffa8ff8dff80ff79ff73ff7aff87ff94ffaaffc0ffd3ffefff0f002b0054008400b200ed002b016201a401e90128027302c00208035e03bb0312047704e2044005a30507065a06b10606074f07a307f80742089c08ff085509b309130a5f0aae0af70a290b600b960bbc0beb0b1b0c410c790cb20cdd0c130d430d5e0d820d9d0da10db10dbb0db50dc30dcf0dcd0de40dfa0d010e1d0e330e380e530e640e640e7e0e900e950eba0ed90eea0e1e0f4d0f690fa30fd40ff10f2a1058107110a810d710f610391174119d11ec1134126a12be12051335138013bf13ea1332146e149814e314211549158f15c615e1150f16281625163516341622162a16241612161e161b1604160116e815b21587154415eb14a5144e14f013af1365131613e2129d124a1201129b111f11ac101d10850f040f770eef0d8b0d200db70c6b0c100cab0b560be30a640afc097e090109a8084b08f707ce079f076f075f073d070d07f306c506880669064206180618061906190642066a068806c206f306150750078207a707e90729085e08b5080c095209b1090c0a530ab20a0e0b570bb60b150c660ccf0c380d8c0df40d550e9a0eee0e3e0f760fbf0f0a1048109c10ef1035118f11df111212541286129712b612cd12cf12ee121113291362139a13c413081439144a146e147a1465146a1467145314681480148f14cc14051528156a1596159f15bf15c515a915b015ae159d15be15e015f91545168a16bb160d1745175a178a179d179217a717ad17a317c517de17eb171e1841184e1875187f186a18681848180f18ed17ba177b1758172c17f916e016b81683165e161e16ca157c1513159b142d14a2130d138b12f9116611e4105210c10f3e0fa40e060e730dc50c0f0c640ba40ae50933097208b90715076506c0052d058b04f1036703cb023102a40105016800dbff44ffb7fe3cfebafd46fdedfc91fc3ffc04fcc6fb8ffb69fb3bfb0dfbeefacbfaabfa9bfa8ffa8bfaa0fac0faeafa29fb71fbb8fb06fc4ffc8bfccafc06fd35fd6bfdacfdeffd4bfec0fe39ffc5ff6300f2007e010a027c02df023c038503d00328047d04e5046605e805730606078607fd076708af08ed08240947097209a809e109310a8f0aec0a560bba0b040c4c0c810c970cab0cb40cb00cc10cd60ceb0c1c0d520d810dc30dfb0d1d0e470e5d0e5c0e6b0e700e650e720e7e0e840ea30ec00ed20ef80e130f1f0f390f470f440f4f0f4c0f3c0f370f240f080ffd0ee70ecb0ec00ead0e960e8f0e7d0e640e4e0e250ef20dbb0d6f0d1f0dce0c6c0c140cc40b670b150bc90a6c0a110aad092d09ac081c086e07c6061c066105b90417046e03df025302b80129019200e0ff30ff71fe9afdccfcf6fb18fb50fa86f9bdf80ff860f7abf60cf662f5aaf4fff346f381f2cdf115f15ef0bfef22ef90ee1aeea8ed3aeddfec81ec25ecd6eb7ceb29ebe5ea99ea5aea31ea09eaf3e9f1e9eee9fae917ea2dea4fea7bea9fead3ea11eb46eb91ebeeeb45ecb0ec29ed98ed19eea4ee1defa6ef36f0b7f047f1daf15bf2eef288f30ff4a3f43af5bbf546f6d3f64af7cef755f8c8f848f9cbf93cfab9fa35fb99fb05fc6afcb1fcfefc48fd7afdb3fdeefd1dfe57fe93febffef3fe23ff3fff5bff71ff72ff73ff72ff69ff6aff72ff77ff86ff98ffa3ffb1ffbaffafff9cff85ff63ff43ff27ff0cff00ff03ff08ff1aff32ff3dff41ff41ff2eff0effedfec0fe92fe72fe57fe48fe4efe50fe53fe5cfe53fe39fe1afedffd98fd57fd04fdb6fc80fc3ffc05fce7fbb6fb78fb47fbf9fa96fa38fabbf934f9c2f839f8b1f749f7d0f654f6f2f572f5e4f467f4c2f310f373f2b5f1f1f04cf08fefd5ee3fee8fede1ec51ec9eebe6ea4cea95e9dde847e898e7f0e669e6cce538e5c2e431e4a8e33ae3b0e22fe2cbe152e1ebe0a6e052e014e0f5dfc4dfa8dfa7df8edf87df9adf97dfa9dfd6dff4df2ce081e0c9e02fe1ace112e294e22be3a3e32ce4c6e448e5dee584e613e7c1e783e82ee9f5e9ccea82eb48ec15edb9ed6aee1fefaaef48f0f5f07ff121f2d6f269f30ff4bcf439f5bff541f68af6d5f623f743f770f7abf7c2f7eef72bf843f865f88ef888f87df871f836f8fbf7cbf77ff73ff716f7dff6b5f69af66cf643f61af6d2f588f53ef5e0f489f443f4fbf3caf3b0f394f387f38af381f378f372f35cf345f336f321f319f326f339f361f39cf3d4f319f463f498f4d2f40ff534f560f598f5c3f500f654f69bf6f0f655f7a2f7eff73ef866f88cf8b4f8b4f8b9f8cef8c5f8c8f8e4f8e4f8eaf801f9f1f8daf8c6f882f836f8f2f785f716f7bbf645f6d7f580f511f5a8f44ff4d3f355f3e1f246f2a4f10ff15df0abef10ef68eecded4bedbfec44ecddeb65ebf4ea8eea14eaa1e93ae9c4e85ee80fe8bfe788e76de755e758e772e788e7afe7e3e70ce841e87fe8b5e8fee853e9a8e91deaa4ea2bebd2eb8aec38edfaedbeee71ef37f0f9f0a7f16bf232f3e5f3b3f48ff559f636f715f8ddf8b3f981fa2cfbdffb8bfc14fda7fd37fea9fe2affacff10007b00e20024016701a101b401c601d401c001ad019a016c0142011a01db009d0060000e00b8ff61fffcfe94fe29feb3fd3efdcbfc53fce0fb6efbfdfa96fa36fad9f981f930f9e9f8a8f869f837f80bf8e2f7caf7bbf7b4f7c6f7e9f714f854f8a3f8f5f857f9c2f92afa9ffa18fb8dfb13fca6fc36fdd8fd8dfe41ff0300d00096015e022903e5039b045405ff05a1064907ea0786082709c109500ade0a620bda0b480ca50cf30c3a0d6e0d920dad0db50dac0d9c0d830d5b0d280def0cb10c6a0c1d0ccc0b6d0b040b990a1b0a92090c097908dd074f07c0063306bc054505d0047004070498033b03d1025d0201029f013e010701da00b400ba00c700d5000701350157019401ce01f9013f028d02da024c03ca034804eb0497053606e80699073808e2088a09230aca0a740b160cc70c7c0d250ed40e7e0f1510a8102b119b1108126412b012ff1246137d13b513e413051420142b1424141614f413c2138e134a13f712a8124e12e911891119119e102a10a70f1b0f9d0e100e780df30c640cce0b500bc80a350abe094009ba085508e90773072607da0686065d0635060306ff05fd05ee050d062b0637067306b106db0634079307e1075e08dc084509df097e0a030bb20b640cfc0cba0d790e1f0fe80fb31067113c121013cb13a21473152716f216b2175118ff18a019211aaf1a321b9c1b141c7c1cce1c351d8e1dcb1d141e491e611e811e891e721e641e401e031ed51d941d421d071db91c571c101cb41b411be41a6f1adf196719d9183518b31720177c1602167f15ef148e142014a5135513f2127b123112d41165112511db1087106c104b10221031103810301056106c106d109110a1109f10c410de10f21038117d11bc1127128c12e1125113ac13e9132b145414671488149a14a214c714e7140115311558156b1582157c1554152615dd147a141b14b1134213e8128a122912d611761105119110fb0f4a0f980ec80de80c1b0c490b7b0ad2092c098c080f088a07ff068806f8055705cc042b048103fc027502f201a4015d011d010d01fe00ee0002010a0107012301340137015d0180019f01e80137028602000384030404a7044b05e1058f063707c5076308f9087709080a9a0a1e0bbb0b610cfb0caa0d5d0efa0e9c0f3110a61017117411af11eb1124124e128712ca120c136013b81303144b147d14921493146c142514d51372130713ab124f120112cd11951161113711f110911023108e0fe20e2e0e600d990ceb0b3f0bab0a3d0acd09690913099f081a088e07d7060b06420567049603ea024902c70171012501eb00bc0076002200c6ff43ffb2fe24fe8cfd03fd9bfc4afc1bfc10fc15fc2afc43fc4dfc4afc2cfcf3fbb2fb60fb04fbbafa7bfa4cfa3ffa40fa4dfa6dfa7ffa86fa8bfa6efa3bfa04fab1f956f90cf9b3f863f82df8edf7b4f78ef74df705f7c2f65df6e8f575f5e4f451f4cdf335f3a5f22ef2acf139f1def074f010f0beef57efefee90ee19eea0ed2ceda6ec28ecc0eb56eb02ebccea99ea80ea84ea86ea95eaafeabceaceeae3eae6eaf3ea0feb25eb54eb9febf3eb64eceeec76ed0deeaaee2eefb3ef33f096f0fbf065f1c2f135f2bbf240f3e4f399f43df5f1f5a3f62ef7b7f731f87cf8c9f816f945f985f9d8f91dfa7dfaf0fa49fba8fb05fc33fc52fc64fc44fc1afcedfba2fb62fb3dfb0dfbf4faf7faedfaecfaf5fadafab0fa80fa24fab9f953f9d2f850f8e8f77bf71ff7dff697f653f61cf6c8f56af510f594f40cf48df3fcf273f20af29af13af102f1c2f084f05cf021f0deefa4ef4defebee94ee29eec5ed78ed22eddcecb5ec81ec5dec54ec37ec1fec1becfbebddebd1ebaaeb88eb78eb4feb36eb39eb28eb29eb49eb54eb72ebabebc4ebe4eb14ec1bec23ec38ec25ec18ec1dec06ec05ec22ec2cec4eec87eca2ecccecffec02ed0aed16edf5ecddecd6ecb1eca4ecb3ecacecbdece3eceaecf8ec0bedf5ecddecc2ec86ec59ec3dec13ec05ec13ec1dec46ec82ecaaecdeec13ed2aed45ed5eed60ed71ed8eeda3edd5ed1cee63eec6ee37ef9bef0ef084f0e7f056f1c5f124f293f20cf37bf302f497f423f5c5f56ef603f7a4f746f8cbf855f9ddf948fab8fa28fb84fbedfb5afcb3fc1afd86fddafd38fe95fed4fe13ff49ff5eff73ff86ff7dff75ff70ff5eff56ff54ff41ff35ff2cff0dffe8fec0fe80fe36fee7fd89fd2cfdd6fc7bfc2dfcf0fbb3fb7bfb52fb29fbfdfad4faa8fa7afa4ffa20faf4f9d2f9b4f99bf98ff986f980f981f980f980f985f988f98af992f999f9a6f9b9f9ccf9e9f90efa33fa5ffa90fabffaf3fa27fb53fb83fbb0fbcffbeffb0dfc1afc29fc3bfc42fc4dfc5dfc67fc79fc8efc98fca6fcb6fcb6fcb3fcaffca0fc8efc82fc71fc64fc5efc5afc5dfc63fc64fc66fc65fc59fc49fc38fc1ffc07fcf5fbe5fbddfbddfbe2fbeefbfafb07fc19fc28fc33fc44fc53fc63fc7efc9cfcc0fcf3fc27fd5efd9ffddbfd17fe59fe95fecdfe0bff44ff80ffc2fffdff40008f00d70025018101d90133029902fa025f03c80329048b04ef0444059905ef053a068606d80623077407ca071a086e08c208070946098109b009da09fe09190a390a5a0a760a960ab60ace0ae40af20aed0adc0ac10a990a680a2e0aee09b20974093409fa08ba0872082c08d8077c072507c0065506fa059b053c05f004a0044c040b04c50377033603ec02980259021902d601ae01890164015a01510144014c01530155016b0181019701c601f9012d027d02d10223038603e40337049704ef0437058905da0520066d06bc06050752079907d507150851087f08ad08d808f80818093109410950095a0955094d093c091b09fa08d4089f086b083608f607b90779072e07e40694063b06e40589052a05da048b043a040104cf039c037c035b03370326031003ef02e202d502bf02c002c602ca02e60204031f0353038b03b803f8033a047004b904060549059d05f6054506a10601075807bb071e087508d3082e097b09cc09170a510a8d0ac30ae90a110b360b500b6f0b8a0b9d0bb20bbd0bbc0bbc0bb30b9a0b800b5c0b2f0b080bdf0ab20a8c0a620a300a030ace098c094809fa08a1084b08ed078f074007f206a90672063906fe05ce0592054e051205cc047c043904f803bc03950370034f0341032e0314030603eb02c102a2027b024b022e02170204020b021b022e0258028302a402ce02f102070325033a0343035a0372038403a803d60302043b047404a804e704230552058505b505d705fc052106450670069b06c406f506260753078307ac07cc07e907f807f807f407e707cf07b907a2078a07780768075607470733071807fc06d1069b0669063006f305c505960567054f053d05280521051605ff04f204db04b50499047a0454044304380430043f04530468049104ba04dc040c0539055d058f05be05e705230662069e06e5062b076d07b407f10723085b088608a108be08d508e308f308fe08060914091f0924092509200915090109df08b60883083f08f507a7074f07f4069d064006eb059b054205e80496043904d2036903f3027a0207028e011901b5005500fdffbdff81ff48ff21fffbfed1feaffe8afe63fe48fe2cfe14fe11fe14fe1bfe38fe5afe7ffeb3fee8fe17ff4eff83ffb1ffe5ff1c0053009400d7001c016b01bc0109025902a502e90227035d038803ad03c703d903ee0300040e041f042f043f0451045e04620461045b044b042f040c04e303b3037d0348031503e202b20285025a022d02fe01cb01920157011a01dd00a100670035000f00edffcdffb9ffabff9aff8aff7bff69ff57ff42ff2eff24ff1dff1bff26ff37ff4dff6bff8affa7ffc7ffe3fff7ff0a001b002b0042005a0075009a00c500f5002c0163019901cf0101022d0251026c02830295029e02a602ae02b302b802bb02be02c402c202ba02b302a4028d02740250022702ff01ce019a016b013601ff00cc008d0048000700bbff64ff0effaffe4afeedfd89fd22fdc7fc6dfc10fcbbfb61fb03fbadfa54faf4f99bf93ff9e3f897f84bf802f8c8f792f75ff73cf71bf7f7f6def6c9f6b3f6a6f69bf690f68cf68cf691f69ff6adf6bff6d8f6f0f610f73cf764f793f7cff70cf84df895f8d7f81df966f9a4f9e6f928fa5cfa95fad4fa01fb32fb69fb8ffbb7fbe3fb01fc23fc47fc5afc73fc8efc93fc9bfca8fca0fc99fc8ffc6cfc49fc28fceefbb7fb8bfb50fb16fbe8fab0fa7ffa54fa1afae2f9aff96df92bf9eef8a5f85ff81ff8d7f798f762f728f7f9f6d2f6a3f67ff667f649f633f627f61bf61af620f622f631f643f64cf661f67df68ff6aaf6cef6e9f60ff73ff769f79bf7d7f709f842f880f8b2f8e7f823f950f97ff9b2f9d6f9faf924fa3cfa4ffa68fa73fa7dfa8bfa89fa8cfa98fa95fa94fa99fa8bfa7dfa75fa5afa39fa1cfaecf9b8f98cf94ef90ef9d7f892f84ef815f8ccf784f746f7fff6bef68df651f618f6ecf5baf58cf564f52df5f9f4c9f48df455f425f4f2f3ccf3b6f3a0f39df3a9f3b0f3c2f3def3edf3fff312f416f420f42ef432f441f45af46df48df4bbf4e4f416f54ff57ff5b9f5f6f528f662f6a1f6d4f612f754f788f7c3f7fff729f859f889f8a6f8c6f8e8f8f8f812f932f947f968f990f9a9f9cff9fff91dfa40fa65fa78fa8bfa9afa94fa94fa95fa82fa76fa72fa67fa67fa70fa72fa81fa98faa2fab1fabefabbfabafab6faa1fa91fa81fa68fa56fa4cfa3efa3cfa40fa3dfa43fa4dfa4bfa50fa5dfa64fa73fa89fa9cfab9faddfafcfa1cfb39fb4bfb5dfb6cfb70fb75fb7afb7dfb8bfba3fbc1fbf0fb29fc62fca7fceffc2ffd70fdaafdd1fdf7fd18fe2afe39fe47fe4ffe62fe7cfe90feadfed4fef6fe1dff4bff6cff87ffa3ffb8ffc2ffc4ffbeffb5ffa6ff90ff7dff6cff56ff42ff32ff1fff0cfffafee8fed7fec7feb6fea7fe9afe8dfe83fe7bfe71fe64fe52fe40fe2cfe12fef6fddbfdc1fdaefda3fda1fdb0fdcbfdedfd1bfe50fe84febbfef0fe1cff43ff65ff81ff9dffb5ffccffeeff180045007e00c3000d015d01b10106025c02ae02f8023f038303c003f503270457048104a504c604e704010517052d0543055405680581059a05b805db05fa051b063b065406670671066b065b063f061806f005c40593056f0553053c0539053e05420555056b05770587058d05810578056805480530051805fd04f604f404f0040405200538055f058805aa05d405fa0516063c065b066e068e06a806b706d106e606f00608071e072a0743075d0773079b07c607ee0726085f089208cf0805092c09520969096e09720968094f093c0925090909fc08f308ed08fc080e091d093e09570964097a09870981097e096f09500939091709e908ca08a60879085f08460827081d081208020808080b0805081008120808080c080308e907dd07c807a407930781076907680769076a078607a507c007f40727084e088608b608d6080209230933095309690971098b09a409b809e609150a400a870ad20a120b660bb60bf30b3a0c780ca30cd20cf00cfb0c100d1c0d190d240d290d230d2f0d3a0d3c0d4d0d5a0d600d760d820d830d8e0d890d720d650d450d100de10ca40c580c190cd00b800b470b0a0bc90aa20a7b0a4f0a380a1e0afa09e709cb09a3098b09670935091209e308a808800851081c080208e807cd07d307da07df0703082808450876089f08b608d808ee08f508070910091109250939094c097709a109c709030a3b0a6b0aa80adb0a020b320b530b630b770b7b0b6e0b680b560b380b240b080be80ad60ac00aab0aa70a9d0a8f0a8d0a820a6b0a560a310afd09cc098c094109fb08a6084b08fe07a7074e070907c0067a064c061c06ef05da05c205a6059b0587056805540533050305df04b1047e045e043f041f04190419041a0431044c0465048e04b504d404fd04200539055b0578058e05ab05c105d305ec05000610062906450663068c06b906e6061a074a0773079b07b807c907d307cd07b907a30782075b0734070807dd06bb069b067c06630647062d061706f905d405ad057b053c05f504a1044304dd036c03fd0291022202be0163010d01c500840042000800d0ff8eff4eff0effc4fe7bfe32fee0fd95fd4ffd04fdc1fc87fc4bfc13fce7fbbffb9ffb88fb7bfb77fb79fb83fb95fba8fbbafbcbfbd5fbddfbe1fbdcfbd8fbd9fbd9fbdefbeffb05fc21fc47fc70fc9dfccefcf9fc26fd50fd6bfd84fd9bfda4fda9fdacfda0fd93fd89fd74fd62fd56fd42fd33fd2efd20fd13fd0afdf4fcd9fcbbfc8dfc5afc22fcd6fb86fb38fbdafa7afa21fabbf95af905f9a8f852f80cf8c1f77ff74df715f7dff6b6f680f643f609f6bff56cf51df5bff462f415f4c8f385f35af335f321f324f322f327f33cf348f352f362f365f36bf37af37df389f3a2f3aef3c3f3eaf300f41bf444f45af478f4a7f4c0f4e3f419f539f55ef591f5a8f5c4f5e8f5ecf5eef5f8f5e3f5d2f5cff5aff596f592f574f55ef55df545f533f530f513f5f7f4e6f4b2f47cf44df4fcf3a8f35ff3f9f297f248f2e8f191f154f109f1cdf0a6f06ef03ef01ff0e6efaeef80ef3aeff8eec5ee7bee3bee0eeeceed98ed78ed45ed18ed00edd8ecbbecb6eca0ec96eca8ecacecbcece0ecefec02ed20ed24ed2aed3eed38ed3bed4fed52ed64ed8deda9edd8ed1cee4dee8aeed2eefdee2eef6aef87efaaefd6efe1eff6ef1bf027f03ff06bf07ef0a0f0d6f0f3f01bf153f16df18af1b2f1b9f1c1f1d5f1caf1c4f1cef1c2f1c0f1ccf1bff1bff1cff1c4f1bff1c6f1b1f1a2f19df184f179f181f171f16ef17af16df165f166f14af12ef117f1e4f0bbf0a3f07df06cf073f070f07ff0a6f0c0f0e0f009f11ef131f145f13ff13ff147f13ef141f152f157f170f19cf1baf1e4f11df248f27df2bcf2e7f21bf358f37ff3adf3e4f308f434f469f48af4b5f4eaf410f540f578f59af5c8f502f624f651f688f6a9f6d5f60af728f74cf77af790f7a8f7c1f7c1f7c5f7cdf7c3f7c5f7d4f7d8f7ecf70ff829f854f887f8a5f8c5f8e5f8ecf8f1f8f1f8def8d0f8c8f8b7f8b5f8bff8c3f8d3f8eff802f91bf937f94bf966f982f996f9b2f9d2f9ecf910fa38fa55fa76fa97faaffaccfaeafafffa1cfb3ffb62fb8ffbc2fbf4fb2efc6bfca3fcdffc18fd4afd7ffdaffddbfd08fe2ffe53fe7efea5fec8fef4fe24ff56ff90ffcdff10005c00a500ec00300169019a01c401e101fa0110021f0233024f026c029102bf02ee0224035d038d03be03ee0312043604590472048e04a704b604cb04dd04e304ef04fa04fc040605140520053d055d057905a405cf05ed05120630063b064d0659065206510651064a06510658065c0674068c069c06bf06e60603072d07550774079f07c607df0700081808220835083f083f085208650873089608bc08e1081a094e097709b109e4090a0a3d0a660a810aab0acd0ae20a080b250b310b4c0b600b660b830b9e0bad0bd60b080c2f0c680ca10ccb0c030d2e0d400d560d5d0d4c0d470d390d1d0d180d170d110d240d350d3e0d640d850d970dbd0dd80de40d060e1e0e220e3a0e440e390e3e0e370e1d0e1b0e120efc0d050e110e150e3c0e670e860ebf0ef30e140f460f6a0f770f950fa70fa20fb50fc40fc30fdc0ff10ffc0f241047105c109010c110e1101b114a1161119011af11af11c311cb11b911bb11b511a011a611a8119e11b111be11bb11d011da11cf11da11d711c011c011b0118f1186116f1142112811fb10bd10931058100e10e10fb00f7d0f6e0f5c0f460f4f0f500f400f430f320f090fee0ec10e7f0e530e1f0ee20dc20da00d7b0d780d730d650d750d800d7f0d960da50da70dba0dbf0db50dbd0db60d9b0d960d870d6b0d6a0d670d5a0d6d0d800d8b0db20dd40de50d070e1e0e200e300e320e1f0e180e050ee60dd70dbb0d940d830d660d410d370d2a0d140d190d190d0f0d190d170d060dff0ce30cb10c8c0c520c050cce0b8f0b480b1e0bf40ac90abc0aac0a930a930a880a6f0a6b0a5d0a3d0a2f0a180af309da09b90991097809510922090909eb08ca08c108b808b208c608d508e20805091f0930094b09570957095f0955093f09370925090b09ff08ec08d608d608d608d508e708f90809092809430950095d095f094f0939091109de08aa086e0833080408d207a7079007790761075707440725070907e306ad0675063206e7059c054905f404a60452040004b7036d032503e802a90274024b021d02f401d301aa0180015b012801f000bc007c003d000500c5ff8aff5dff2eff08fff4fee2fed9fedefee2feedfe02ff12ff23ff39ff45ff4cff55ff54ff4cff44ff3aff32ff31ff33ff3cff4dff64ff82ffa3ffc2ffdffff7ff090016001800170013000500f5ffe8ffd3ffbcffa9ff8fff73ff5bff3dff20ff06ffe7fecbfeb8fe9dfe7ffe66fe43fe19feedfdb5fd75fd33fdeafc9dfc57fc12fcd2fb9ffb75fb53fb3efb2efb22fb1afb0ffb03fbf4fadcfabcfa9afa72fa48fa22fafef9dff9cbf9c1f9c2f9d0f9e5f901fa28fa4ffa77fa9dfab9fad3faecfaf8fa00fb0cfb0ffb15fb24fb29fb33fb48fb51fb5ffb77fb81fb8afba0fba7fbb0fbc6fbc9fbcafbd5fbcbfbbcfbb1fb8dfb64fb41fb07fbc9fa97fa56fa1afaeef9bbf98ff971f945f91ef900f9cff89bf86ef82bf8e0f79bf744f7edf6a1f64cf600f6c4f581f547f521f5f7f4d3f4bdf49ef481f46ff453f435f41ef4fdf3dff3c6f3a1f382f370f355f341f33ff335f335f347f352f36af395f3b5f3dff318f446f476f4acf4cef4f1f416f522f530f545f545f54ff568f573f58af5b2f5d2f503f642f66df6a1f6dcf6fef620f740f741f743f747f730f71ef715f7f8f6e4f6dcf6c4f6baf6bdf6acf6a0f69cf683f66cf65bf632f60df6eff5baf58af566f531f503f5e1f4acf47ff460f42ff404f4e9f3c1f3a1f390f376f363f35ef34df343f344f336f329f326f316f308f304f3f6f2f2f2faf200f314f334f351f382f3bef3ecf322f462f491f4c4f4fbf41ef544f570f58af5a7f5cff5ecf510f63ef663f68ef6c3f6eef61ff758f780f7a8f7d3f7e7f7fbf712f812f812f816f806f8f8f7f2f7d7f7c2f7b9f79ef788f77cf75ef746f736f711f7f2f6dcf6aef681f65ff628f6f0f5c1f582f547f517f5daf4a5f481f456f437f426f40bf4fdf3f9f3e4f3d5f3cdf3b3f39ff393f375f35ef355f347f344f34ef352f369f38ef3acf3d7f30ef439f470f4adf4d9f40df546f56bf597f5c9f5e8f511f642f665f693f6cdf6faf631f775f7abf7ecf733f869f8a6f8ebf81af94ef988f9abf9cff9f8f90cfa22fa39fa3cfa44fa4ffa49fa49fa53fa53fa5efa72fa7bfa8dfaa1faa7fab3fabdfaaefa9efa8dfa68fa44fa23faf5f9cff9b2f98ff979f971f962f95af95af950f94bf94af93cf931f926f90ef9faf8e8f8cbf8b5f8a7f893f887f88bf88ef89bf8b0f8c6f8e8f811f933f959f983f9a7f9ccf9eef906fa24fa44fa5cfa78fa96fab2fad8fa00fb25fb55fb8bfbbefbfcfb3efc79fcbdfc03fd3dfd79fdb1fdd9fdfefd1ffe2ffe3efe4cfe52fe5cfe6dfe7afe8bfea5febafed4fef1fe05ff18ff28ff2cff2cff29ff17ff04fff0fed2feb4fe98fe77fe5bfe43fe27fe0ffefcfde6fdd5fdc4fdaffd9efd8ffd7afd64fd4efd33fd18fdfdfce4fccdfcb6fca6fc9cfc93fc90fc93fc98fca9fcc2fcdafcf6fc18fd3bfd5cfd7dfd9afdb6fdd3fde9fdf9fd0cfe21fe39fe56fe7dfeaffee9fe28ff6cffbbff090051009900da000b0138015f0177018c01a301b501c901e001f9011a023c025c028402ac02cc02ef0211032a0341035403600369036a0365035f03520340032d031403fd02ea02d502c802bf02b402b302ba02bc02c002c502c502c502bf02b002a00287026a0254023b02200211020502fd0104020f0220023e025a0274029702b202c702e002ee02f402ff02030302030c03170322033c035a037703a103d203ff03330468049904cd04fe042705520576059005ab05c005ce05df05ed05f105fe05100621063b0659067a06a606d006f606280752076c078a07a007a507aa07a4079007820772075a074b073f07340738073b073e0750076007690779078207830785077b0768075d07460726071007f706db06cf06c106b306b706ba06b906c806d206d406e406f106ef06f506fa06f806fd06f906ed06f206f306ee06f906000703071b07320745076c079207af07db0701081d0844085f086c088408930893089f08a708a808bb08cd08db08fe08220941096b098f09ad09d609f609080a1f0a2e0a2e0a330a310a270a280a220a160a190a170a100a1d0a280a2d0a410a510a590a6c0a760a730a7b0a780a670a600a500a370a2a0a180a010afd09f409e709f009f309f109030a100a130a250a2f0a2e0a3b0a3d0a320a370a320a230a240a1c0a0d0a140a170a130a230a330a3d0a580a6d0a7b0a960aa60aaa0abb0ac00aba0ac10abe0ab10ab50ab40aab0aba0ac40ac90ae70a010b110b350b530b660b870b9e0ba40bb70bbf0bb90bbf0bba0bac0bb10bb00ba80bb70bc50bca0be40bfc0b0c0c2d0c460c530c700c840c8b0ca10ca90ca10caa0caa0c970c920c890c740c6e0c610c4b0c4d0c4b0c420c4c0c510c4c0c590c5b0c4f0c500c400c1c0c0b0cef0bc00ba30b800b530b3c0b200bfc0af00ae10ac70ac30ab80a9e0a950a800a5f0a500a320a060aee09d009a7099309790959094e093d092a092e092b0922092e0933093009410945093d0947094a0943094c094b094009440945093e09440948094909570962096d098909a109b309d109e809f6090a0a130a100a140a0b0af809ef09db09c309bc09b209a309a509a509a109a809a4099609940984096609510932090709e308b9088808610832080108dd07b00781075f0731070107e006b7068c066c0644061b06fd05d405aa058c05620532051005e404b40492046c0444042b041304fa03ef03e703dd03dd03da03d403d403ce03bf03b703ae039e0394038f038b0391039903a403ba03d203ea0306041e04310442044f0457045e045c045704580454044e044f044a0442043d0433042804230416040604f903e803d603c303ab039203760350032903f902be0283024502fc01b50170012501dd00990055001800ddffa1ff6aff30fff1feb3fe70fe26fedefd95fd48fdfffcb7fc6efc2bfceefbb6fb85fb57fb2dfb0afbe8fac8faaefa94fa77fa5ffa47fa2efa1cfa09faf5f9eaf9e3f9dcf9dcf9def9e1f9ebf9f5f905fa1bfa2bfa3efa5bfa6ffa82fa9dfaaefabbfad0fadafae0faeafaeafae7faebfae5fae2fae9fae6fae4faedfaebfae8faecfae0fad2fac8faabfa8bfa6efa3cfa09fae1f9a8f96df93df902f9ccf8a1f868f835f80ef8d9f7a7f77ff744f70cf7e2f6a4f663f630f6eff5aff57af53bf500f5d5f4a0f46ff44df422f400f4edf3d1f3bff3b9f3a5f39af3a0f395f38ef397f38ff38bf397f393f395f3a8f3abf3b6f3d1f3e1f3faf324f440f463f492f4aef4cef4fcf414f52bf54bf557f568f582f587f595f5aef5b3f5c2f5dff5e4f5f2f50cf60bf60ff620f616f60ef610f6f3f5d7f5c8f59ef576f55bf526f5f6f4d5f4a0f470f44ef419f4ecf3cff39bf36ff351f31bf3eaf2c8f28ff25af231f2f2f1b9f191f155f11ef1f8f0c4f099f07ef056f03bf032f019f00bf00ff005f000f00af004f006f013f011f015f025f027f035f051f05ef077f09ef0baf0e2f019f13df16cf1a8f1cff1fcf134f257f282f2b6f2d2f2f6f225f33ff366f398f3b1f3d8f30bf423f446f477f48df4adf4d9f4e7f4faf41bf521f52af53cf535f534f53bf52bf523f523f50df504f507f5f2f4e9f4eef4dff4d7f4d9f4c9f4c0f4bef4a7f494f489f46ef45bf44df430f41df414f400f4fdf304f4fef307f41cf421f431f44ef45cf472f48ff49ff4b5f4d5f4e8f405f52cf547f56cf599f5bdf5edf524f64df683f6c2f6f3f62ef771f7a7f7e7f72cf85ff899f8d8f809f944f97ff9a9f9dcf914fa39fa68fa9cfac3faf1fa24fb48fb71fb9bfbb7fbd7fbf4fb02fc14fc26fc28fc2dfc36fc34fc37fc3efc3cfc3efc44fc43fc48fc4ffc4dfc4bfc4afc43fc3cfc34fc26fc1cfc11fcfffbf4fbeafbdbfbd2fbcefbc8fbc9fbcefbd1fbdcfbecfbfbfb0ffc23fc36fc51fc6bfc82fc9dfcb7fccefceafc06fd21fd41fd64fd87fdb4fde0fd0cfe40fe74fea7fedffe14ff47ff7cffadffd9ff080033005c008700ae00d400fd0026014e017a01a601d001f8011d02440269028802a902c802dd02f3020a031b032b033d034903560366037003790385038d039903a803b203be03ce03d903e403f003f503fd030604030405040c04070406040d040f04150420042a043d045304610478049104a104b704cd04dc04f00401050a051e0530053d0557056e057c059805b805cd05ec050e0628064c0670068d06b306d706f30619073a0750076f078b079e07b607c807d307e907fc0708081f08340843085b086f087c089308a208a808b908c208c208cc08ce08c808d108d408cc08d408d808d008d408d408c808c908c608b308ab08a208900887087c086b0867085d084d084a084208340835082e082108250821081708220823081c082c083708360846084f084c08590861085c0867086d086a087708800881089408a408ad08c608d908e208fa080b091209260934093a094c0959095e0970097a097d0990099a099909a409a7099e09a309a1099309950990097e097b097509680966095f094e0948093e09290920091309fd08f108df08c708bf08b408a10899088d087908710864084e0844083608210818080a08f807f307e907dd07e007da07ce07d307d007c507c807c407b807be07bd07b707c307c907c707d607de07df07f007f807f80707080a080608100810080808120814080e08150814080d0812080d0800080008f707e807e207d407c407c007b1079f079c07910780077807660750074707350718070207e806c806b30695066f06550637061006f105cf05a9058c056a05440529050905e604d004b7049a04890476045f0451043e042a041e040b04f403e903d903c403b903aa0398038f038303750371036a0361035f0359035303550353035003560359035a03620367036c0377037e0383038c038f0393039b039e039f03a403a2039d039c0395038a037f037203610350033a0323030e03f402dc02c702b002990284026c02510238021d020102e301c1019f017b0152012a010101d300a8007e0050002400faffcdffa3ff7bff50ff2aff08ffe3fec0fea1fe82fe66fe4dfe32fe1afe06feeefddbfdccfdbefdb5fdadfda6fda5fda6fda6fdabfdb4fdbafdc2fdcafdd0fdd8fde1fde5fde9fdeffdf4fdfcfd04fe0efe1bfe26fe31fe41fe4dfe56fe64fe70fe7bfe88fe8ffe93fe99fe9bfe9bfe9cfe97fe8ffe88fe79fe66fe54fe3bfe1ffe06fee6fdc5fdabfd89fd67fd4afd24fdfefcdefcb6fc8cfc67fc3afc0dfce8fbbbfb8dfb6afb43fb1efb02fbe5facafab2fa94fa7afa63fa45fa28fa0ffaeff9d2f9bcf9a2f98ff980f96ef965f966f960f960f96af970f97af98af996f9a9f9c0f9d3f9eff90efa26fa42fa60fa76fa92faaefabefad4faeefafbfa0afb1ffb2dfb3ffb53fb5dfb70fb85fb8afb95fba7fba9fbacfbb4fbaefbacfbb0fba7fba2fba5fb99fb8ffb8ffb80fb70fb65fb4bfb30fb19fbf3faccfaabfa7efa52fa2cfafbf9ccf9a5f974f946f920f9f2f8c8f8a7f87ef859f83ef81df8fff7ecf7d5f7c2f7b3f79df78cf781f76df75bf74ef73cf72cf725f71bf716f718f719f720f72df739f74cf761f771f789f7a3f7b5f7d0f7f0f709f82bf854f875f89df8ccf8f5f826f959f980f9adf9ddf900fa24fa4cfa68fa86faa4fab9fad3faecfaf9fa0afb1efb25fb30fb3efb3efb43fb4afb46fb47fb4dfb44fb40fb40fb37fb30fb2afb18fb09fbfafadffac7fab2fa92fa75fa5bfa38fa1bfa01fadff9c5f9aff98ff977f967f94df938f92bf919f90df908f900f9fff803f906f912f922f932f94bf965f97cf99bf9bbf9d7f9fbf91ffa3efa65fa8cfaacfad3fafbfa1cfb44fb6efb93fbc0fbedfb14fc44fc76fca2fcd6fc0dfd3cfd6efda1fdccfdfafd26fe49fe70fe93fea9fec1fed9fee8fef6fe02ff07ff0dff10ff0bff09ff04fff5fee9fedcfec8feb7fea5fe8dfe79fe67fe52fe40fe30fe1dfe0ffe01feeffde0fdd4fdc3fdb1fda0fd8efd7efd6afd55fd43fd32fd1ffd10fd01fdf3fce9fce0fcd9fcd8fcd9fcddfce6fcf0fcfffc14fd2bfd45fd62fd7ffd9efdc0fde2fd07fe2cfe4efe74fe9afebbfedefe05ff26ff48ff6eff91ffb5ffdbfffdff1f00430066008800ad00cd00ee0012013301520173019201b201d401f201120231024d026b0285029902ab02bb02c502cf02d502d402d402d402cd02c702c202bb02b502b002ab02aa02a802a402a302a0029c029f02a1029f02a402a702a602ad02b402b602be02c402c502cd02d302d302dd02e502e502ed02f802fd02070312031a032a033b0346035a03710382039c03b903d003f10314043004530476049504b804d804f1040d05280539054c055f056a0573057c0583058a058e058e059005920591059105920590058e058c0588058705830580057e05790571056c05620556054c053d052a0519050305ea04d504bb04a0048a046f0453043c0421040304eb03d203b803a50392037f03720365035b035a03560354035a035a0358035f035f0359035a0355034b0347033e0332032e0326031c031c031a03140317031803150319031c031d0327032d032e033a0345034b035a0367036f037f038b039203a103ab03ae03b803c003c203c803cd03cd03d303d403d203d803d803d403d903dc03dd03e603ed03f203020411041e0436044b045c0476048d049d04b504ca04d804ea04fa0402050f0519051e0527052e05300538053c053d054805500552055c0567056f057e058a059305a205ac05b305c005c805cc05d505da05db05e105e305e005e205e105dc05da05d205c505bb05ab05970585056d055405400527050f05fd04e804d404c804ba04ac04a30497048a048304770467045c044e043b0429041404ff03ea03cf03b20399037c035d03410324030703ed02d102b602a1028c027702670257024602380228021b020f02ff01f201e701da01cd01c101b301a50199018801760164014e01380122010801ee00d400b8009f0087006d00580043002b0017000500f2ffe3ffd5ffc4ffb8ffaeffa0ff94ff88ff78ff69ff5aff45ff30ff19fffcfee0fec4fea3fe84fe69fe4cfe33fe1dfe08fef7fde9fdd9fdccfdc2fdb6fdaefda7fd9ffd98fd95fd93fd92fd96fd9cfda2fdadfdb8fdc3fdcefdd9fde1fdebfdf5fdfbfd02fe0bfe15fe1ffe2dfe3cfe4efe63fe78fe91feaffeccfeeafe0dff2eff50ff76ff9cffc1ffeaff120037005e008300a400c400e000f7000e01220130013f014e015901640171017c01870193019c01a601ae01b301b801bc01bb01b901b801b401af01ab01a6019f0198018f01830176016701550141012a011101f700db00bd009f0081006200430025000600e8ffcbffaeff95ff7dff67ff54ff44ff36ff2bff22ff1bff14ff0cff02fff8feeafedbfecafeb7fea2fe8dfe77fe63fe50fe3dfe2dfe21fe12fe04fefbfdeefddffdd4fdc5fdb6fdaafd9afd8cfd82fd75fd67fd60fd53fd43fd3afd2afd15fd03fdeafccefcb4fc92fc6efc50fc2dfc06fce5fbbdfb94fb73fb4bfb1ffbf9facefaa1fa7dfa53fa29fa0afae8f9c5f9adf992f977f962f94af92ef918f9fcf8ddf8c1f8a0f880f864f845f828f811f8f9f7e5f7d7f7c8f7c0f7bcf7b7f7b8f7bdf7bff7c9f7d7f7e4f7f9f711f828f848f868f886f8aff8d8f8fbf828f957f980f9b1f9e3f911fa47fa7cfaaefae9fa23fb57fb95fbd2fb08fc47fc85fcbdfcfffc42fd80fdc6fd0bfe4cfe96feddfe1eff65ffa9ffe4ff22005d009000c500f4001d0148016f019001b601d601f2010f0229023e0254026802780289029602a302b102bc02c702d402dd02e702f002f502fa02fd02fa02f902f602ed02e602de02d202c802bf02b202a8029d028f02830276026402550248023702270219020c020002f601ef01e901e301df01dd01d701d201ca01bf01b301a4018f017b01640147012c010e01ec00cd00ab00840061003a000f00e9ffbdff8bff61ff31fffafecbfe97fe5dfe2bfef4fdb6fd81fd45fd02fdc9fc89fc41fc02fcbefb72fb30fbe9fa9bfa57fa0efac2f980f938f9eff8b1f86ef82bf8f2f7b7f77cf74bf719f7ebf6c4f69cf67af660f643f62df61ef60df602f6fcf5f4f5f2f5f5f5f4f5fcf508f60ff622f638f64bf66af68df6aef6dcf60df73cf77bf7b9f7f5f741f88cf8d2f827f97cf9cbf927fa80fad5fa36fb94fbebfb51fcb2fc0dfd74fdd7fd33fe9cfefffe5dffc6ff27008400ec004b01a5010a026602be0220037b03d20331048704dd043a058c05de0534067e06c806150755079507d6070b08410876089f08cc08f80818093c09600979099609b209c309db09f009fa090d0a1c0a210a2e0a380a390a420a460a420a430a3d0a300a290a180a000aed09d209b209960973094c092a090009d508ae087e084d082008e807af0778073607f506b6066c062506e10591054705fe04aa045c040f04b4035e030703a3024402e20174010d01a3002e00c3ff57ffe1fe76fe0afe96fd2cfdc1fc4ffce8fb7efb0efbabfa45fadaf97bf91af9b6f85ef802f8a5f753f7fcf6a5f659f607f6b7f573f529f5e4f4abf46ef438f40df4dff3b9f39ef37ef367f35bf349f341f341f33df345f353f35df376f394f3adf3d6f303f42af461f49bf4d0f413f557f597f5e6f534f67ef6d8f631f786f7ebf74df8adf81df989f9f4f970fae6fa5cfbe4fb65fce6fc78fd02fe8bfe23ffb0ff3c00d5005f01ea018102080391032604ac043505cb055306de067407fa078508170998091c0aa60a1e0b980b170c840cf50c6a0dcd0d360ea10efa0e590fb70f04105410a210de101d1157118011ad11d311e911051217121b122512241216120c12f711d611ba1191115e113311f810b7107e103610e80fa20f4b0fef0e980e300ec30d5b0ddf0c610ce80b5d0bd20a4e0abb092a09a1080a087807ed065406c1053405980401047103d2023902a60107016f00ddff40ffaefe20fe8afdfefc77fce7fb63fbe1fa59fadcf95ff9dcf865f8ebf770f700f78ff61df6b7f550f5eaf492f437f4e0f398f34bf304f3ccf28ef256f22bf2faf1cff1aef186f165f14ef12ef117f109f1f4f0e9f0e9f0e3f0e7f0f6f000f117f135f14ff177f1a4f1ccf103f23ef275f2b9f202f348f39cf3f1f346f4aaf40df570f5e3f553f6c4f644f7c1f740f8cef856f9e1f97bfa0dfba2fb47fce0fc7dfd29fec9fe6dff1f00c4006f012902d40287034804fa04b20577062a07e207a3085109020ab80a590bfe0ba70c3a0dd20d6e0ef60e830f131091101311961106127a12ea124613a613fd1340148614c214eb141615371547155b1562155b155a1549152b151215e914b41483144014f213a9134c13e61287121212961123119a100d10890ff20e580ec90d270d860cf00b460ba00a060a5909af0810085f07b2060f065905a90403044c039c02f80143019900faff4fffaffe1afe7bfde9fc60fccdfb49fbcbfa43fac9f954f9d6f866f8f9f786f71ff7bbf653f6f9f5a0f544f5f9f4adf45ff421f4e1f3a1f36ef337f300f3d4f2a3f272f24ef221f2f6f1daf1b5f194f182f16af158f154f14bf14af155f159f165f17bf189f19ef1bbf1d0f1ebf10df228f24df277f29cf2ccf203f335f375f3bbf3fdf34df4a0f4f1f44ff5aef50bf676f6def645f7baf72cf89ef81df997f913fa9efa21fba6fb3afcc5fc52fdeefd80fe14ffb6ff4b00e30087011d02b5025803ec0381042005af053f06d8066207ef07830807098f091c0a990a190b9d0b0f0c830cf60c580db90d170e640eb20efa0e310f6a0f9d0fc20fe90f0a101e10371047104b105410511043103a1023100110e30fb60f7f0f4c0f090fc00e7c0e290ed00d7f0d200dbe0c620cf70b8b0b270bb20a3b0acb094a09c9084e08c3073807b506230695050f057c04ee036a03db025302d2014601c2004400baff3affbefe36feb7fd3cfdb7fc3bfcc2fb41fbcbfa57fadcf96ef901f98ef828f8c3f75af7fff6a2f643f6f1f59bf543f5f9f4aaf458f414f4caf37ef341f3fcf2b8f283f249f211f2e7f1b7f18bf16ff14cf12bf118f1fcf0e6f0daf0c4f0b4f0aef09ef096f099f092f094f0a3f0abf0bef0dcf0f2f016f142f166f198f1d2f101f23bf27bf2b2f2f5f23af377f3c1f30df451f4a5f4faf447f5a7f508f663f6cef639f79df711f882f8edf867f9daf946fabffa33fb9efb17fc8afcf7fc71fde5fd54fecffe43ffb4ff3100a50014018d01fc016702d8024003a3030b046a04c60426057b05cf0527067606c30614075d07a507ef0730087208b508ef08280960098f09bd09e709080a290a460a5a0a6d0a7a0a810a890a8d0a8c0a8c0a870a7e0a780a6b0a5b0a4c0a330a170afc09d409aa0980094a091209db08990857081608cc0783073d07ed069f065206fa05a7055105f00492043304c8036203f80283021602a6012d01bc004900ceff5effeafe6ffefffd8cfd12fda4fc31fcb5fb46fbd5fa5afaebf97af903f998f828f8b6f752f7e9f67ef623f6c5f565f512f5bef46bf424f4d8f390f354f312f3d3f2a1f269f234f20cf2ddf1b4f198f176f15cf14ef139f12ef12ff129f12cf13af140f151f16bf17af194f1b5f1ccf1eff119f238f262f294f2bcf2f0f22cf35ef39cf3e1f31df466f4b3f4f5f444f597f5dcf52ef682f6c9f61bf770f7b9f70cf862f8aef805f95df9aff90afa66fabbfa19fb76fbcefb2dfc88fcdefc3bfd93fde8fd43fe98feebfe46ff9cfff1ff4c00a300fc005a01b3010d026c02c4021e037c03cf0324047f04d00421057405c0050e065d06a406ee0639077d07c307080847088a08ca08040940097909aa09dd090d0a340a5e0a820a9e0aba0acf0ade0aef0af90afd0a030b020bfc0af60ae90adb0acc0ab20a960a7a0a500a250af909be0983094809fe08b6086f081a08c80779071d07c60670060e06b3055805ef048b042904b8034c03e2026d02fd018d0111019d002d00b5ff43ffd5fe5efef1fd88fd19fdb2fc4efce5fb86fb2dfbcdfa74fa21fac9f979f92df9e1f89cf859f818f8e0f7a9f775f74af724f701f7e4f6c8f6b2f6a4f695f68af686f680f67ff686f68af693f6a3f6b1f6c7f6e3f6fcf61df745f76af797f7c8f7f7f72df867f89df8d9f817f951f991f9d1f90cfa4efa8ffacafa0dfb50fb8efbd3fb18fc5bfca5fcedfc36fd86fdd3fd1efe6ffebefe0dff5effabfff9ff48009100de002f017801c60117026002b00204034f03a103f5033e048d04df0425057305c00501064c069906d7061d076607a507ed0736087408ba0800093c098109c509fe093d0a7c0ab00aea0a1f0b4a0b7b0ba70bc70bef0b120c2b0c490c610c700c870c970ca00cb00cb90cba0cc20cc10cb90cb60ca80c960c8a0c6e0c4c0c300c080cdc0bb30b7b0b430b120bd20a900a540a090abf097c092809d40885082708c80770070a07a5064506d9056f050c059d043104ce036303fc029a023102cc016c010601a2004600e5ff83ff27ffc8fe6afe10feb7fd63fd12fdbffc73fc2dfce8fba9fb71fb3dfb0cfbe1fabafa99fa7dfa65fa50fa3efa30fa25fa1ffa1efa1efa22fa2bfa36fa45fa5bfa70fa89faabfaccfaedfa19fb43fb6bfb9cfbcdfbfcfb33fc67fc9cfcd8fc11fd4bfd8efdccfd0cfe55fe96fed9fe27ff6dffb2ff000047008c00d8001b015c01a101df011b025b029302c902020334036903a103d10306043f046d04a104da0408053a056f059805c705f7051a0642066c068b06ab06cd06e806070725073c07590775078907a207ba07cc07e307f6070208140822082a0838084308470852085b085e0867086c086d0874087608720874087108680865085a0849083d0829081008fb07de07bb079d0776074d072807fa06cb06a20670063e061106db05a50573053805fc04c2047e043904f403a60359030c03b4025f020c02b1015601fe00a0004500e9ff89ff2dffd0fe6ffe14feb6fd54fdf8fc9cfc3efce7fb8dfb36fbe6fa93fa40faf9f9b3f96bf92cf9eef8b2f87df847f815f8eaf7bef796f773f750f732f71af701f7eff6e4f6d6f6d3f6d8f6ddf6ecf602f717f736f75cf782f7aef7e0f711f847f881f8bbf8faf838f978f9c0f907fa4cfa9afae6fa30fb83fbd3fb22fc7afccefc1ffd76fdcbfd1efe76fec9fe1bff73ffc1ff10006500b100fa004b019401d90127026a02a802ed022b036603a403d90309043a0462048704ae04cc04e50400051405240536054805570562056a0576057f0584058c05920592058f058b0584057b056d055e0550053c0522050a05ef04d304b704970478045b0438041504f403cf03ab038903660341031b03f202cc02a7027e0256022e020002d701b101830155012a01fd00d200a4006f003f000e00d5ffa1ff6bff2ffff5febafe7afe3dfefdfdbafd7dfd3efdfbfcbffc7efc3cfc02fcc4fb82fb49fb0cfbcafa8ffa4efa0cfad0f98cf945f909f9c7f883f847f806f8c2f788f74cf713f7e0f6a7f674f64bf61cf6f0f5cdf5a7f586f56df54ff537f526f50ff502f5fdf4f2f4eff4f2f4f0f4f8f408f512f526f540f554f56ff592f5b2f5daf506f62ef660f696f6c7f603f744f781f7c8f711f859f8abf8fdf84bf9a4f9fef952fab0fa0cfb62fbc3fb1efc73fcd4fc30fd82fdddfd36fe86fedffe32ff7dffd3ff24006b00ba00050147019101d701130253028f02c602ff0231035b038703af03d003f0030c0423043904490453045d04620463046404600456044704370424040e04f703db03bb039e0380035b0337031003e702c1029d02720247021c02ed01c1019301620135010701d1009e006e0038000500d2ff9fff6fff3eff0bffddfeaffe7efe54fe2afefffdd8fdb3fd8cfd6cfd4afd23fd04fde7fcc6fca9fc8dfc6efc52fc36fc17fcfefbe4fbc9fbb3fb9afb7efb68fb4ffb37fb24fb0cfbf4fae3facafab2faa2fa8dfa76fa69fa54fa3ffa35fa23fa0efa06fafaf9e7f9dbf9cdf9bff9b6f9a8f999f991f983f976f96ef961f955f950f947f940f93df939f939f93df93ef944f94ff956f963f975f983f995f9abf9bef9d7f9f3f90afa27fa49fa64fa85faadfad0faf7fa23fb4dfb7afbaafbdafb0cfc41fc75fcadfce6fc1bfd57fd94fdcffd0efe4cfe87fec9fe0cff49ff8bffcbff070047008900c800090145017e01bb01f5012a0262029502c402f50223034c0374039903bd03e103030422043f04590473048a049c04b004c004c904d304dc04e004e104de04d804d304c804ba04af04a1048c0479046504500439041e040504ef03d203b4039703770359033e031b03f902dc02ba0298027a02570237021e020002e001c601aa018f0179015e01460134011e010501f400e200cc00bc00ae009f00920086007b0073006c00660063006000600062006400660069006c0073007c00820088008e0093009c00a800b000b700c000c900d400e000eb00f800060112011e012901340140014c0154015e0168016f0174017c01830188018d019101960199019c019e01a001a101a201a501a501a1019e019a01960192018d0185017f0176016d0167015e01550151014b0143013c0136012f012b01260122011f011901130112010f010a0109010801040106010a010a010a010e0116011e0124012b01350140014a015801670173017f018d019b01ab01bd01cc01dc01ee01ff0115022a023a0250026a0280029802b002c402dc02f8020f03230338034c036303780388039c03b003c003d303e403f103040416042204340441044a045a0467046c047804820486048f04960496049b04a104a004a304a604a604a904a904a504a704a804a304a704a7049f049e049c049604970494048c048e048e0488048c048d0488048f04970498049f04a404a704b904c404c404d304e304e804f60401050705180525052c053e054c0554056605760580059305a505b005c005cd05d905eb05f405fa050a06130617061f0621061d06210621061d061d0613060306fc05ee05da05cb05b7059b058105630542052005f904d204aa04780448041d04e703b00380034a030f03d8029b025f022502e401a40167012201df009c0053000e00cdff84ff3ffffdfeb7fe76fe36fef2fdb8fd80fd42fd0efddefca8fc78fc4efc22fcfcfbdafbb6fb9afb80fb64fb51fb44fb33fb26fb20fb1cfb1cfb20fb27fb31fb3ffb51fb64fb79fb93fbaffbcefbedfb0ffc38fc62fc88fcb6fceafc19fd4dfd89fdbefdf6fd39fe76feb1fef2fe2dff6affadffe8ff240064009d00d700150146017801b501ec011c0251028202b302e60212033f036f039703bd03eb0310043104560473048b04aa04c704dd04f10405051b052c053805470553055e056a0573057705810586058505880588058405860585057f057d05770571056f056a056505630559054f054e0547053c053405260519050d05f704e304d304ba04a1048b046d044f0435041204f203d403ad03890366033c031603ed02bb028c025d022702f201bb017c0140010101bc0079003200e8ffa0ff50fffefeb5fe63fe0bfebcfd64fd09fdb7fc5ffc01fcaffb56fbf7fa9efa43fae9f99af943f9ebf8a0f850f8fef7b9f770f726f7e8f6a7f664f62df6f6f5c0f591f560f534f512f5edf4cef4bbf4a3f491f48cf488f489f493f49df4adf4c9f4e6f409f531f55af58ff5c6f5faf53af67df6bef60bf75af7a5f7fcf752f8a6f809f96bf9c6f92efa95faf8fa64fbcefb36fca8fc14fd7afdeafd56febcfe2aff92fff5ff5f00c10020018601e20139029902ed023a038f03da0319045e049b04cf0409053d0564058b05af05cc05e805ff050f0620062c06320637063a0636062d06240616060406f105da05bb059d057f0556052d050605d504a404750440040a04d6039c0361032703e802ad0274023202f201b60173013401f600b0006f003200edffaeff70ff2bffedfeb0fe6cfe2efef1fdadfd70fd2ffde9fcabfc6cfc27fce8fba4fb60fb25fbe3fa9ffa62fa21fae1f9a8f966f926f9f1f8b2f873f83ff803f8caf796f756f71df7edf6aff675f648f610f6d9f5abf574f542f51bf5e9f4bcf49af46ff44bf430f40ef4f0f3dbf3c2f3b0f3a4f393f38cf38bf384f387f391f399f3a9f3baf3caf3e9f30bf426f44ff47cf4a3f4d7f410f545f586f5c9f506f652f6a2f6ecf642f79bf7f0f753f8b5f813f97ff9e9f950fac3fa34fba1fb17fc8cfcfcfc75fde8fd58fecffe3fffabff1f008b00f4006301c9012a029402f5024d03ab0302045104a304f00435057b05ba05f00526065a068506ac06ce06e706fd0612071f072507290725071a070e07fa06e106c706a5067c0652062406f005bb057e053d05fd04b80470042a04dd038a033b03ea0293024002ea018f013801de0081002900ceff6eff16ffb9fe5afe04feaafd4efdfafca3fc4afcfdfbaffb5cfb13fbc9fa81fa42fafef9baf982f945f90af9dbf8a7f873f849f81af8eff7cff7a8f785f76df74bf72ef71ef706f7f1f6e5f6d2f6c3f6bdf6b0f6a9f6aaf6a1f6a1f6a9f6a5f6a8f6b4f6b6f6bff6d3f6dff6edf600f70ff725f73cf74ef76af785f799f7b9f7d9f7eff711f835f851f876f89ef8bff8eaf815f93cf96cf99df9caf9fff933fa63fa9dfad6fa0bfb4afb86fbc0fb02fc3efc7bfcc3fc05fd44fd8cfdccfd0dfe5bfea1fee2fe30ff78ffbdff0c0054009900e6002c016f01bb01010244028c02d002110355039403d10310044b048604c204f60429055c058a05b805e00504062b064e06670682069c06af06c106d106dc06e706eb06ec06ed06ea06e506df06d106c106b2069c0683066a064b062b060c06e405ba059305650538050d05db04a70475043f040904d5039c0366033303f902c0028a024f021502e201ac01740141010c01d800a700750046001a00eaffbfff9cff73ff4bff2aff08ffe9fed2feb6fe9bfe89fe74fe5ffe55fe49fe3dfe3afe36fe31fe36fe39fe3afe44fe53fe5dfe6dfe7ffe90fea4febbfed3feeefe09ff23ff45ff65ff82ffa5ffcbffedff14003e0062008900b600df00070132015c018a01b701dc010502320259028002ab02d102f7021e03410365038903a903c903e70301042204400455046e0488049a04b004c504d404e804fb04040512051f05260532053d05410548054b054b05500552054f05530553054b054a05480540053f053b05320530052b0520051e051a05120512050e05060507050205fa04fc04fa04f404f904f804f104f804f704f104fd040105fb0406050c05090515051e051e052d053705380547055505590568057705810593059e05a705bc05c905d105e605f405fc0510061e062406370644064b065b0665066706760680068306900697069806a506ac06ac06b606bb06ba06c206c606c406cc06cc06c706d206d406c906cc06ce06c606c806c706bd06bf06bd06b406b506b306ab06ab06a806a006a206a0069c06a306a1069906a206a506a006a606a906a906b406b506b206bd06c206c006cb06d006ce06d806dc06d906e306e906e706ed06f006ed06f306f106ed06f306f006e906ed06e806dc06d906d306c506bf06b306a10691067f066a0656063b0622060b06e705c205a4057c05540531050105d004a704750442041404dd03a40372033a030103cd02930256022002e601a8016e013501fb00c20087004e001700ddffa6ff73ff3eff0cffe0feb2fe85fe5cfe33fe0efef1fdd2fdb3fd9cfd87fd72fd68fd61fd57fd54fd55fd54fd58fd61fd6dfd80fd94fda5fdbefddcfdf7fd19fe3ffe61fe8bfeb7fedefe0dff40ff6dff9fffd8ff0e004a008600bb00f80039017101b001f3012e026b02aa02e40221035d039003ca030404330467049b04c704f504220544056d059505b005d005f3050a0623063d064f066106730681068f0698069b06a006a406a306a2069e0695068c067f067106640651063c0628060d06f105d905ba0598057705520530051005e804c00498046c0443041e04f203c7039c0369033c031103de02ac027c0246021302df01a60170013601f900c100840042000900caff84ff48ff09ffbffe81fe40fef7fdb6fd74fd2afde7fca1fc5afc19fccefb80fb3ffbf8faabfa69fa1ffad1f98ff944f9f6f8b4f86af81ff8dff794f74af70df7c6f67ff648f607f6c5f592f558f51ef5f3f4c1f48ff46bf442f41ef401f4dbf3bff3aff393f37ff377f367f35ff360f356f354f360f365f372f387f395f3adf3cbf3e3f309f436f459f488f4bef4edf426f566f59ff5e0f527f66cf6b8f604f749f79cf7eff73bf892f8e9f838f992f9ecf93dfa98faf2fa42fb9cfbf7fb4afca2fcf9fc49fda0fdf3fd40fe97fee9fe30ff80ffceff120059009f00dd001e015b018f01c501f80121024c0275029602b802d602ea02ff0212031b032503300330032e0330032a031e0313030003ec02dc02c002a10286025f0234021402e801b40187014f011001dc00a00059001a00d2ff85ff46fff9fea2fe5afe0afeb1fd63fd0efdb2fc64fc0dfcaefb5cfb05fba9fa58fafcf99df94df9f4f896f847f8ebf78bf73cf7e4f686f637f6e0f588f53df5e9f492f44cf4fcf3aef36ff323f3d8f2a2f261f21ef2eff1b6f17df154f124f1f8f0d8f0acf088f074f052f036f02cf014f003f0feefefefeaeff1efeaefeeefffef00f010f02ef039f051f077f08ff0b4f0e4f007f137f170f19df1daf11ef255f29af2e2f220f36ff3bff301f456f4adf4f5f44ef5a9f5f5f552f6b2f603f764f7c5f717f87cf8e2f838f99cf901fa59fac1fa2afb83fbe7fb4efca9fc0dfd6ffdc6fd25fe82fed6fe31ff88ffd8ff2f008100c70014015f01a201e9012a0262029f02d60207033d036e039603c203e9030704280448046004750488049704a204aa04af04af04a8049f0495048604710458043f041f04fa03d503ad037f0351031e03e502af0275023402f701b80173013101ea009d0057000c00bbff70ff1fffc9fe7dfe2bfed3fd83fd2efdd3fc85fc33fcd9fb8bfb39fbe3fa96fa46faf5f9aff965f91bf9daf895f853f81bf8def7a9f77cf748f718f7f5f6cdf6a9f68ff670f656f64af639f62af625f61df618f61ef623f62cf63af647f65af675f690f6b0f6d6f6fbf626f758f78af7bff7f5f72ff871f8b2f8f3f83df984f9ccf91dfa6bfab5fa08fb5bfbacfb04fc56fca8fc04fd5afda9fd05fe5ffeb2fe0bff63ffb9ff13006600ba0016016801b90110026202b20208035503a103f00336047f04cb040d054e059405d0050d064a067f06b906f2061c074d078107a907d207fe0723084c0872088f08b108d308ea0805091f0934094b095d0969097c0989098d099909a0099f09a309a20999099609910985097c096d095a094c0936091d090d09f308d008b9089c0878085b0837080e08ee07c6079807750749071507ee06c006870658062706ee05ba0582054a051805db049b0468042f04f303c00386034a031803e102a9027c0248021102e701bc018d0165013c011301f200ce00ad00940076005600460033001d0014000900fbfffafffcfff9ff01000c00130025003800490067008600a000c700f200140142017601a301db01150247028602ca02030347038d03c90311045d049c04e80436057605c10512065606a106ef0633077f07cc070c0855089f08dc08240967099d09e009230a540a8b0ac50af20a220b4f0b710b9c0bc30bdc0bfd0b1a0c2a0c430c570c5c0c6b0c760c750c7a0c7a0c730c740c6b0c560c500c400c240c160c020ce10bc90bad0b890b6f0b490b1b0bfc0ad30aa00a7a0a4f0a1a0af209c4098d0961092f09f608c90895085f083308ff07c8079d076b0737070c07da06a9067f064b061a06f605c6059305700548051905f304cb04a20480045c0436041604f103ce03b503970374035d03450327031103fc02e502d302c002ac029f028e027d0276026c025c02580253024702440243023a023b023d0239023d02430246024d0255025d026c0277027e029002a102ae02c702de02ed0205032003350352036e038503a403c303dc030004210439045f0484049d04bf04e404010528054c0567058e05b205cc05ef0511062a064e0671068806a606c506da06f4060e07200738074a075507670775077e078c078f078e0795079207890787077c076d07650752073c072c071107f406da06b6069106710646061906f005be058b055b052005e704af046d043004f503ab0364032003d5028e024802f601a8015d010c01c10072001c00d0ff83ff2dffe1fe94fe3ffef3fdabfd5dfd13fdc7fc7afc37fcf3fba9fb6afb2cfbe8faadfa73fa38fa05fad2f99cf970f945f917f9f3f8d0f8acf890f875f85cf849f834f823f81cf810f806f808f807f808f811f818f821f831f840f854f86ef885f89ef8bcf8dbf8fff824f947f970f999f9c0f9f0f921fa4dfa80fab4fae4fa1cfb52fb84fbbcfbf4fb27fc61fc9cfcd1fc0bfd42fd78fdb3fde8fd17fe4efe82feb2fee8fe18ff41ff72ff9fffc5fff0ff19003c00600082009e00be00dc00f3000b0123013301420151015c0166016e016f01730175016e016801650157014a013f012a0115010401e700c900b2009300700051002900ffffdcffb1ff81ff58ff28fff4fec4fe8efe57fe26feecfdb0fd7dfd40fd00fdc9fc8bfc49fc11fcd0fb8bfb51fb10fbccfa92fa52fa0dfad0f990f94ff915f9d4f892f85bf81ff8e0f7aaf770f735f702f7c9f696f66af632f6fef5d8f5a8f57cf55cf531f509f5eef4c9f4a9f495f479f45ef44ef439f42bf424f414f40cf40ff409f40af413f414f420f434f43df44ff46df481f49af4bcf4dbf402f52ef552f57ff5b3f5def515f651f683f6bff602f73ef781f7c9f70bf858f8a5f8e8f838f98af9d1f922fa7bfac9fa1afb6ffbbefb15fc6bfcb7fc09fd60fdaefd00fe50fe98fee9fe37ff78ffc2ff0c0049008b00cd0002013c017701a601d80109022e02540279029502b302cc02dc02ef020003030308030e030b030303f902e902da02c702ab028f0273024b022302ff01d1019e016e013601fd00c800890046000a00c6ff7fff3cfff1fea4fe60fe15fec3fd7bfd30fddffc96fc49fcfafbb2fb67fb19fbd4fa8afa40fafcf9b5f971f937f9f5f8b4f87ff846f80cf8def7adf779f750f726f7fdf6dcf6bdf69ff686f66df65af64af638f62df627f61ff61ef622f621f62bf63cf646f654f668f67cf697f6b6f6d1f6f4f61cf740f76af798f7c5f7f7f729f85af896f8cff805f949f98cf9c7f90bfa52fa96fae1fa29fb6ffbbdfb0bfc5afcaefcfcfc4afda0fdf1fd43fe9dfeebfe3cff99ffecff3d009900eb003b019701ea013a029002e10230038503d3031f046e04b70403054f059105d7051f065c069d06de0614074e078807b707ea071d0844086c089508b608d708f30806091e0931093c094a0952095309570954094909420935091f090a09f008d408b7089008680843081308de07ae0777073a07fd06ba0678063606eb05a10557050505b60467040f04b90365030903b1025d020002a4014a01eb0092003b00dcff82ff2dffd1fe7bfe2afed3fd80fd31fddefc94fc4cfcfffbbafb7bfb36fbf8fabffa85fa51fa1efaeaf9c0f99bf974f954f939f91df905f9f4f8e6f8daf8d2f8ccf8cbf8cdf8d4f8def8e9f8f9f80df923f93df95bf97bf9a0f9c2f9e8f916fa44fa74faa9fadafa0ffb4efb89fbc1fb03fc42fc81fccafc0cfd4bfd94fddcfd26fe74febafefffe4eff98ffe3ff32007a00c20012015b01a501f3013a028102ce0212035803a203e60328046e04ac04eb042f056c05a805e6051b0654068f06bf06f106250752078007ae07d207fa072208420864088808a108bd08d908ec080109150923093409400946094f0953095309590956094e094d09410931092b091b090509f908e208c508b508990876085e083d081408f607d007a307800756072707ff06cf069e06740640060b06df05a905710544050c05d204a2046c0435040304c903950366032b03f302c5028e0258022b02f701c301980168013a011301e400b60094006a00420024000100dbffbdff9eff80ff68ff4fff34ff1eff0afff8fee7fed7fecdfec5febafeb2feadfea8fea8fea9fea7fea9feaffeb5febbfec4fecffedafee7fef8fe0bff19ff29ff3eff53ff68ff7fff93ffaaffc4ffddfff7ff11002900440061007c009700b100ce00ed00070121013f015a0173019001aa01c301dd01f601100229023d0255026e027e029102a802b802c802db02ea02f9020703110320032e0335033f0348034e0355035d03600363036403640367036603600360035d03560355035103460341033b0332032903200314030b030003f002e502d902ca02bd02af029f029402860276026b025c024c0240023202230218020a02fa01ee01e201d501cb01bd01b301aa019b018e0187017b016f016c01630156014f01470140013d0135012d01280123011e011b01170113010f01060102010201fd00f700f300f200f200f000ec00e900e800e300de00db00d900d500d100ce00cb00c700c300be00b900b500b000aa00a4009f009c00990091008a00860081007a0074006b0062005f00590050004b0045003c0038003200260020001c0013000a0007000000f8fff2ffecffe7ffe3ffddffd4ffcfffcbffc5ffc0ffbaffb5ffb3ffb0ffaaffa7ffa4ffa1ff9fff9cff98ff96ff93ff90ff8fff8cff88ff87ff86ff84ff83ff80ff7eff7dff7aff77ff75ff72ff71ff71ff6eff6bff6aff67ff63ff63ff5fff58ff54ff54ff4fff4aff46ff42ff3dff36ff2fff2cff26ff1eff1cff18ff10ff0bff08ff03fffdfef4feedfeecfee5fedafed6fed2fecbfec7fec1febbfeb9feb6feaefea9fea6fea1fe9dfe99fe96fe95fe91fe8ffe90fe8bfe85fe85fe86fe87fe86fe83fe81fe84fe84fe84fe88fe88fe87fe8bfe8dfe8dfe90fe92fe92fe96fe99fe9afe9cfe9efe9efea1fea2fea1fea4fea5fea5fea6fea8fea7fea7fea8fea7fea5fea2fea1fea0fe9bfe96fe94fe8bfe84fe83fe7cfe73fe6efe65fe5afe54fe4afe3ffe36fe29fe1efe15fe06fef6fdecfddbfdcbfdbffdaefd9cfd8ffd7efd6dfd60fd4efd3dfd2efd1afd09fdfdfce9fcd6fccafcb8fca5fc97fc86fc72fc63fc54fc44fc37fc27fc18fc0efcfffbeffbe5fbdbfbcefbc5fbb8fbadfba9fba4fb9cfb97fb91fb8cfb88fb84fb82fb82fb80fb80fb83fb85fb87fb8bfb8ffb97fb9efba1fba9fbb4fbbbfbc2fbcdfbdafbe6fbf1fbfbfb0afc1bfc2cfc3cfc4bfc59fc6cfc80fc91fca5fcbbfccffce3fcf7fc0dfd25fd3dfd52fd69fd7efd94fdadfdc5fddbfdf1fd0bfe25fe3ffe58fe71fe8cfea6febdfed8fef4fe09ff20ff3bff54ff6dff86ff9fffb9ffd3ffeaff010019002f004800610077008c00a300b900ce00e200f6000a011c012e014401580169017b018c019b01ac01ba01c601d301e101ed01f80100020a0215021d0223022b02320237023c024002430245024502430241023e023d023a0234022f022a0222021b0215020c020002f301e601d801c901b801a8019701840171015e014a0134011f010a01f000d700be00a40089006e00520035001a00ffffe1ffc2ffa3ff84ff66ff46ff27ff0bffecfecafeaafe8dfe6ffe4ffe2ffe12fef4fdd3fdb6fd9bfd7dfd61fd49fd2dfd10fdf7fce0fccafcb5fc9efc88fc76fc63fc4ffc3ffc30fc23fc18fc0cfc02fcfbfbf1fbeafbe7fbe3fbe2fbe2fbe0fbe0fbe5fbe7fbecfbf5fbfcfb05fc11fc1cfc2bfc3cfc4bfc5dfc70fc83fc99fcaefcc2fcdafcf5fc10fd2afd45fd60fd7efd9bfdbbfddbfdf7fd17fe3cfe5efe7ffea3fec3fee5fe0bff2bff4dff73ff96ffb9ffdfffffff2000470069008a00ae00d000f10011013001520175019401b301d001eb01080224023e025c0279028f02a802c202d902ef02060319032d033f034e03600372037f038e039d03a903b603c303cb03d403df03e603ec03f103f503f803fa03fc03ff03ff03fd03fd03fa03f603f403ed03e303de03d603cb03c103b303a6039b038d037f036f035b034a033b03260313030403ef02d802c402ad0295027e026302490234021c020202e701cd01b4019d01820166014c0131011301f600dd00c700ae0092007900610047002d001400fdffe7ffd0ffb8ffa1ff8bff74ff5fff4bff39ff2bff1eff0fff01fff2fee3fed7fecdfec1feb7feb1fea9fea1fe9bfe97fe94fe93fe94fe94fe94fe94fe96fe97fe9bfea3feacfeb5febdfec5fecdfed7fee1feecfefafe07ff14ff23ff34ff44ff53ff63ff75ff85ff97ffaaffbcffceffe2fff5ff07001a002c003e0052006300750088009900ab00bf00d200e500f8000801170129013801460156016401730181018d019801a401b101be01ca01d201d901e401ed01f301fc01030206020b02100216021a021d021e02200222022202240224022402230222021f021b02150211020f020b0207020402fd01f601f101eb01e301dc01d501cc01c301ba01b001a801a001990193018c0184017a016e0163015601490141013a01320127011c01130109010001f800f100e700dd00d500cc00c300bb00b300ad00a5009d0096008e0086007f00790075006f00680063005f0059005500540050004d004c004700430042003e003c003d003b00380038003600370038003600370039003a003c003e003e0041004500460046004a004d005000530057005d00610066006b006e007200770079007b008000850088008c008e00900095009a009d00a300a800ad00b300b600b900c000c400c600ca00cc00cd00d100d500da00e000e300e400e700ea00ed00f000f000f100f400f400f300f500f700fa00fd00fc00fb00fc00fb00fb00fd00f900f600f700f400f100f100f000ee00ec00e800e500e500e300df00dc00d900d700d300ce00cb00c900c500c100be00ba00b600b100ac00a800a3009e009a00950090008d008b008800860083007f007c0079007500730070006e006b00680064006400640063006100610060005e005b005a005b005a0058005800590058005a005d005c005b005c005e0062006500660067006800670069006c006d007000730075007700760075007700780077007800790079007b007b007a007b007c007a007900780076007400730070006e006d006a00670062005d00580053004d004a00480043003c0035002d00270022001a0014000c000300fbfff2ffe7ffe0ffd9ffcfffc5ffbbffb0ffa5ff9bff93ff8dff83ff77ff6fff69ff60ff57ff4dff45ff3dff36ff2dff23ff1aff13ff0bff04fffdfef8fef1fee9fee4fee0fedefedbfed8fed4fed0fecbfec7fec4fec3fec1fec2fec3fec2fec3fec4fec4fec5fec6fec7fec8fecbfecbfecefed3fed7fedcfee2fee7feebfef0fef4fefbfe03ff09ff10ff18ff1fff27ff2eff34ff3dff46ff4eff58ff61ff66ff6dff75ff7dff85ff8cff92ff9bffa3ffaaffb4ffbdffc5ffceffd9ffe2ffedfff6fffbff020008000d0013001a0021002a00310036003c00410047004c0050005300570059005c00620067006b006d006e006f00710072007400770077007800790077007500750072006e006d006900660064005f005d005b0054004d004800400039003200280021001c0014000d000500f9ffefffe6ffdcffd3ffcbffbfffb4ffa9ff9bff8fff85ff77ff6bff61ff55ff4aff3eff30ff23ff15ff08fffdfef0fee1fed6fecbfebcfeb1fea7fe9cfe91fe85fe78fe6efe63fe58fe51fe48fe3dfe37fe2ffe25fe1ffe17fe0ffe0afe05fe00fefbfdf5fdeffdeefdeafde5fde3fde2fde3fde6fde8fdeafdedfdedfdecfdf0fdf3fdf7fdfefd02fe07fe10fe16fe1bfe24fe29fe2ffe3bfe44fe4bfe55fe5ffe6afe75fe7dfe85fe91fe9afea1feadfeb7fec0fecbfed8fee8fef8fe02ff0cff18ff20ff28ff32ff3aff43ff50ff5bff66ff72ff7bff82ff89ff90ff99ffa2ffa8ffafffb8ffbdffc1ffc6ffcbffd0ffd6ffd9ffddffe3ffe7ffebffeeffeffff0fff3fff3fff3fff4fff4fff4fff5fff4fff3fff2ffefffebffe8ffe5ffe1ffdfffdbffd5ffd1ffccffc4ffbeffbaffb5ffb1ffafffaaffa6ffa3ff9fff99ff93ff8dff86ff7fff78ff72ff6dff65ff5eff58ff51ff49ff40ff37ff31ff2bff24ff1eff17ff0fff09ff03fffdfef7fef0fee9fee3feddfed7fed4fed0fecbfec8fec6fec2febffeb9feb4feb1feaefeaafea7fea3fe9ffe9efe9cfe9afe9cfe9bfe9bfe9cfe9cfe9efea0fe9ffea0fea4fea4fea5feaafeadfeb0feb5febafebffec7feccfed3fedbfee1fee7feedfef2fef9fe02ff08ff0fff18ff20ff2aff34ff3dff47ff51ff58ff60ff68ff71ff7bff85ff8fff9bffa7ffb1ffbcffc7ffd1ffddffe8fff3ffffff09000f00180023002b0034003c0044004d0056005f006900710078007f0085008b0094009a009f00a500ac00b300bc00c100c600cd00d200d600db00de00e000e500e700e900eb00eb00ec00ee00ee00ef00f100f100f300f500f500f300f200ee00ed00ec00ea00ea00e900e500e400e300e000df00db00d500d200d000cb00c500c100bb00b700b300ad00a800a4009e009a00960090008d00890082007c0076006e0069006600620061005e0058005600520049004400420040003e003d003a00390037003400340032002d002900260022002100220020001f00200021002400260027002c00300031003500380039003d004100430048004d0053005d0066006c0074007b007e0084008a008e0095009e00a500af00b800bd00c400cd00d600e300f000fb00070112011b01260130013801400146014d0159016601720181018e019801a301aa01af01b601bd01c101c901d501e001ee01fa01050212021c0223022c0234023b0244024c02500255025a025e0264026b027402820290029a02a602ad02ac02ad02ab02a802a802ab02ab02af02b302b702be02c502c902d102d402d102d102d102ce02ce02cd02cb02cc02ca02c502c602c902c902cc02cc02c702c302bc02b002a7029e0293028b0283027c027b02770270026b0264025b0255024c02400237022c02200217020b02fd01f101e601dc01d601cf01c601c101b701a9019c018b01750160014a0136012a011f0118011801160110010901fc00eb00dd00cc00bb00ad009f0095008f00870081007e0078007300730070006a0064005b00520049003d0032002a0021001b001b001a001d0025002a002d002e002c002a00290026002600290029002b002f00300035003b003f0045004e0054005a005d005e00610060005b00580059005c0063006b0071007a00830089009000950095009600960096009c00a100a400ab00b100b500b900bc00c000c600c900c900c900c500be00ba00b400ad00ab00ab00ac00b000b300b500b600b100aa00a700a2009c009b009a009a009e009e009900920087007d0077006f006b006e006c00670065005f00580050004100330027001a0011000e000900070007000200fcfffafff4ffefffecffe8ffe3ffdcffcfffc1ffb5ffa8ff9fff9eff9effa1ffa6ffa5ffa2ff9dff91ff81ff72ff62ff56ff4eff45ff41ff41ff3eff3bff38ff32ff2eff2dff2aff29ff2cff2cff2aff25ff18ff0cff01fff3fee9fee7fee8feebfef2fef6fef8fefafef6feeefee4fed5fec7febcfeb1feabfeacfeaffeb4febffec7fecefed3fed5fed9fedbfed4fecbfec0feaffea0fe99fe97fe9bfea7feb3fec1fecefed2fed2fecdfec1feb3fea7fe98fe8cfe87fe85fe87fe90fe98fea0feabfeb2feb8febbfeb5feaefea9fe9efe92fe89fe7cfe74fe70fe6bfe6cfe76fe7ffe88fe90fe8ffe89fe7efe68fe51fe3bfe23fe10fe06fe03fe08fe15fe1ffe29fe31fe31fe31fe2efe24fe18fe0afef2fdd8fdc2fdb1fdabfdb1fdbbfdc9fdd7fddbfddbfdd6fdc5fdb0fd99fd7efd6afd5efd57fd5afd64fd71fd82fd90fd95fd99fd9cfd96fd8ffd88fd7dfd76fd72fd70fd75fd7dfd83fd8bfd90fd92fd99fda0fda5fdadfdb6fdbbfdbffdbefdbbfdbcfdbefdc1fdccfddbfdecfd05fe1dfe34fe4bfe5ffe6cfe76fe79fe78fe77fe77fe7afe87fe99feb1fecefeebfe04ff1dff2fff3cff47ff4fff54ff57ff58ff5dff68ff76ff8affa8ffcaffecff0c00240035003f0040003e003d0040004b005f0078009900be00da00ec00f600f700f000e400d800d400d700e200f5000f0128013f0153015e016401650163015d0157015201520156015d016b017d018d019a01a201a1019a018e017f01700161015301480141013c013d013f013f0141014301430142013e0136012e0124011a0111010701fa00ec00dd00cf00c600c200c100c400c900cb00c700ba00a20082005b0033001200fdfff5ff0000170030004600550058004e0038001600efffc5ff9dff7fff6fff70ff86ffaaffd2fff8ff13001a000c00ecffc0ff90ff60ff35ff1bff14ff1cff35ff5dff87ffafffccffd7ffd1ffbeffa1ff83ff69ff57ff53ff5bff6cff88ffa8ffc3ffdaffecfff6fffdfffffffdfffdfffdfff8ffefffe4ffd6ffd0ffd3ffdefff7ff1a0042006f009b00be00d900e600e300d600c200aa009b0096009c00b600df000f0146017e01af01d501e601dc01c00194015f0134011b01170132016901b101050255029102b302b40297026b0236020402e701de01e7010502320265029a02c402de02e902e102c802a7027c024d0228020f0203020c0226024b0274029502a902af02a20282025c0232020b02f301e701e501ed01f601f901f501e901da01cd01c101b801b801b701ad01980172013c01ff00c3009500800083009c00c200ec000c0117010101cc0083003000e4ffb2ffa1ffb0ffd6ff03002b00450046002e000100c6ff87ff4dff1dfffcfeedfeedfef7fe06ff17ff24ff2aff28ff1dff08ffeafec3fe9bfe78fe63fe63fe7cfea4fed2fef9fe0fff0affebfeb8fe7dfe44fe15fef9fdf4fd04fe26fe54fe80fe9dfeaafea3fe8bfe68fe43fe23fe10fe0afe13fe28fe40fe55fe69fe77fe7ffe86fe8afe8afe89fe85fe82fe81fe80fe80fe83fe83fe80fe7ffe7ffe80fe87fe90fe9dfeadfebbfec4fec6fec1feb4fea4fe91fe80fe77fe73fe79fe94fec3fe02ff4bff90ffc4ffddffcfff99ff40ffd1fe62fe0afedafde1fd23fe94fe1bff9fff02002d001300b9ff34ff9dfe13feb3fd92fdb3fd0ffe96fe2cffb6ff1d0050004800070096ff09ff77fef5fd97fd6bfd73fdadfd11fe8bfe03ff62ff95ff91ff54ffecfe6dfef2fd93fd63fd6bfda2fdf4fd4bfe94febefec5feadfe82fe51fe27fe0cfe02fe07fe0efe0dfef6fdc8fd8efd59fd38fd3dfd6cfdbdfd1ffe7cfebdfed4feb8fe6cfefdfd81fd10fdc2fca6fcbdfc04fd71fdeefd6cfed9fe25ff44ff30ffe6fe71fedffd47fdc8fc7efc7bfcc9fc60fd23fef1fe9fff04000900acff01ff32fe6bfdd9fca2fcd1fc58fd1afef2feb1ff35006a004b00ebff66ffd8fe63fe1afe06fe2bfe7bfee3fe51ffb4fff9ff18001200ecffb3ff77ff45ff2fff39ff60ffa1fff0ff3b0076009700960078004000fcffbfff9cffa0ffd7ff3a00b80035018d01a501720101016c00dbff75ff56ff89ff0700b50070010d0267026a0213027801be0013009dff7affafff2d00d2007901fe0148024f021b02bf015301eb009a006e0069008a00cb001f017201b501d901d301a4015701fd00a9006d0056006d00ad0005016701c101ff011402fb01b2014901d8007c004f006000ad002901b5012d0277027d023502ab01fb004500b3ff69ff79ffe6ff990067012302a502d202af024f02cb014501d6008700610063008600c6001c017f01e9014c029502b802a6025402ca011a015f00c7ff79ff8fff1200ea00e801d7027f03b5037503d002f3011f01890050007e00fc009c0131029702bb02a6026b022102e901d001d501f4011b02330231020d02cc0184014e0141016f01d4015a02e9025d03970392035303eb027a021a02d901c001c701e401160255029c02ef0249039c03dc03f503d5037603e1022a027801f300c000f9009b018c02a203a5045c05a3057005cb04dd03dc02fd0170015201a3014d022803ff03a704ff04fb04a60418046c03c5024202f401e7011c0284020e03a10321048004b504c004ab0483044c041004ce0383033103e702b702b302e5023f03b0031704510451041c04c1035c030703cc02b102b402ce02ff0244039503ed033d047204840472043904e90391033a03ec02ab027702590259027602b402080355038803930372033603f302b6028c02790276028402a502d20208033a0354034b032103db028f0253022a0217020f020102e901c5019e0187018f01ba01020254029102a8028e024402dd0172011501da00c900dd0015016101b101fc01330245023202fa01a1013301bd004900e5ff9dff7fff9dfffeff98005301040278028a022a026401630065ffa7fe59fe87fe23ff09000101d1015002610200024401550064ffa1fe2efe1afe5dfeddfe7bff18009d00f90029012801f6009600100076ffe0fe6cfe33fe49feaefe52ff1600d00053017f014301a700c8ffd7fe07fe87fd75fdd4fd8cfe6fff4500dd001201dd00510097ffe8fe76fe63feb6fe57ff1600b6000301e100560089ffb3fe13fed1fdf8fd72fe12ffa6ff07001f00f5ffa5ff4cff09ffeffe04ff3dff8cffdfff23005100620055003000f8ffb8ff77ff33ffebfea0fe58fe1ffe06fe1efe6cfee3fe69ffdcff21002400e8ff7fff00ff89fe35fe18fe3cfea4fe47ff0c00ca004e016501ef00eeff8bfe18fdeffb59fb7bfb40fc6afda5fe9fff200019009effddfe10fe6dfd16fd19fd6afde8fd71fee5fe2bff40ff29ffeefe9efe42feddfd71fd03fd95fc33fcf0fbdefb0efc7dfc11fda8fd1afe46fe27fed0fd5ffdfbfcbffcb4fcd5fc10fd4bfd78fd8afd78fd4afd0dfdc7fc8dfc6bfc65fc80fcb3fceafc13fd14fddafc6cfce2fb5afb02fbf8fa3efbcbfb81fc36fdc9fd1dfe1ffed8fd54fdacfc06fc80fb27fb0dfb32fb8afb0ffcaefc48fdc6fd08fef0fd79fdacfca7fba4fadbf974f990f92bfa21fb44fc57fd21fe83fe6efee8fd17fd28fc4bfbb7fa8bfac7fa5ffb25fce0fc6bfdacfd9bfd4efddafc4dfcbefb38fbc1fa6efa4cfa5efaacfa28fbb6fb40fcaffceffc07fd03fdecfcd5fcc1fca8fc8afc63fc2cfcf1fbb9fb81fb51fb2afb0dfb08fb25fb62fbbcfb1dfc68fc8ffc88fc4cfcecfb77fbfdfa9bfa6bfa7efae3fa90fb61fc2cfdb7fdd3fd72fd9efc7cfb51fa60f9d9f8dbf85af92bfa1cfbf8fb93fce2fce6fcaafc46fcc9fb3cfbb3fa3bfadff9b0f9b6f9edf950fac8fa35fb84fba0fb7efb2afbb8fa3bfad2f98ef974f98bf9cff92efa9cfa08fb5afb8bfb94fb71fb2efbd7fa71fa11fac7f999f991f9a7f9c5f9ddf9e5f9d5f9c1f9bdf9d9f923fa8efafefa56fb79fb52fbeefa6dfaf6f9b9f9cdf928faaffa31fb7cfb7bfb2ffbacfa25fac7f9aff9eff97cfa2efbdafb53fc75fc44fcd4fb45fbc6fa73fa56fa73fabefa24fb98fb07fc5bfc8bfc94fc7bfc5afc45fc45fc5ffc85fc9ffca8fc9ffc91fc97fcbefc04fd5efdb0fde1fde4fdbafd6cfd13fdc0fc7efc58fc4dfc5afc86fccffc32fdacfd30feaffe26ff8effe8ff31005a004e0001006effa8fedffd47fd0ffd4ffdf6fdd8feb6ff51007e0031007bff89fe9cfdeefcb2fc01fdd0fdf9fe430072015502d302e202920201024a018b00e0ff59ff04ffe6fefafe38ff91ffebff3500610066004e002400f5ffd0ffbeffc0ffdaff0b004d00a10000015e01b8010402350244022b02e70189012b01e900da00fb002d014a012801b500080055ffd9fed4fe5cff5c009e01c80281039303f302cb017a0069ffeffe3eff4200b2012f035004cc049404c20392025b016100cfffb7ff04008f003701d0013f027e028a026a023802ff01ca01a5018c017a017d019b01dc015002e9028c0322048904a80487042b04a4030b036c02d3015e011c011e0178011c02e802b5034b047f045704e903670318031f037e032104cd04480580056b051f05cc048d0472048904bb04e9040505f204a9044704e2039c03a003ed0373041e05be053106780691068d068f069a06a906b906b106850649060906dc05e1050c0645067f069d06940680066a06620679069c06b306be06ad068306650660068906f906a10761082209a909cb098309ce08ce07c606e20548051e055805e105ae0692076708190979096c0900093f0858079c063c065c060b0715083409300ac00ac20a430a51091808e706f30571058e0534062d073d08090959093709b6080d08850732071b073f077807b207f60739088508ef086509d709390a600a300ab609f3080908330783060d06df05df05fe0541069206ec065b07c60723087d08c108ea080509f908bc085908ca072a07b2068006b4066407600868093b0a880a2b0a3909cc0724068f04390355022102ae02ff03fb053008190a410b450b2a0a5b086006d30427045c04350552063907a807a8075107e1069c06850690069f067606f3051e050404da02f3018101b10197020404b0054e077c080309db080e08d006710523041d038c026e02ba025c031c04cc044c0575053e05b904f30313034c02b40163016801a60108028102f6026803e3035d04d0042b0544050605730494039a02c6013f011f016101d101360267024102d0013c01a70037000600090037008800e2003e019801e1011a02480265027802840277024a02f7017301d00027008fff25fffcfe08ff39ff75ff9affa0ff8eff6fff5aff5eff6eff7fff86ff76ff61ff61ff88ffe2ff6300e10039014701f600540079ff87feaefd13fdcffceffc67fd12fec4fe4cff84ff66fffdfe62fec1fd39fde4fcdbfc27fdbffd94fe7aff3d00b400be005c00adffd4fef7fd38fd9bfc21fcccfb93fb79fb86fbbdfb22fcbdfc7dfd49fef8fe4eff1dff5afe1cfdb3fb92fa1afa83fac8fb88fd47ff8a00f300750046ffb7fd2afcecfa16fab1f9b2f9faf977fa19fbb7fb34fc7afc6ffc25fcc4fb6bfb41fb58fb95fbe1fb21fc39fc30fc1efc0efc1cfc56fca9fc04fd49fd40fdccfce9fb9dfa2af9e7f713f7ecf680f79af8fcf959fb5afcdafcd7fc5cfca9fb09fba5faa5fafcfa61fb94fb66fbbdfad8f916f9c2f818f911fa49fb59fcdefc8dfc76fbe3f927f8b5f6e5f5cbf577f6cff786f95afbf9fcfcfd32fe93fd37fc87fa00f9f6f7a9f714f8e4f8cbf97ffabffa94fa1bfa66f9aef81ef8c7f7d5f757f828f922fa02fb6dfb4bfbacfab7f9d5f863f87df82bf936fa2dfbc6fbd2fb3ffb56fa71f9c9f897f8d4f832f975f96df9f6f83ff894f729f73cf7d9f7c5f8cdf9affa1efb16fbabfaf6f93ef9bbf877f885f8daf846f9c0f93cfa99fad7faeffabdfa48faa2f9daf82ef8d0f7cbf729f8caf865f9cff9e3f986f9ebf853f8f6f727f8fff844fab1fbd8fc3efdcafc9efb00fa79f873f709f73bf7d4f77cf80af96df994f99ef9a3f99df9aaf9d6f90dfa59faabfad0fac0fa7bfafdf982f949f96ff918fa38fb84fcb6fd76fe6bfe87fde5fbbff993f7d2f5c3f4a4f475f5f1f6d6f8c6fa56fc55fda7fd4ffd9bfce5fb66fb62fbe0fb9efc62fde1fdd6fd44fd4bfc1efb18fa79f952f9a8f942fac3fafbfaccfa2ffa6af9c3f85af859f8c9f88ff9b1fa2efce2fda3ff26010402050227019affd4fd46fc37fbcffaf0fa58fbdbfb52fc9cfcbcfcaefc62fce8fb4efba9fa2ffa01fa22fa94fa41fb00fcccfcabfd9efea9ffaa005f018e010301beff1cfe8bfc76fb3bfbdbfbf8fc27fef7fe12ff7ffe7efd6bfcacfb7ffbeafbd4fcf8fd03ffc8ff2c002b00f2ffb1ff85ff83ffa4ffc8ffd1ffa6ff3fffb1fe0ffe71fdf6fcacfc9bfccdfc31fda7fd13fe4efe48fe14feccfd96fd94fdbbfdf7fd45fe99fefcfe93ff6a0060014802e202f20263024501ceff41fecdfca1fbe3fa9efaddfaaffbfffc96fe340085013f024402a00191006eff84fe0efe23fea9fe6eff3500c200f000bb0039009eff21ffe0fedcfef3feeffeaafe16fe4bfd95fc37fc5efc26fd72fef1ff5b01730201030503a602100284012e010e011e01450150012e01e90081000700a3ff6dff6dffa9ff2400ca007001f10137022702b8010f015100a4ff46ff5affe5ffd700f401e80274036c03d102e501f80048000b003a00a3001901690171014101f100a2009600f600cf011c03a4040906ff063e07b20699053e04f2021102b901d0014602f502b10373042805ab05e905bf050e05ee038c0226011a009aff9eff1100bf006c010d02b6028703a104f20549076308ef08cf081a08e8067c0537043e03ad02b2022b03da03a8046205db052b0657065c064a0609068105dc044004d003cf033f04e30494053106ac062707ba075e08f2082109b508c70786063f055904df039b036003fc026502e201b8011202f90223043205f10536061b06fd05110672062d07ff079308ca088808e5074e07100751071b081e09ed09390abc097e08d206fb04560354020c026f027503c504f905e9066b078307740755072e07240722070a07f906ea06ba066406d2050005260487036603f20300053e065c07fb070408af072c07c106ba061f07e8070609330a340bea0b160cac0bde0ac30991089c07ee06820659063506e2056305a404c503280307039003e804c006a008340a210b480bf10a5e0ac90966092309da0884080b086d07c4060a065005c50477047b04ef04b405a406a6077f080f0955093709c7084b08f007f8079c08b409f40a140cbe0cdd0ca70c430cd10b5c0bac0a9709200853067c04fc02f3017801920100029e026d03520446055b066207230885086708e7076707310787078508d109fa0ab30bb20bf50ad509aa08c507600767079507a007370749060b05dd0337036d0375041206c507f608660921094e08560799062506000614061c06fd05b3052105530474039a02fa01d6012702d102a8034d047e043c04a7030a03c4020103c803f6043a064f07100863085b082708eb07ca07d007dc07cd076f078e062f056803590156ffc1fde5fc13fd70febf008c03350601087f08a707cc05890384013700d2ff1b00a800190116018100aeff11ff11ff0600d001d2035505b3059004350258ffc1fc18fb9dfa30fb99fca3fe1801d3038a06b608d809a5092e08ea0584038e015100b6ff7fff6eff5aff46ff4bff6cffabff020049006f006b0014005fff75fe74fd9afc27fc0dfc19fc2dfc27fc0bfc26fcabfc92fdaffea1ff0200a6ff9dfe3afdf8fb3bfb49fb29fc91fd17ff4b00d300b0002f00afff8effebff7d00e800dd002e0005ffc7fdb9fc03fc9afb43fbe2fa7afa12fad1f9c5f9bbf988f91af968f8bcf77ef7ecf722f9f7faf0fc99fe94ffa0ffdafe8bfdebfb59fa2cf982f87cf815f9faf9e0fa7dfb7afbd4fac9f99ff8c6f7a0f731f859f9b8faaffbcafbecfa43f966f713f6c3f59bf658f860fa2efc55fda3fd43fd68fc4dfb5afab9f946f9f1f885f8aff79ef6bbf557f5b1f58bf618f7bbf63af5dbf29ef07aefbaef2cf117f391f458f5caf571f6eef779fa98fd900098020903bb01ecfe20fb3cf705f4e3f100f104f146f166f152f131f17bf15ef297f3d6f4a1f594f5ebf405f413f34ef2a3f1b5f084ef56ee8eedcbed70ef4cf2daf527f92cfb72fbfff95df7a0f49df299f199f132f2cff264f31bf411f57bf61ff853f9aff90cf991f7f2f5c4f410f4a6f3f3f24ef1caee04ecc1e9eae8dfe916eca9eea5f06bf127f181f03df0f2f085f245f47ef593f566f4a9f233f1b3f09af184f373f595f644f668f4e3f1b9ef97eeebee55f0cef1b0f2bff217f25ff122f16bf113f2c5f234f390f327f413f559f696f72af8d6f7a9f6f0f450f34bf20af28ff284f350f489f4def354f28ef040efe7eeb5ef0cf1c9f13cf14defadece3ea33ebd1edfdf127f6abf8d7f806f74af4fbf1dcf0e7f0bef1c3f297f385f4e5f5d3f73afa7cfcbdfd90fde6fb30f975f679f46df333f329f38bf256f108f04cefdfefe6f1abf441f7d0f8f0f8fbf7a8f694f528f558f5c2f524f655f645f61ff607f607f63cf6b3f658f7fef746f8e4f7d0f618f515f36bf178f05af02cf1b3f298f4c6f60ef91ffbd3fceffd36fec8fde0fcabfb61fa02f95af775f597f334f2f8f145f3e4f528f91dfceffd74fe14fe7bfd4ffdbffd7bfefefec8fea8fddafbb4f982f79af53af48cf3bcf3bbf423f65ff7d6f743f7ecf572f48af3aaf3b6f428f68df7b3f8c6f93cfb63fd1c00e40209051b063006b2052805e004b8044a04430385014bff11fd31fbd5f902f98cf84ef854f8a3f828f9e5f9d3fad8fbf8fc44fe96ffa4001e01b40041ff0efdb1facef8fef787f822fa45fc77fe65001702f0033406c1081a0b6b0c010cdd09a4064e03d20091ff2eff03ff99fef5fda3fd50fe3e001203f005eb0796081608eb0698055c042403c301470024ffdffebaff9101bf035b05e905790560043303820256028002fd02d7032305fa062109250ba50c6f0da70da50d8d0d3e0d640c970add07b30499010cff4bfd15fc37fbe2fa6efb48fdbc006805870a5b0f3313cf1562170618c317c81628150e13d910a80e510ca40980061f032e005dfe12fe38ff1e01f5023a04c70400057d0590066308f20af70d4e11c914d117e019911a8019001715148c11fa0f7f0f3d0f2f0ee50b5d0852040e0151ff2cff5200fe01990338052707d009720d97118615a7185e1a671a04196e160913910fb70c290b5c0b050d5a0f5f1111123811850fe50d630da00e0d117f13d6143114ba11c70eca0ce60c6c0f4913e61615194a191f18cd16e6153415e613c310820b5805070059fd37feb8010b069409550bcc0b8b0c9b0e2e12aa16801a7c1c9a1c651be0192d1982196a1a5e1ba21bc51adb18f01546127a0e050b7c0884072a082c0a360da210f413f4163a197c1aa81a9f19d61739165f15af152817eb181e1a631a8d1900186616d0142f1377113f0f9e0c400a8108e7071409b80b150f71128c1467140f12320e310ac307c107f4094f0df10f6410940e5d0b4008b20600076a08be09ee094e099509ad0c1e1418208e2e5b3c9046f54aea4879412636a628ad1a6c0d1e0229fa70f650f758fccc037d0b451128136f10e7092a0197f8adf2a4f081f283f743fea205360d93142f1b0c20a7214b1fa4193212450bf5068905fd051607af079807c3070309990b370fea12ea152d18d319071b001c8e1c751cec1b581bf91a981a7b19ed16a7123b0d6208f405b406420ae40ee0115d11440de806f10015fe38ff53032108f30a520acb062b02b1fee5fd7ffffa01a7034a03f500f7fdacfbddfa82fb9dfcfefc16fc38faa6f8f7f82ffc7002d20a8513c61a8a1f7c2113212a1f611c1c198e15bc11d60d470a6707730585046e04d3043505fd04d703e001a4ff12fefdfd81ffeb011b042505d604b303950208029f01760041fe72fb19f9b9f80ffb2bff35037505d604660134fc60f6abf0a1ebdee72de64de74ceb3af19df727fd4e018b04b407b60a2c0c560a5b0462fbf2f267ef80f3e2fe160efc1b77242a2672222d1ccb15df0f8709c401c5f87df0bceb68ec59f214fbb002e3056b032ffc95f23fe9d6e1ccdcd4d9a1d876d9badc6ce2eee9b4f197f71cfa0af935f564f0a4ec54ebc2ec26f010f40ef703f8b7f62cf4f1f18bf12cf4d5f93c01a2083d0ece106210b80da50905052000b8fa01f597ef5febc2e9aaeba6f069f7ecfdee013602d8fed3f8eff1b4ebcce679e37ce15be02ce020e1dae2e2e48fe609e727e691e445e350e311e508e846eb71ed85edb9ebefe865e6ece5c0e8bfeee4f620ffd0042b069302b0fa7ef017e6eadc20d64cd2b3d108d598dc9be792f40401500a4e0f0810410d5f08e5012df910ee57e1e9d43acc5fca19d0e0db02eaccf516fc2dfc70f7d2f021ebcde725e75fe84aea51ecf5eda2ee30ee3dec59e802e3f5dcbcd633d1daccb0c919c879c8e7ca76cf7ad5b5db89e1afe630ebccefa7f4cef846fb30fb86f80df5f6f293f330f735fcd7ff52002efd28f749f034ea37e545e109de4fdbe1d98cda50ddd1e1f1e659ebc3ee54f112f346f498f41cf3b2efd0ea21e5dcdfb7db5dd876d5bdd22fd097cea8ce4cd00ad3e7d522d830da02dd74e1ece730ef06f512f80ff81df6c4f4b4f58bf8bdfbe9fc58faeef421ef44ebbbeaa5ec60eee8edccea55e625e3f3e246e563e820ea5ce956e754e6fae7a6ec94f2d5f6bdf753f503f12ded36eb8aeaaae905e716e255dcffd7c3d62ed9e7dd7ce255e515e695e5bae5c0e76febd1ef7ff385f53cf65bf62bf69ef5edf34cf046eb6ae6b2e3ece435ead2f168f987feb9ff79fd38f983f4dcf0b6ee75ed85ec52eb9ce939e83ae823eaf2ed84f2d8f573f6e8f31fef52ea9ee7ede7f5ea34efd2f2eaf484f52df5bbf46ff4ebf3edf26af1a0ef1aeef6eccdeb27ea8de72ae433e10be0a2e157e647edaaf4effa04ff98004b00fafe54fdf2fb0afb99fab1fa2ffbb8fb01fcb8fbeefa64fad6fa9afc84ff7102d103e002bcff38fba1f6c9f295ef8fec50e9f0e545e340e22fe3bce52ae9e5ece8f08af50cfb2801d106df0af40c9e0d0d0e5d0f9a118a135113670fb207cefd4af493edf3ea06ec36ef9df2c8f451f5ccf436f4b0f419f79dfbce01b808dc0eb2124e139f109a0b0e06d401e9ff19004c012a02c4011a00ecfdf3fb65fa08f969f756f563f3a1f2faf3adf725fd61038809360f66140e19841c891dd51add13920951fefaf4e4efdcefaff30bf9cdfdc7004202860385054e081d0bb30c770c150bc7098e09a70a1c0c830c490bf408ce060806a7067b07f806220476ffb2fa7df797f6b2f7acf9a7fbacfd3900c70332087f0cd40f23120814a316cb1a112046253429bc2a6f298225111f5f16330ca0015df840f2f2efe3f0b7f38cf642f844f9c8fa2efe4204750c66158d1d8023b92694277526e4238320a51cc7188a15021303112e0fba0c9009b1065305bd069f0bc912e619b51e8d1f6d1c0c175c11d10c190ad708a2089609d80b710fd8139e179919a1194318c71635160b1607152b12540d4308eb052e08220fd0187221fa25d7257f22e41ef31d52208e244f282e294f26e620c71a97152212d40fd40ddc0bfd09dc081b09150a8e0aae092d073a045a0394067b0eb419e224762c572e562aa422b11af5148f122713c1149b153a15b313e7114311531202151f19dc1d4522ad253b278926ef23e41f461b151779135210b10d950b7f0a2f0b840df510ab144e17921899197e1b4a1f8225da2c27339d36ae35ea2f6326931a6a0e4004d2fd41fcd2ff1d07e80feb17011d7a1e3c1d6b1a55171e15d9138513a7147c17331cb622a829152f5931562f72297b216b194c1373105f10d0117913af13af111f0efc099d066d05cc06870a201088161a1dd4235e2a6c30d035b539393bbb3980347e2b9c1f2a1269051cfce6f72ff90bffef062d0e281321159514ac12de0f660ce60826069b05fe08a510361bf3254b2ddc2e902a2522b2183611da0c6e0b120c540d5f0e440fea0f271005108b0f500f6a106a133d18d71d0222012388206c1bbe15fe1143110a13b715091791157111cf0bbb062b049f047507540b3a0ec50ed20cda080604c1ff9afc9bfacef91dfafefb9200810895137420662c7d34d236d932d229521ec812df083c0179fb1af71ef4dcf22ff4c7f85100da090114ed1c66234127c128b9284328c72705276625f0210f1c1c14170ba50275fc26f960f820f9d1f92ef9e9f65ef377ef5becefeaf0ebd5ef70f631ff2609b712611a481f1b214520c41d711adb165a13f60fdd0c8a0a6209a409390b390d360ecb0cfc070400abf682ee09eadaeaaff06bf949022209280dd10e290fce0e2f0dfd089901edf756ee18e8c7e7a8ed9cf715026b097e0b79083f0282fbbdf636f502f77dfb5a010007210bc10c1c0b2b06eefef3f6f6ef95ebb4ea1aedaef104f7c9fb05ff390079ff38fd1dfa0af70cf5edf4eaf6a3fa15ff1203d0050407e206f6057d042f02a1fe8cf919f317ecc6e58de194e02de3cae83df0a1f708fd6dffd6fe2bfc0df9e3f62ff6b9f6d7f7edf8faf936fb98fcbafddafd72fcfef9b2f7dbf62ff8fbfa7cfd11fe00fc06f8f8f329f198ef5aee00ece9e766e3b9e08fe137e6f6eceef237f6adf6daf517f67ff8f8fb37fe01fda9f709f02ae97ae5cfe5cbe8eeebafed08ee1eee8cefabf209f6a8f714f67cf122eca6e877e84debd0eef6ef4eed60e73ce0bbda93d88ad96cdcbfdfc8e253e668eb24f280f922ffa9008ffd14f7b3ef55ea4be805e956ebd9edb3ef41f19bf2e7f24df10bed50e653dfe2dab1dae7de76e50eeb8aed92ec88e922e74de733ea05ef47f4b8f86dfca9ff130205032b0165fb64f21ee8e0debbd8d6d53fd4c3d1e8cc1cc65ac026bf9ac4ddd04ae1a8f1dbfe7f07e10bcd0d970e350e380c09088f011bfa31f392ed88e986e6aae303e10edf2bdeb3de2de085e14ae255e2bde133e1dee03fe05edf6cdebfdd77de34e147e5b5e933ed8eeef2ed60ecbaeacae976e9c3e834e706e521e344e3a5e6eeecacf475fbf1fe67fe88fadcf46aef27ebb2e78ce420e12fddb7d9bbd763d791d894da6cdcfbdd72dfd6e07de23ee491e5cee695e830eb04ef82f305f773f870f76df40bf19fee18edadeb00e910e4d8dd88d835d630d89cddc7e340e89fe934e85ae643e67be84decbfefc3f043ef94ec6cea89ea26edc7f002f4e0f509f648f555f40bf327f16aee13eb8fe85fe81feb67f03ff60ffa73fa52f7e6f1a7ec85e9f6e88aeae2ec5aee4beebbec1bea70e780e599e416e5bee6c0e886ea72eb18eb17ea7be9f9e9e9ebaeeebbf0def0d6ee61eb37e800e74fe88feb47ef04f254f3b2f322f4a9f572f8cafbd0fea700c30024ffd5fbe3f6d2f06deab7e4fde0ebdf17e192e338e623e87ee913eb7eedf6f011f5e1f8d1fbcdfdecfe3fff49fe21fb86f552ee76e7a4e3cde4b0ea23f3f5fa48ff24ffa2fbe6f6f8f283f0e3ee49ed49eb36e93ce801e9d8eaa5ec54ed76ec32eb78eb6bee02f4d9faa400c303fe033a021600defeeafe0900cc01c103df050a08a909f5092a08020421fe89f723f1aeeb35e779e3d8e010e0d3e1a0e6ecede3f584fc65005601b1007500fa014c05ff08010b200ac406cb02a100b20161056e094c0b9f091405fcffd5fc82fcc1fd35fe00fc19f7cef167effcf141f98a022e0ab20dfa0cec0927074c0600078a071c060d0249fcc2f65af3f9f236f5f6f80afd6f00aa029e031103f700e1fda6fa59f823f870fabefe0a041409d60cf00e7d0fd90e5a0dfb0a8d071a0307fe2df99ff52df40ef5b4f70ffb43fe0501a703fb069a0b2c119616651a5a1b3619c6144d0f070a9f0518025bff8cfd08fd4efe7201a2059809320cd10cbc0bed09420811074d06e7052a06be073c0b7510e41527192f184712b1087ffe21f7aef455f776fd490484095e0c3d0d430db60d380fc9112715cb182e1cdf1e1420271f2d1cb017aa124c0e0e0b8c082a067703d60093ffdb002505ef0b61137219361d8e1e0c1e9e1c6d1a11178112240d3d08a6054806c109b70ef6120a154415c3140b154d17d31ab11d611e101c7417df124e1060104712ba13a612d70eb609eb0504065a0a39111018321cac1cb81a0618ed15da14be137e11250e6f0ac4076b072409e20bc10e0711f21272159b18b91bc31d8d1d231bed176d15c9140a167117ff16c313ed0d5607bd02d90103052f0bfb1147171c1a821acd19cd19621ba11ec022f125e0264f259221f81c3319fb165816e6169517c0178517e816231681158f14e4129b10b80d9e0a2308c20602079109810ea8157c1e6327ac2e44335b344d328c2e162a8d255721f71c25188f13ee0f220eef0ec4117215f2180e1b651ba11a0c19e1169014e111e80ea30cb80b940c7d0f8913a317621b4b1e662039224b23dd22ca20041d6918c714061323137614661521157914b2145317371ddf24cc2bf62ff22f5b2cac27e123052202221d22b6206c1d9b18ae134910b50ea70e7e0ff10f870fab0e690d310cb50beb0b070d690f8812b8155118351937183e162b142913ef13b015701784185e1895174e17cc17f318481acd1a871a7b1a741b2d1e7722722628286926dd20f8184611b80b9109ef0a700ea912a51696199c1b491da91ecd1fa72094205a1f461d831aa5175e1598130a1265102c0e940b8109a7089d09510c7f0fda119d126811010fe00cd00b1c0cb60ddc0f1f12cf143718a51c3c223228522d8e30d430c22dd927d21fb516a70d3905d4fd12f87df4def3f8f67cfd2306f40e8a157b180718721582129110820f720e950c860901067303b102cf0346060809800bcc0df50fe2112213d512b1107a0d610aa808d908110ac90ad7090207830330013301b0038007ac0a000c6e0baa09fd074e0761078207f3062305500240ff9dfc0dfbf9fa4ffcdffe3c0298053b08b209f509970946095709c409060a910988086e07ce06fb0675071f072c057501b4fc73f811f621f668f8d7fb27ff7701440274015aff5efc08f907f6e2f3eaf238f399f4e9f628fa4bfe340359088c0c8a0e540d8708e300e2f710eff3e769e36be1bde1e1e309e7b6ea8aee1ff292f533f918fd510179059f080e0a820939074e04df015b00bcff48fffefdb6fbe1f82bf6a1f4aef4aef5c1f6c1f678f4c1ef3ce9e8e185db85d739d64fd7a5d9a8dbd9dcbedd3cdf7ce29be721ed5af106f3ecf1a9ef5cee19efd3f104f56af614f597f181ed12eb9aebb3ee3ff395f71efa9dfa6df9e6f6e9f307f120ee6deb02e983e646e4d6e28ce247e473e841ee85f48ff96dfb9bf9cff45aee52e82fe4f5e133e1eee0fedf61de9cdcffda20daffd9ead9bfd982d936d9b4d98cdb8adebce2b7e76dec79f06cf384f4e7f3e9f1b2ee4beba1e8d7e640e6a0e608e752e7a6e709e83be98deb32ee60f006f125ef41eb80e6e5e1b5de04dd92dba1d9bed6dfd280cf1cce0dcf6bd243d7b2dbd1de2be05fdf36dd90dab4d776d55cd42ad412d500d749d90ddc6cdf09e32ae7d7eb5ef083f4f1f7f1f993faf2f9e1f7d3f4e2f09eeb58e56ede30d707d13acd22cc12ce61d258d7eddb45df84e006e04bde71db60d8dfd5f9d31fd367d33bd4abd5f0d7f3daefde7fe355e794e9aae997e7e7e440e35ee38fe5d1e844eb09ecf1ea45e86be55be300e266e148e13ce1e8e1e7e311e72ceb2aef65f14af1f7eee8ea79e69ee24cdf88dc22dae0d757d6dcd518d6d2d685d7dbd7d2d899dbbbe03ce89df060f7f6facafa66f7c9f291ee30ebc1e8a1e6fae31ee1a1decadc2cdcdddc78de35e145e56aea6cf067f6fbfa7efdc4fd1bfc95f9cdf698f3c6effaea44e5dfdf0bdc73da39db34ddb1de05df4fde78dd28de17e1aee5f1ea78ef41f2adf37df431f526f6e9f695f6e0f4dcf116eeb4ea85e8e3e718e9b8ebf5ee35f2aef4def51af6e2f5ddf5bef653f8d4f997fad5f964f725f407f1cdee19ee9eee7fef0ff09befd7ed41eb82e864e6c9e502e7e6e913eeadf2ebf67efa47fd78ff70010f03f203ba03fd01f1fe8efbc6f850f757f7f9f7f9f786f660f34cefddeb5cea6eebeeeeadf328f852fbc3fc02fd4efdcafeff018106d60a460dc30c5109340457ff20fce2facefa6efabaf8a5f5ecf1bdeef6ec99ec3ced8cee6af02ef355f7ccfcf9020c091f0ea811a2131614fc1256102d0cec067401c4fcadf98cf82ff932fb44fe18026f06cb0a270e7d0f3f0e7e0a3705e0ff6dfb24f8a7f542f3def049ef83ef3df23df7f6fc8401b8037403ce014e00c0ff07006d0028003eff76fe8efed9ffea01c103ca043505aa05f6064609d30bb90d6e0e070e680d4f0d960d970d610c54091205ec0004fe10fdd5fd6fff6801d5032407ea0bea110b181d1d2420e7203020b31ea71cf6190516a810e50a17067703a903a70596072b08dd068d045e03c404f308050fc6143d180419b517d815371541164418241a5c1a3a186214b40f5c0b8208310724073b08c7096a0b330d9f0e6f0ff80f33107d108e113a1328153d17e918301ae81b4f1e5d21c0240527e92634241b1fd6182913d10edd0bf209f1075a05c602f4001b0157045d0a29125c1ae2206724d3246b226b1e9d1add17a31616174c1879195e1a721aa9198318ea16e214ae12f80fb90ca00937078306c808230eeb15d91eaf26c92be62d662db02b832a432aa82a2e2ba62aa628d5258322451fec1c521b801a091bb61c5a1ffb2292263b29c82a9c2aad28db258922801f111e6d1e59207423292659273927252657256e2654293e2d58310634b3342e34bc32e1306a2fe72d4e2c7d2b722b442c452e6730f3315d33ad3465366639d93c8c3fed401540383dc839523619335d30382d6529e8255b239d227a24f627d12b612fa331ad32b7331a3538377a3af33dd640fd4288433d42bf3f103ca73779337d2fb92b9c28d32576232b22c62129226d23ff24da26bc29d52d5a33203a91402f4531472d462c431140c53d973c173ca43a6137c132872d3c293a2723270a28122952293a29372af82c8831ed36cd3a4b3be137f43050282c209c1915157312cc10cd0fa20f23107a11b8133616b218271b281dbc1ef71f4c208b1fbc1d801a14161011bc0bdd066803a001b00161038e0526076c07ce05b2022eff2dfc92faaafaccfb34fd3dfe7efe65fea9fe9eff600180032205e505c705e804bf037d02f3002dff5afdb5fb94fad5f9c7f8d0f6c7f367f04aeef5ee13f3fdf9a501b207820a7d096a05c5ffabf9eff3fceeb8ea5de762e5d6e4c6e507e8ccea88edf8efaaf1a2f217f3f0f284f26cf2edf275f424f734facbfc0afe0efd04fae4f5c1f125ef1eef75f172f5bef95cfc28fcd5f889f29aeab2e2b6db6bd610d30ad139d0e0d0fad2d2d66cdcd3e22fe9e3ee49f38af602f964fa60fa8ef86ef491ee48e8cde256df36de6dded9de82ded0dc7ddad0d89dd885da43de79e20fe63ee878e82ae7f9e402e28ddeb6da54d6f7d163cee9cbe6ca24cbcacb8ccc75cd9bce90d050d3dbd555d7fdd695d463d1f4ce16ce2ecf59d1e9d25ed314d3ded256d4e6d71adc4edfd8dfc8dc8ad742d247ce7dcc3dccd4cbffca7dca70cba1cf54d79de05de961ef22f152ef23eb42e5aade99d7f5cff0c899c326c0bebe42befcbce5bac5b8c3b7a5b98fbebcc471ca00ceb2ce0ecedfcd27cf79d2edd6f8da2dde82e033e2f1e36fe5bae561e414e149dc76d7a7d38ad198d150d315d67bd977dc32de5fdec4dc41da8cd8c6d88adb5de04ce5b5e8e8e90be9a7e73ee7fae77de9beeaa3eab5e933e914ea51ed69f275f744fbf2fc2afc5cfae0f85ff8fff915fe2d048b0c9e16e7208e2a4432bb365738b93792357c333832c13189322e34033631385b3a323c6e3e4041bd4462497c4ef7526e5628583058db57d7577e580e5a745ba25b8c5a2958215597529650d74e114d8c4a69478c4498428242d144db48eb4df05253568a5790568d53e94fe14cb34aa949084931478e43d53de435012d4424361c011614120e10f30ff610c3110d1288113310280fa50e180e200d890a7e05d0fe47f7ddefebe904e517e040db9dd6ded299d1f0d2c3d5c4d8dbd9c8d759d3d6cdbcc854c537c34fc1fbbed2bb7db838b656b589b5efb531b50fb354b0f9ad48adb5ae54b13bb492b6d1b7bcb822ba00bc35bed7bfa0bf87bd19ba3fb6a8b330b3a0b4b6b76fbbb3be8cc1f5c305c68fc887cb63ce35d165d387d477d59ad632d820db08dff8e2ede64feaa0ecabee7ff0a7f19bf22df321f394f312f580f741fbb1ffa5031b07cc092d0b910bbd0a48083705ba02bf016b0347075a0b180e3a0e820bbb07ad040203dc02f1025f01d6fde4f869f31eefe0ec23ec73ec16ed09ed52ec1feb1ae993e6f8e34de14bdfa5de3bdf0de1bbe325e6b9e71ce8b7e6d1e3fbdf5adba9d69ed244cf02cdf8cb72cb15cb73cac1c833c66bc3cac04cbf7abfc1c0c9c2fcc465c62bc7bfc713c898c841c903c95cc7f5c37cbefbb7dfb117adc8aa08ababacf5ae36b1ffb268b561b9f0be23c6d6cd0bd427d8e4d911d9bad645d32dce07c880c14abb82b763b74eba68bfbac410c88bc934ca16cbe9cdb1d2b2d701dcd7dee5dfaee0f7e104e354e3aae1efdc70d6e9cf8ccacec77fc712c80ac90dcaefcae3cc7ed052d55adbeae1c9e78fec9cef1cf031ee0cea03e418dde1d5aece1dc85fc2a6bd4cbacbb74cb534b2d2ad83a8b1a37ca0d09fdea156a5e9a8f1ab40ae0fb11bb638bed9c97ad869e86cf865071814491ea6258529572a9828aa243c20871cfa19b519d61b761f85240b2a652e8e316c33ce331e34cb34ed3463344c32f32d38291e260226652a4132c83a5542bf47564b8e4f5855285c5a63ab686a6a9b695a67ff6466642565166641673b685869196c55702175f979617db47ecf7ee67d587cba7a72788e75157378719771f57332771d7af37bd17ba47af979017a077b857c857c8b7a0377fa71ce6c78681364445f9c59125276490a412b390733fe2ec22be228d4257021671c9217c012a60e550bb7074904d3016a002f01570423086c0b090dac0b08085003b9fde0f7c4f175ea4be23adabfd2e1cc2ec9e7c6abc56bc5bfc5ecc663c9a9cc5ed06ed45bd81ddc2de037e4ade753ea66eb8aeaace8a0e63be5d3e57ce846ecc6f0eef4a9f785f9e5faa8fb92fc93fdf2fd5efe4effc900f30307090b0fe215f01c39234029302fa0343d3a1940c345e64b8352f358685f6265086abe6d7c70f171b772c472e77103717e708570ae7159736f74a2748c737d71c96ffa6e1b6fe16f0a700c6f886d196cf96be86da270bb72f9720c70b76aee64be5f6b5c645b355b1e5bea5adc596c581b570e5522524f4ef048e942533d2638dd333330b42b2d26c51fa0187812710e4d0c110c8a0cb80b4909280578fff0f96ef5c8f163ef8bed13eb2de8bfe4a0e0c4dc62d93cd6ccd3c6d19acf6ccdd9ca7ec7adc36ebf23bbc0b7afb542b58fb6a2b89bbafdbb55bc17bc1fbcb6bc01bea2bfacc0cbc009c0a0be52bd7bbcf8bbf2bb32bc7dbc50bdbabe94c04ec3c6c6a2ca1ccfa0d335d7b7d9abdae5d9afd8e4d7bed7e8d8e2da77dcb4dd93def0deeedf20e22de55ee944eeaff266f6ecf886f9f0f8e2f7aff696f60ef86cfa9dfd01014c035e040f04d4016efea9fac2f6c2f32df250f1d0f01cf04aeea6ebe4e84ee69de4f3e356e35be2e4e0b3dea1dcb3dbeadb45dd4bdf9de0b2e093dff8dc68d988d50ad14fcc07c818c41dc1c4bf6fbfe0bffac0d4c17dc25fc3edc34ac497c4e9c36ac2a6c04fbe07bc52ba7bb8b1b628b541b394b1a2b0e1afc3af62b0f5b0eeb175b3ceb465b61cb8fbb862b952b9f7b7cab5f6b20daf1fab1da84ca693a6c9a898ab31ae8caffcae52ad4fab89a9c8a88aa8f8a7f5a61ba59fa270a0689e2e9cc7997d968d92768ff68dda8ed292c498819f9ba635ad6db360ba47c288cba7d6f3e2daefcdfc36082b115d175d1a551b051c261dbf1f0e249d28b12cd12fe8304230542ea02ac1257f20ee1a37164d13f4118312e1144718fb1cf922a4291831de384c40d747654faf56045e58647a68836a316afe67b965e6639e627362b3620d637e64fa66586adb6e68730877e679bf7bbe7c737d5a7dfd7b57794175a870e46ca26ab26a026d4470c073a276cf77a977b876d474b37286706e6d726986642b5e27571350bb48b2411c3b7334442ee7280524ea1f261c99173412dd0b7a0434fd9df682f051ebb1e6f9e1ddddbcda71d8aad741d84ad9c3da60dc8eddb7ded2df1ce06ddf7fddeed932d5dfcf49caf0c401c06ebb4db7b3b3b9b078aed5accfab70abd4ab56adfeaf71b330b781ba04bd07bf03c1a5c357c7b4cb35d05cd48cd7f4d904dcb3dd50dffce051e2b4e394e5a3e725ea21edd1ef64f245f530f891fbb2ffef034408c30cf2101b158119a51d6e21a824bf26e7278828f7281e2a872c24301935f23ace407046934be14f9b53c356fc58345a445a1c5938571c553c53fd514251bc501950fa4e6f4dbd4b094ad548704898485949784a2d4b5b4b074be849774822478b45bd439641673e7f3a83368d32312f8f2cb12919269f21371c9d164311340c1a08e304da0138ff04fd03fbe1f9abf9c7f951faddfaa0fad5f963f8f9f542f390f0d6ed92eb93e940e79fe475e19dddb7d927d637d365d182d036d051d04bd0fccfb5cf86cfc9cfd9d057d2eed33dd593d5ebd4acd3fad14cd0facec2cd9ccc7ccb28caf1c828c8dec778c810ca70cca5cf40d380d63ed92adb21dcf8dc13de4edfdfe031e237e203e1bbde80db7ad849d6bcd432d478d4d4d4a1d506d788d88eda19dd5fdf88e1a1e327e58ee61fe868e9bbea32ec25edb5edebed53ed5dec54ebece98ae83ae75de536e301e182de57dccfda69d946d856d714d6f2d459d406d437d4d4d439d599d51bd678d610d7ccd7dcd73bd7d7d566d3add02ace99cb66c9c8c774c61ac633c741c90dccdece6dd09bd0c1cf46ce78cd07cea1cf32d20ad51bd781d84cd941d905d9a8d8a9d76dd6f8d4dbd2a3d08dce6dccfeca92caeaca5dcc9acec5d001d340d538d78ed944dc93de45e0cee09cdf84dd64dbbed98bd9b0dafddbb5dcfadb50d9cdd597d278d073d054d213d572d8f8db35dfc4e284e687e99beb4dec3deb7fe909e820e743e7f5e705e823e726e514e2f8de8bdceeda80dafddaa8db2fdc1cdc14db6ed97dd7afd591d414d4ffd31ad4d7d317d302d279d0c3ce2dcd94cb49ca7cc9b6c8f4c710c780c5a1c30bc22dc150c24ec6fecc50d65ae176ecf8f64900e507980ea7149719c01dfa20f522d4244127362a642e37334237683a213cd73bbb3a583994379a36733641367e36d3366d3655361837c2389a3c4d42f947114d2351cc53fd5510580a5a9f5c4d5f7161bc6320668968b36b026fc5716c74937633783d7a477cb87daa7e477e597cc5798e76fa72c96f9b6c876938677065616456646b644664ed63c4622b61b15f065e905c865b375ae058885753557452ff4e664a6f45c4403e3c9e381236b933a831b22f082dfd29ab269e22661e201a48154110f40ac50434fe8af7cdf0f9ea77e60be302e1f1dfeedeeadd8fdc67daf9d78bd514d327d1e9cf04cf8ece51cecfcd18cd2bccd8ca67c926c81ec776c64dc675c6b5c6f7c609c7bbc63bc6ccc593c504c664c767c9e3cb87ce9bd00fd229d3f4d30ed502d796d9e8dceae0e9e4cfe884ec5def85f16ff32af594f767fb4b001c066c0c35125717f51bca1f312342268728522ae12b142d7f2e51300e32db33c2358937b939a33c0040cc439847b94a384d1f4f6e509751a0523f5375531a532d5229515150d14fc84fda4fc94f7e4fbe4ecd4d174d7f4c154cc64be54a2c498e46d442863e503a6a365b333c31692fb32dd72b39292326e4225f1f121c2f19471694131e117f0e170c160a3308e40661064d06e006d20727089107c4055f0217feb0f974f5f1f12cef9cec3eea12e809e685e490e3b4e2b8e15fe08fdec9dc85dbfada3adbeddba4dc2edd64dd54dd36dd04ddaadc41dcecdbe4db6bdca5dd74df77e14fe3d1e4d6e56ee6d8e61fe765e7efe7d0e825ea17ec63eeb1f0bcf212f48cf486f44ef44af404f599f6faf805fc27ffd401d603ed04280519052c0597058e06d5070e09280a190bf80b140d4e0e390fb20f9f0f060f650e070ec90d930d2f0d5a0c750b070b3f0b3c0c9a0d580edb0d1b0c54094706c40307021801c50088003700d9ff2cff37fe28fdf4fbfdfac8fa29fbccfb3cfc9bfb9df99df6f7f25def66ecdfe9afe7e6e54be41be3bde2d5e201e3ece202e259e07ddea9dc37db37da08d97dd7bdd5d4d376d23dd2dbd20cd478d56ed6ecd648d793d712d8bfd821d937d9fcd83dd86ed7d1d641d621d68dd622d7ffd7fad872d971d9f5d8b8d74ed634d565d45bd420d51ad64cd789d84fd9fcd9c9da71db50dc53ddd3ddf2dda6dd9bdc87dbd4da59dab5da06dca1dd99df95e1b0e22ae320e34ee28fe15ee14ce194e110e2f2e170e1c2e0acdfbcde3eded3dda7dd93ddfcdceedb6dda47d8f5d5e2d32cd222d196d018d08ecfb5ce69cdfacb69cac3c84bc7e6c5adc4fcc3c3c316c40bc534c674c706c9dfca45cd95d0a6d474d905dffce443ebbcf1d3f745fdc701e80400078508a009fa0ade0cf70e6a1107142416df171e1945199b184c172015da120e11ac0f3c0fde0f0311ca121e158f17751ad31d462118250f299f2c0a302c33be355238093bd63d3a410345cc48d94ce650bb54c058ab5c166011631365c865876546643562e35f4b5d8a5a0758ad558853a651a44f624dd04ad94706459e428040e43e753daa3bd63902380a365a3494321130252dc229e3258b22f31fc31d491c0d1b531945177d147610890b920589fe5ff76cf0d4e942e484df3edbcbd7e7d44bd238d025ce9bcbeec806c605c395c096bed0bc68bbedb939b8b7b657b523b43cb326b2b6b029af7ead25acb3ab33aca3adc6af01b2feb375b52cb652b6fbb563b522b541b5b2b5a0b697b75fb865b99fba3dbca5be36c16ec34dc575c646c7bbc8f1ca14ce48d2acd6e6da27df19e319e7beeb93f072f552fa7ffe2302de05ba09640e4d14bb1a42216a27322cab2f603258342c363a38f8393c3b003c0b3cee3b483c223d963e4c408c412e423a42ca417f41be4195420b44c8456e47f148324a514b8f4cb14d884ede4e284e784c3b4a9c4731456c43f041af40a83f623e0f3de53b613a6638d3351e32972db82889239c1e3f1a22169712b90f1e0d040b50096107700593038301cfff9cfe68fd57fc46fbbff92ef8caf65bf528f40cf383f1bfefcfed90eb6de986e7b2e52ae4e5e2b5e1bae0dbdfe8dee8ddb1dc3adbbad94ad827d792d683d6f4d6c7d798d837d988d970d923d9c7d85cd808d8bdd75dd71fd722d787d7a3d859da59dc7bde57e0c0e10ce366e4f1e5ece7f3e982eb82eccfeca0ecb0ec57edb3eeddf04ff37cf555f79ff850f9dff96ffa0cfb18fc92fd51ff68017d0320056e0666070e08d108a109050ae1091509a0073d069c05f0054b072c09a00a290ba30a1109fc06eb04f102210169ff84fd82fb99f9dff7a0f623f63ff6b4f625f7f8f6e7f515f4caf199efffed00ed8fec82ec86eca6ec0aed8aed19ee8bee6ceea9ed6decd0ea47e92de85fe7f0e6dae6b1e658e6c7e5aae429e3b4e17fe0f3df42e008e1ffe1dde23ce34ce351e33ce33de337e3a0e28ae133e0b2de90ddfedc81dcebdbf0da29d91cd762d53dd44bd494d560d77ad99ddb4ddddede81e0c4e1ace21fe3cae23be2fee121e21be3d2e484e601e8ffe811e9afe81fe845e7a1e649e6d0e57de55de51de516e557e570e579e559e5b1e4c5e3cde2d4e145e134e14ae15fe128e172e073df59de6dddf0dca5dc4cdca8db5bdaa1d8e7d630d5c1d3d2d219d2b7d1dfd15bd26fd368d525d8e1dbb2e034e661ecfbf26bf9c2ffe405550b2a102d14df16b3180d1a291b091df21f56230e27402ad52b152c2f2b352940279b25dc238922a321d920fb2035220924a3266f299f2b992d662f0531633384360f3a613eef422a477b4b8b4f2353f656d25a9e5e00639067ee6b58700d74a37687785379f378e077a07523720a6e6769df646a61fe5ea65d395dbf5ce05b885a6058ef5576538c50b24d1b4b5248e245f243e141fe3f183e603b52383035a7318c2e3b2c282aa6288c27f225f5238021101e201ace15ae10320b6b0503ffb3f8edf2aeed90e98de6f0e399e125df11dccfd8a3d598d249d0d1ced0cd46cde8cc47cc80cb92ca69c971c8d1c761c74dc7adc761c897c97ecbdbcd5bd0c2d29ad491d5edd5f9d5dbd508d6a2d64bd70fd8ded85fd9e1d99cda49db46dcc5dd5adf46e1a2e3d9e539e808ebeaed4bf14df532f9fffcb000e5036f07fd0b73112d18c31ffe26b22dab337638b83c98409a4323464348be496c4b9e4df74fa05211556856d5566a5647555854f3530c54ec542f566757b858cf597d5a0b5b1e5b8d5aab595558cc56ab55d2546254a75415557955d95592559e5453537a517e4fd94d2f4ca14a48497b4764455f432b41363fae3dd43b9139cc36fe32ba2e882a32263122a01ee01a4d172e142d119d0e410c2209330563009dfa06f57ff030ed86eb06eb91eae2e9a2e8afe6dce487e3a7e295e2f5e22fe34ce305e315e2dee074dfe7dda6dcb9db12dbc0da6fda03da8fd9e6d82ad881d79dd671d5fad3f9d1bacfafcdf7cbf4cabfca06cbc3cbe3cc2bcedbcf07d269d4f5d65ad933dbbcdc1cde4ddfa4e003e2f4e278e374e3cbe20ae294e187e14ae2cce3ade5ffe77beab0eccbee9ff0cdf198f2edf28af2fcf182f1e5f092f097f082f08ef0d9f026f1d7f104f344f4acf518f712f8e9f8caf976fa34fbf2fb1bfcbefbd8fa1df9eff696f4eaf152ef16ed13eba0e9d6e848e8fae7d2e767e7f3e696e6f6e528e51fe469e24ee034de23dca7da0edae9d928dab1daf6da03dbf8da84daded957d9dcd8d9d893d9aeda1bdc80dd15dee3dd0fdd76dbafd928d8afd694d5e1d41fd493d354d3f1d2afd28fd209d266d1bfd0aacf93ceb0cdb2cc19cc14cc34ccd5ccf3cde1cebfcf7dd09ad095d0c8d006d1c5d1f6d2ddd383d4bed43dd4c1d3b9d3f0d3b4d4a4d5e5d5a3d5ead4a2d3b1d272d280d20bd3c2d3f5d3fed30ed401d46ed470d596d603d878d96fda1fdb71db17db6eda9ad9a7d820d824d88dd868d93dda90da53da46d98ed7c4d51bd4e9d28dd2b4d240d34fd489d5fed6f4d818db5cddd9df45e2e3e429e815ece9f092f650fcd401be066f0a290d360f9010e4119d13b115a118651c59207c2462283e2b402d672e692ed32dc22cf32afc280627f2246d239122112256222a232024a7259f27ca29b22c2b30d9330d385e3c4c40134445478949494b5b4cda4ca14dda4ec450e653b657bc5beb5f7563f4659967fc672c67aa655c63a060fe5d3b5b6f58b6559a52534f374c16494e46f9438d41323ff43c803a4638633648340832672fef2b37289024de20ab1dd61acd17f0143d126f0f190d270bf308a106ee037f00fcfcacf973f6c6f371f1eeee7eec0eea6de70ee5d4e258e0b2dd9ddae0d6edd2e5ced5ca30c702c430c1f1be34bddfbb10bba6ba85bacbba77bb8ebc1ebe0cc020c20cc493c5a5c63cc782c7b8c7dbc704c85bc8d5c8b1c93bcb51cdfccf1cd317d6d2d84fdb32ddcfde7de0ffe1b1e3e9e53be8cfeabaed57f0bdf21bf5fbf6a8f87efa2efc1dfeb900ca03b0079e0cec117017f01cc8212c26712a7a2ead322437693b7a3f3443484604498b4bb54da54f17517f51c850d24eb84b454814458042d1409e3f533eba3ca53a54385836e1340f34df33df33ff335834b1341e359735ae35713500352734323346321231c92f852e022d7d2be729bf271925fc215f1e061b55180f1644147812f90f080dd8098c06bd03460196feabfb3bf83bf45ff0b6ec13e993e5aee119dd70d8f3d304d054cda6cba1ca5dca73cac1ca8ecb82cc69cd56cef2ce49cfa8cfe1cffbcf0dd0c8cf46cfb7cef1cd21cd5ecc70cb97caf0c948c9b8c813c806c7e4c5d9c407c4f6c37dc40bc59fc5edc5b9c5a3c5e4c558c63fc761c871c9dbcab0ccc4ce4fd1fed35dd6add8ecda1addb4df99e26fe568e851ebf6edb0f03ff32ef58af612f7adf601f658f5dbf404f595f529f6f6f6d9f7b9f80bfaadfb40fde5fe50002b01c9012a0221020702dd0170010501a4000f0064ffa8fed0fd3bfd39fdddfd44ff36013403f3043306c106bc0649065e0516048a02af00a3fe8efc74fa77f8a8f6e5f429f36cf18defaced01ec94ea8fe906e9bde890e862e8f7e76fe702e7b5e6cae672e784e805eaeeebecede1efbaf127f32ff4dff407f5bef40ff4c3f216f15eefc9edccec9eecf8ecb0ed6bee9bee3eee67ed10ecaaea71e936e813e7efe581e404e39fe13be023df5fde9cddfddc87dc08dcd0db0edca0dcbedd5edf22e10ee3f4e475e6bee7e5e8e6e91aeb88eceaed3fef46f0c1f0f5f0fcf0d1f0b0f069f0beefe2eee6edeeec4eecd6eb33eb3eeabde8efe670e580e459e4e2e474e5c5e5d0e587e56fe5dce56fe606e751e7c2e6ade58de49ee3b3e336e5ebe712ec78f164f7e3fdb704460bd8115218121e41239f27a92af22ccd2e54306d321e35c537893ade3c073e783e223ec93c433ba039ad374436583586347534df3446354736a237f338d33ae23cb33ee6401f430d456f47f1494e4c364f23529b54175709594d5aec5bfa5dc4602d657b6ae56f5175aa79747c367ea17edd7d8c7c377af3766e73796f7f6b316827656d623560d45d595bfa581156b352f84e4e4a28450e40df3a42367532be2e492b1b28c22406225920411f031f461ff61e351e0d1d111bdd189c16ba139a10560d9009f105b50259ff1efcecf846f5a5f150ee10eb39e8a9e5c7e29fdf25dc3ad867d4fed007ced0cb44ca04c900c8fbc6b5c556c4ebc276c135c04dbfc9bed2be6bbf77c0e0c195c399c50dc82fcb03cf3ed38ad762db48de60e0e7e1e6e2c0e389e4e5e410e550e599e57fe641e857eab4ec2def2ef10ff326f523f752f9cafb06fe5b0024033c061c0ae50ef21331196d1e182372279d2b512fd1321936cf384d3bbd3d07409e427a453a48ff4a8b4d8d4f5651d452de53b55427550b55c254385467539c528451e84fff4d984bd24821466943c9409b3ea83c153b233a75390739e838a1385a3854383c38433879384438c6372f3735365635de3463341e34fb33563360321c31122fa92c072ac62645238c1f2f1b9416e611090da808eb04770170fe70fbddf707f405f0e5eb4ce830e53de2a0df0edd5dda15d845d6e2d442d41bd41ed475d4ead45dd504d6a5d611d76ed796d796d7b3d7e3d72dd892d8c7d8b0d836d823d7a4d5e8d3ffd148d0e9cec6cd0acda5cc5bcc65ccb5cc04cd83cd12ce62cebbce29cf82cf21d003d1e4d115d397d43cd668d80ddbcfddd3e0dfe38fe629e9a4ebceed06f03ff23af44af656f813fac8fb48fd39feedfe61ff7dffcaff60000301e201a102a302fd01990060fef5fbbbf9b9f752f677f5b5f413f476f395f2b3f1f3f025f079ef01ef7cee18eefdedf6ed22ee89eecbeeeeee12ef08ef06ef41ef73efa0efdfefe9efe5ef0ef020f01ff004f05bef31eebfecdfeae4e818e73ce579e3fbe16fe003dfcddd60dcdbda65d9b7d72fd613d504d432d3b0d212d2add1cfd11dd2c9d2ccd374d4dcd437d539d556d5e7d570d607d7add7ced79cd74dd77ed672d55bd4ded26ad167d0a2cf81cf13d0b4d071d12fd268d281d2a5d260d209d29bd189d040cfe7cd18cc63cafac878c774c61fc6fdc57bc683c75bc854c986ca8ccbfdcc02cf13d15dd39fd525d739d8fad83ad98cd910da60da9dda7cda88d90ed825d6dbd3cfd11fd0b6cedccd56cde5ccbecc9fcc63cc49cc21cceccb0ccc60cce8cce3cd02cf37d0d7d1e2d396d655dad5dedee33de947eecdf2eef688fae8fd6901e60492088a0c77106f146e18071c541f4d228b2441267827e527e927ba273227c5267e26f5255f259a2454230c22f320f21f801f901fcf1f9320c22124230f2542275529742b642d162f1d3184335436e639e03dfb415c46964a764e1a5206550e576558d858a4584c58c6574657f4565b565755d3536851364e794a2646a741393db53865344b301b2c0d280524aa1f3e1bb616ec11780d89090c068403d5019200f3ffa9ff28ffacfefbfdb4fc49fbc7f9fef766f6f2f441f39ff1fbef1bee6cecfdea91e95ce829e79de5d2e39fe1d4dea4db0cd810d407d00acc37c8c1c48ec193bef0bba1b9dbb7ddb698b604b7edb7feb824ba5fbbb7bc5cbe4bc068c2a8c4d3c6edc82ccb94cd5fd0b3d34fd73edb84dfb7e3dee7edeb55ef2cf294f443f6bdf76af9fbfac2fccefe6f00c701e90255038503f1036a049205bc07610a9e0d5811e7149418931c8820b9241329ee2c693092333f360039133c353fa24234468549d44c0450c1522d550457fc576e586658f8579f574a57cf566456bb55ac547753e9510b50444e754cb44a37498947854543438240a33d373b2939b137cd36c23584342a336c31d02fb12ea82de82c5f2c6f2b662a6d291d28e026c7254224a6220021db1ea81c811af617741503133310600d850a3a07e8039f0018fdb8f968f6c1f200ef12ebd0e6b8e2e5de38dbeed7d7d4b0d1c3ce23ccecc986c8ebc7edc78dc88ac9bfca4ccc29ce46d0a3d200d521d7e5d826daecda54db75db83db9fdbd9db5ddc26dd26de72dfe2e051e2d0e330e54ae634e7b9e7b4e752e77de639e5eae3a6e28be10be12de1e9e174e385e5c7e73eeaa8ece6ee56f105f4f9f672fa28fec20148057a08430bf40d8510dd12211513178418a319621ab91ae51ad51a7f1a1a1aab193019c9185218951790163e15ae131912a110370fcb0d410c720a6408420622041b025400c3fe6cfd7cfcedfbbbfbf8fb5efcaefcebfcf4fcd8fcf1fc47fdd2fd95fe24ff21ff8dfe55fdb3fb3afa1ef97af863f870f856f810f873f796f6a8f57cf400f337f1f3ee67ecf0e99ee7a6e520e4b8e264e127e0cdde88dd8cdcaadbf6da80da00da8dd954d927d92dd983d9d6d918da4ada1bdab5d961d921d951d92ada6edb16ddfcdeb1e041e2aee3c1e4b3e583e6dce6ebe6b0e6f5e521e54fe449e369e2b2e1e2e06ce06fe09fe035e1efe131e227e2e2e15de144e1d4e1bfe202e43de5f1e557e6a4e6f9e6b9e7d6e8ffe91cebf5eb87ec1aedb3ed63ee2fefc5ef16f02cf0dcef59efc5eee7ede6ecdeeba0ea76e998e8e0e79ce7f7e7bde842eaa8eca6ef6ef3ecf79efc86016906b70a8f0ee4117714c7160f19381bc61dbb20b623fc265d2a532d1b307832ea33d0342135b634553434342d34c534b3355736e236f63633363535fb3372325831a8304430c930f93178338d35a13735399c3a893b043cda3c0e3eca3f9542f8458b49484d6b50ac5265546b551a560b57f857e358df59525a425ae759f0589557fc55b353ee50e34d5d4ad0467143da3f2f3c5938ea33452fa22ad4254a21fe1c7b180a14ae0f3a0b4e071c04600162ffd5fd1efc75facbf800f7c4f53cf51cf593f52cf62ff6aff582f47cf234f0d5ed48ebece8abe641e4f8e1cddfa4ddc4db12da4fd882d67bd418d290cfeecc4acad3c774c52dc317c13cbfd3bdffbca9bcbfbcf7bc10bd20bd4abdd5bd1fbf13c187c34bc6edc86dcb18cef9d069d49bd81addcbe192e6f2ea1fef51f325f7cafa40fedf00cc023004b704f7046c05da05b2063308e209010cb50e79117914ba17a01a491dd41f02224d240a27052a672d05314d344137da39f63bf93d094006421a442646f947c549824b1a4db94e30504b51175266522c5297519550384fa94db84b6f49ec460544f140ed3ddf3a00386335bd324330152e052c6c2a5229362811279b2553238f20891d3b1a36179314fa11b10fa00d6f0b7b09ab079f059b037d0114ffecfc0efb51f901f8bef616f54cf341f1f9ee09ed55eba4e915e82ee6b6e304e104dedadaefd711d52cd269cf8bcca6c9f7c653c4d4c1a0bf7cbd9fbb44ba53b90fb986b962baafbb46bdc9be5bc0edc134c360c463c507c6a8c66bc74ec8bcc9b3cbebcd7cd015d352d55cd719d968dab0dbefdc09de49df76e048e1fbe15be246e23fe24ce25ee2e7e2b6e37ae47ee58be668e785e8c0e9d3ea13ec51ed4dee7befdaf044f217f42ff631f852fa76fc6efe9700ea02200555074709940a630bc50bb50b940b730b200baa0aec09a808160765059803fe01b60086ff76fe79fd44fceefa95f913f895f646f5f0f3a9f28df15ef034ef4fee8eed1ded3fedb8ed84eea4efa3f061f1e9f1f1f19df13bf1b3f035f0f0ef9aef33efbdeed9ed9cec34eb78e9bce749e6f7e4e7e319e31ae2ece0a0df04de6bdc12dbc1d99bd89ed76ed631d518d4fbd221d2a9d14ad126d141d153d19ad135d2ddd2c1d3e3d4e3d5e8d6f0d7aad855d9fed955daa2daf2daf3daf8da1adb12db3fdbbbdb36dc03dd25de33df6de0bee1b4e294e35be4abe4dde4fbe4b7e464e406e454e39de2dbe1cae0c1dfd1dee0dd56dd46dd87dd42de44df44e053e14ae20ce3c2e352e4ade4efe4ede4a7e446e4b7e336e30ee331e3cce3e3e406e61fe725e8dbe898e9bbea32ec44eef8f0d3f3e9f646fa97fd1601c80423081c0b990d410f8c10ed116e1397157d189e1b041f782279254828dc2ad92c8e2eec2fa7304731e6315f3241336f3477359b368637c337bc3757377536c6354835d534eb34383557359e35c735b63506369e3677370b390e3b5a3d5340a0431547e34a754e81512c540f563d571d586d584d580b585b577356b055d054f1532053d4511150ee4d2b4b30484d454942693fab3c99395a36e432e32eba2a8c262722041e351a6916fa12df0fba0ce4094a077d04cb0123ff3cfca6f987f7a7f56bf4a0f3b6f2d7f1dff085ef33eee3ec43eb92e9a7e744e5d8e285e040de65dcd8da46d9bcd700d6e2d39bd130cfaacc51ca2ec844c6b8c482c399c200c2a5c17bc170c17ec1b1c101c280c248c337c45bc5c2c63ac8e7c9f4cb2acea7d07cd344d614d90edcf3de13e2b0e571e97dedd3f1e1f5c4f997fdef00090408077b099c0b980d220fa8107b125b14a31674195c1c7c1fc922c02582281d2b482d5e2f88318a33a335d037be399e3b6d3deb3e4c40864175426f438a44c2455a471949a64afa4bca4cfe4ceb4c8b4cf74b6d4baa4aa0497c48f9462e455e434e41233f1a3de73ab138a7366f3441325930672eab2c4b2bcf29622818278225e92360226d204f1e121c5b19a8163914c911b50fe70dd60bc009a507490535038501e3ff8efe53fdbcfb0efa46f837f648f474f277f089ee8aec3feaf4e7b2e568e362e19fdfffdda4dc76db4eda42d937d817d7f6d5cfd4a9d3b0d2ffd1b5d1e8d187d277d37fd461d50cd683d6ebd696d7b2d856da96dc3fdf1fe22de52fe800eba3edd6ef75f1a0f24df3a5f30ff493f43ef53ef651f758f882f9a0faadfbeffc3cfe87ff09018a02ec0359058e0672074a08fe088f09450af50a7d0b070c780cda0c7e0d610e720fba10fb110a130314ea14ca15c016b2177318ef181f19171905191219411972197e1925194118ea1636154c137611c70f380edf0c990b470a0a09ce0790067f057c046b0369024a01fcffb3fe4efdc4fb41fa99f8c9f618f56df3dff1aef0a7efc3ee2deeb1ed51ed35ed12edd3ec8cecf6eb29eb70eaace9fbe880e8e7e724e74be618e5a8e32ee277e0aede10dd7cdb2eda62d9e0d8b4d8dbd8ead8dbd8b2d827d866d798d68fd58bd4b4d3dcd247d216d20dd260d207d39cd345d4f6d465d5e9d596d626d7e0d7b4d848d9f7d9cdda91db9fdce3dde9deeadfd2e05ae1f6e1b3e24ae301e4b1e4fde42ae531e5e7e4ace48ae461e486e4efe46be51ae6cde64de7c1e712e839e860e86ae84de82de8fbe7d6e7e5e7fee71ee83de81be8d9e79de751e730e756e78ce705e8dce8dbe934ebe8ec9aee71f07cf289f4f5f6f1f941fd12014e0575098a0d6811a7148917371a991c231ff421b9249527582a982c972e48306b315232df32db32c132a5327632a532f032e532be32393239315c308e2fa72e092e622d902c2a2c202c682c632d942e9a2fb33089311b32f432e733f53488365d386d3afe3c9c3f09425d442f469a470b49684ad74b704db04e774fc04f3c4f294ebe4ccd4a9948384667436a40513dd8394c36a932a42e852a3b267821a01cc317be121c0eec09e805650241ff1ffc61f9f4f67df447f21df09ded30ebece8bee631e540e48ee33fe308e37fe2e0e119e10ae010df2fde48dd97dcf7db35db71da8fd97ed862d716d67ad499d268d01fce1bcc88ca8bc9fec883c8e8c70cc700c623c594c454c46ac48ac4a3c4fbc495c59bc63cc818ca06cc20ce2ed06bd232d541d89ddb54dff0e27de62deaa1edfef078f4b9f705fba7fe4102f105bf09250d481062132716d718941beb1d0a2029220d24fc250a28b229e52aa52bc02ba52bba2be62b452cc42c032d262d5b2da82d462e382f3b30453145322133f233ad343b35a435e53516365d36a436db36e5368c36f4355535c634883497349e3496346134ca3311332c32c530fa2eb52cd029b82691233d20081dd91968160713b00f2e0cc70850057f01aefdeef93af617f37cf02cee61ece0ea61e922e8e8e66be5e2e327e22be05fdec1dc43db18daf8d8b7d785d64bd51fd448d3a6d236d20ad2e6d1c7d1bcd197d16bd14cd119d1f4d0e3d0b5d085d050d0f2cfa7cf72cf2fcf10cf04cfe9ce0dcf74cffdcfe0d0ebd1d9d2e4d303d523d69dd748d9d1da52dc99dd88de99dfece077e284e4d9e617e96aebb1edc3eff9f13cf44bf65cf849fadafb61fdd5fe090049017c026503450405056505aa05c00573051605af041a04b503880362038303d50303042e043c04e2035a03b102bd01c700ebfffbfe36feb2fd2ffdcdfc8efc22fca5fb34fb9bfa01fa82f9cef8ecf7f7f6b2f550f414f3cdf18df069efffed5becb2ead7e801e771e5e5e376e252e135e04fdfd0de61de10dee1dd6dddd4dc42dc71db94dac5d9a1d858d70fd689d41dd3f3d1bdd0b3cfe0cef8cd49cdf8ccbdccd8cc49cdaecd44ce11cfc5cf9dd091d13fd2dcd26dd3b7d313d499d407d5a3d56ad614d7e7d7e4d8bfd9aeda9ddb35dcb9dc29dd4edd80ddc8ddf1dd4fdee2de63df0de0c1e023e181e1ebe14ee229e38ce425e60be8ede951eb6eec4fede8edb6eed2ef0bf198f24cf4d5f54ef78ef85bf9e9f931fa32fa38fa46fa54fa7ffaa2faabfab0fa98fa6efa41fae8f967f9c1f8d0f7c7f6c4f5c0f405f4a8f37bf3a6f30bf456f4b5f425f57ff525f623f73ef8b2f965fb0ffd06ff5c01db03cd06080a130d0c10d61230158417ea19301caf1e5921e723a9268c293a2ce72e54311b337f346a35b535de35e1359d35813568351535d53452343933ec314530552eda2cd02b272b3f2b982bd92b5a2cc62c142dcb2d992e5b2f75308e31a1322e34e135a237b5399f3b513d303ffe40e24237459247e449464c3a4ec94f1e51dc512b522d5283515850c54e764cb649af4622436c3fa23b6b371533b12efd2970253221f71c0c195f157811a80d060a4f06ee02f2ffedfc1bfa82f7cff468f27af0baee70eda6ecfcebaaebc2ebe7eb36eca8ecd6ece2ecf2ece1ecf9ec6aedfbedb3ee81ef06f02ff0f6ef2defe4ed46ec51ea26e800e6f4e31de2b3e0badf12dfb7de73defbdd5ddda1dcbfdb09dba5da6bda91da1ddbd8db0fdddfdefde09ee3a9e6a0e9c0ec13f04ef3e6f6f1fafffe5903e407160c4e1097148e18ac1cf020d724bb28892cd02f1033603662397d3c893ff34100449b457e463947df4732488248a2484548cf4747479d463846ea457545114595440944d943ec433444cf445445a545f2450246f6451446104603461f461046fb450f46e2458f453d458644a643d642b1417040373f973dd13b193a0338d735b5332331652e9a2b4e28ca242721f91c99183214700fb80a2a066d01e5fcb6f8a0f40cf103ee24ebaae883e662e49ce231e1dcdfcbded7ddb7dcaadbb4dac7d926d9b6d849d8f7d7a8d75ed755d78dd706d8c3d88ed94cdaedda4bdb75db70db2cdbceda59dac3d93ad9b6d828d8b7d751d7e6d6abd691d691d6e1d65dd7e6d79bd849d9dfd9a3da90dbb8dc63de69e09ee20ee569e78be9a7eba8ed95efbbf1fcf34af6daf87dfb19fedf009f033706d808500b7a0d880f4d11a712d013aa141c156b15851554152515f0149e1470144f140c14d21393132e13da12931221128f11ca10990f290eab0c140b8e093508cc0658050404b7028c01b600f1ff1dff50fe55fd35fc42fb57fa5df975f852f7e5f586f421f3c2f1a6f081ef2deee0ec69ebdbe989e83ae7e2e5ace44be3c0e13ce076de73dc69da28d8efd519d476d222d128d01bcf12ce39cd58cca8cb44cbc9ca57ca0fcabbc9b3c91eca96ca2bcbc9cb0dcc46ccabcc07cda0cd76ce1acfc3cf83d00bd19ed132d24dd229d2ddd13ad1cfd0d2d0f9d08ed17dd252d363d4b8d5f0d65dd8ecd91fdb48dc67dd13deb4de46df5adf5bdf5edf15df05df43df6cdfdfdf90e00fe1b4e174e2e8e26be3fce355e4dde496e534e6f8e6c6e75ae8fae89fe91aea9eea05eb1eeb1eebf9eab3ea84ea4beaf3e99fe930e9cbe8b6e8d6e833e9cae93eea90eae1ea0feb5bebfaebb1eca3edebee49f0f7f125f48ef654f976fc7dff6d024105a207cc09fb0b090e4c10ec129b157c18881b591e10219c23982533276d281a29ae29512ad42a7e2b162c332c132ca62bce2a0f2a60298728de2733275326b4253c25c524bf24f0242525b6255c26e326a62775284929972a362c022e253037320834d8357d370a39ba3a453c9a3dd53ec53f97407c413842c9421243ba42ed41c6402f3f703d813b14395c364b33b72f012c2528eb23a01f331b7616d511520dc10884048b009bfc0af9c2f579f27defb6ece9e96fe734e5ece2d5e0cedeaddcdeda79d965d8e3d7b9d793d798d7b6d7dfd75cd808d99ed922da5dda3fda0fdac6d95ed9e5d827d81ed7f7d5bcd491d382d265d12dd0d4ce5dcd00cccfcac8c9fcc847c8aac753c730c751c7d2c769c823c934ca70cb11cd47cfb3d166d47ad78bdacfdd79e118e5d7e8d5eca1f079f492f874fc4e004404e307740b3e0fde128816611af61d7e212f25a528f42b1b2f99318f3343359f36f1375c397c3a3b3b993b783b223bd93a8b3a393acc3923396238af371937a9362f368635b734ca33fa3278321e32db3195310f316e30dc2f352f912ee72de82cc02b912a3229d7278026d6240d2346215b1fa01d201c751acb181c172715471382117a0f5f0d130b4d087805a902b0ffe1fc23fa2cf75bf4abf1f0ee81ec3aeadee7bee5cce3ede16ee01edfc5dd92dc60db23da17d90fd8ebd6c7d588d44fd369d2ced180d173d161d14dd150d16bd1cbd164d204d3aed348d4d3d493d583d67ed78ad86ed917dacdda92db67dc70dd69de2fdffedfcde0b3e1efe23fe46de596e690e771e89be9f8ea73ec34eefbefb6f1b3f3d0f5eff73efa78fc7cfea000cc02ed043a076409260bb80cfc0de90eda0fb4104711d2113a126512a212de12e812f112ed12c012b212c912cf12d812d512971250122412f011b3116111aa108c0f390eae0c0f0b9a092808a8064a05e80379023601eaff72fefffc6bfbb1f923f8a4f621f5caf366f2ddf06eeff5ed70ec21ebd9e98fe877e75ae633e531e41ce3fde109e10fe028df7eded7dd48ddf7dcaddc8bdcaedcd0dcfddc3add39dd1addf7dca0dc40dce9db5ddbc3da2eda77d9d5d862d8f1d7aed7a9d7b4d701d896d834d9ecd9a9da20db7adbbfdbc5dbc9dbcfdba9db98dbafdbccdb3bdcfddccbdddade1ee055e1c9e26ee4f0e581e705e92dea49eb5dec27edf2edb1ee16ef73efd2effdef49f0b1f0f6f05ef1edf177f239f320f4dcf481f5f1f502f6eaf5b5f560f51df5f0f4daf4f5f429f55af56ff532f5a1f4d7f3e1f202f25bf1cff072f033f0e6efb9efbaefc8ef1df0c2f094f1e2f2c3f402f7c2f9dafcdaffd702c9057208120bad0df00f12122214fd1510187e1a001db81f6d22aa24a1264f288629b12ad22bb02cb02dc82ec02f01315d327733953466358e357535e534b8339232663129307a2f0f2f972e752e432ed42dc12dd62df72daa2e9d2fb2307d32bb344f37863ace3dce40c7435e469b48ee4a074dd94ea1500f5241538d54a4557d561c57fa562656e054ff52e050ca4e714c0f4abe4715454242413f923b783726336e2ede29b7259421a91dea19da15cf11f00dda09d805f601cbfdd0f957f631f3cbf02defcaedc9ec30ecafeb9deb03ec68ecd5ec2eed1dedfdec01ed08ed49edacedd5edd3ed9ced06ed3fec50eb25eaebe8bbe790e683e590e49be3a0e2a8e1afe0aedfa2de70ddf2db49da9fd806d7c9d5fdd462d40fd406d420d4b1d4dcd553d73ad982dbd6dd98e001e4cfe73fec2df1f4f5b1fa61ffaa03ed07460c4f1055147118531c562085246528142c822f5432e8346937a139d23bf33db03f364188426643fc433a44f5437843e4424342dc4191412541a440e43fe13eea3df43c023c3c3b6a3a8e39e2383e38ae375e37ff369b3669362a36fa35fb35c2355835e53423345733c43210325731a6308b2f402ef82c622bc6293e285f266d2481224020f81daf1bfa1821162e13d20f710c16096c05c5011ffe3bfa86f614f3bbefd6ec59ea03e810e667e4cce279e15ae04cdf8ade0adeb1dda7ddd3dd19de97de3adff1dfc4e091e143e2e0e269e3f4e393e436e5cde52ee635e6f3e579e5eae480e43ce415e418e435e46ae4e1e488e53ee600e797e7e7e720e84ce875e8cee839e98ee9f1e955eab8ea63eb4fec56ed9beef8ef40f1b3f24cf4ecf5d6f7f1f901fc37fe6e00660256042806a7071809720a830b8c0c8a0d470e050fba0f1b1042100f10330fe10d420c480a490875069704c8021c0153ff89fdecfb3bfa81f8e2f61af53df395f1f5ef6fee3eed0aecbaea78e9eee723e671e4ade2fee0cedfdbde2fde08defcdd08de64deacdee4de3bdf3edff4de9bdee1dd0bdd70dcbbdb0cdb79da7cd934d8d7d619d555d3cdd126d099ce45cdcacb74ca6cc952c862c7a8c6c1c5fec48ac41ec408c44dc476c4b6c412c53bc58cc51ec695c62dc7d9c736c89bc824c995c95dca89cbb7cc28cebbcfefd00ed216d3bad381d485d56ed6a7d71cd956dac5db5eddaede11e056e1ece142e263e214e202e237e23de26be292e249e218e214e2f8e130e295e2b9e2fae253e396e330e40fe5dfe5d4e6c6e781e853e931eaf7ead0eb96ec23eda2ed02ee3eee80eea8eeadeea5ee72ee1ceec5ed5bedf4ecafec6bec33ec06eca5eb16eb6dea9de9f8e8cce81be919eac6ebceed2cf0d0f26ff528f8f5fa84fdf2ff4302510484061509e60b360fe1126416cb19e21c501f6c213c239124e9254c278f28302a142ce32de82fc93112331634963461340f349133d232603200326b31ff305e30492f352ef02c762b622a9e293629a829b42a392c702ee8306833133680389c3aa63c6b3e0e40e341b5438e45844733499a4acb4b804cdc4cf84c8f4ccb4bcb4a5b49c44722462744f6417e3f5f3cd538f7348b30ec2b352727221f1d3e1847139d0e480ae905c101bffd85f96ef593f1c3ed77eac3e75ae57ce304e288e045df30de10dd3ddcaedb29dbf4da02db29dba8db5ddc02dda6dd11de1ede04dec9dd74dd2dddd9dc66dce1db3edb93daf3d95ad9cad82ad865d784d670d53bd414d3ead1e8d041d0cbcfa5cfeccf55d002d110d236d3a5d480d670d8abda50ddfedff1e23fe67de9dfec7ef0f3f389f769fb35ff35038207a80be00f371445184c1c692042241028de2b3c2f4a3208352337da38593a763b763c6c3d163e973ef73e0e3f1c3f393f463f663f843f7a3f6c3f513f1a3fe33e7a3ec13dd73caf3b783a8939c7383538d4373c377336ad35c234f1336a33c832143259313130db2e8c2df42b5a2ae02820275e25b523c021ca1fed1dc81bab199e173315b2122410420d7f0afa0767050d03d10056fef8fbccf9adf7ecf560f49ef2c1f0b2ee61ec3fea65e8b8e656e506e493e225e1bedf6bde61dd96dcfadb9bdb64db4edb5fdb80dba7dbccdbe6db00dc1edc40dc74dcb1dcf0dc44dda2dd00de70dedade3bdfb5df41e0dee0abe182e249e317e4d4e47ce543e611e7d0e79fe863e918ea0eeb4aecc8edb4efd7f1f3f323f646f846fa65fc89fe830077023e04b1051607620878098d0a820b2b0cc10c430d980d000e740ec30e110f490f360ff70e8d0ed70d040d320c430b580a800987087e0786067b0572048e03960289018f0081ff6dfe8cfd9ffc91fb82fa30f9a1f724f699f40df3bef16cf013eff1edd3ecc7eb0deb64eacce971e909e995e83ee8b7e70ae763e685e592e4b9e3bae2ade1aee079df33de05ddb7db7bda77d978d8b7d75ad727d73dd791d7bdd7c9d7b8d75cd7fcd6c5d68ad671d674d64ad61dd606d6d9d5c6d5cbd59fd567d533d5e4d4c6d4edd41ed57cd5fad55dd6e7d6a6d766d85fd97fda82dbabdcfcdd3cdfa7e01ee246e358e449e5ece5a7e681e744e843e96cea7cebb4ecf0edd9eea7ef48f09af006f1a0f14bf241f35bf44ef53af6fbf66cf7b4f7bff77af715f794f60af6a9f563f532f515f5d8f479f4fef349f382f2bcf1e2f028f09aef12efc0eea3ee86eea5ee01ef63ef09f0f2f0e7f13cf314f549f730fabbfd700154052a09800c9e0f9d1250151718f81aa11d65204b23192628295a2c2f2fc531dc3326352636fb36993782388b39593a3b3be93b1b3c3c3c003c1b3bfb396838583692341133db317d3188319831f2311a32df31d831d531e03190329733dc34c536e838223bbb3d3d407d42b7448b460b489e49154b974c604e005064518c520353e35257522051884fc04d814b1b49ad46eb432441643e3c3be6374f3405305e2b76261621cc1bc716c411260de908a104a300edfc28f9aef578f228ef12ec3be96ae610e43fe2b6e0b8df24dfa9de84dea5ded9de61df18e0bce078e12ae2b0e246e3cde322e460e453e4e2e334e339e2fee0b5df53dee4dc80db15daa2d82cd7a4d51cd49ad227d1dacf9fce74cd68cc64cb8dca17cae8c91fcacbcaa3cbc1cc4fce21d077d27ad5ced883dc9de0aae4d0e832ed72f1c1f542fa93feec027e07f10b78103215b519241e9822b4269d2a652ead318b340c37e8384c3a5b3bf03b413c693c3f3cea3b6d3ba53abc39bd38a1379c36ab35be34f9333e338432f5317231f7309e303430bd2f672f152fed2e1e2f6c2fde2f803002317d310d326e32c03211331233ef32c2324832c031363157305a2f442ec12c122b3629dd265524a8219a1e851b6218da142b113f0dd8085f04e7ff4efbf5f6d0f2a4eec0ea14e77be341e054dd8dda2ed822d650d4f8d2fdd148d100d1fbd026d19dd130d2d8d2b4d3a2d4b3d500d753d8aed90edb3ddc5cdd89dea0dfbbe0c8e179e2dce2f6e2ade24ce2eae15ee1cde02ce04ddf6cde92dd99dcb2dbc2da92d95fd82dd7f6d518d596d457d49ad443d528d683d72cd9efdafedc22df24e14ae370e57ae7c6e942eccbeeadf1b0f48df77afa47fdc5ff5602ec045807df09510c5a0e3110bb11b7126513ac133d135212fb101a0f180d260b1d09330774059d03da014800adfe1cfd9ffbe7f90bf838f651f484f200f18bef2aeef5ecb6eb81ea83e98ce8b5e728e7bce699e6ede67ce744e83fe90ceaabea32eb65eb72eb7deb47ebfceac2ea5beafce9bfe94be9bae817e80ce7d4e5a2e439e3dde1b5e06bdf2dde1adddcdba7da9cd965d833d728d6f5d4d9d3fcd210d24dd1cdd03dd0cecf9ccf5bcf43cf6dcf8ccfe0cf7ed018d1eed106d306d425d55cd655d755d85cd91fdaf6daeadbb4dca7ddbcde8bdf55e005e141e16ce194e178e17ce19ce184e184e19be17fe187e1b4e1bce1ebe13ee279e2e1e273e3f2e395e450e5ece599e643e7bce725e867e871e872e861e842e83fe83ce83ee85ee870e87fe89ce895e88ae8a2e8b6e8fbe889e915eab7ea78eb0decb3ec98ed85eec0ef6cf13ff37df541f830fb74fefc0148057308830b290ec0107113fb15ad18901b4c1e28211b24c1264829882b1e2d612e572fe52f9330623116320433f73399344135ac358e354435983468334c3239312230872f1f2fa42e6f2e2f2ebe2d902d6d2d3f2d7f2dfc2dae2e0630b2318033a335af378439723b3d3dec3ec4407342f3437c45c846ee471e49014a9c4afd4acb4a2d4a4849d74715461d44a341f13e203cea3897352a32452e302af5254f21ac1c26187b130f0feb0ab806cd0221ff53fbb3f73af49cf044ed45ea64e7ffe416e35fe124e062dfd2deabdecaded5deebdefbdedadecedee7de07df54dfbcdf17e079e0d8e019e141e142e106e19ae00de06ddfc6de25de83ddcbdc05dc38db56da77d9add8ded72bd7b0d64fd637d680d6f1d6add7c8d8ffd983db6bdd6ddfbae166e41ce713ea63edaaf01df4ccf754fbf3fec5026706170ae80d7411fd14a518121c901f3723a626172a962dc030c433a236f638eb3a8b3c983d663e153f793fd23f19401640fc3fc43f5a3ffa3e963e103e973d0c3d673ce73b6c3bf73aaa3a423ab93933396e3881379e3685355c345e334e326031c1301630812f192f7c2edd2d5b2d9a2cd32b232b2f2a3d296f2865275c265725e8235222a420881e531c141a7217c1140f12190f3e0c82099406b703dc00b8fda2faa6f793f4c3f133efa5ec60ea53e843e66ce4b7e2efe04edfd0dd5adc36db65daccd995d9a3d9c4d905da3bda43da30daf9d9a1d957d926d91cd94dd9abd930dad6da80db31dce2dc7fdd1ddebfde63df2be00fe1f8e1f7e2e6e3a4e451e5d7e52ce686e6dae624e7a7e756e824e942ea83ebb9ec0fee5bef81f0c2f103f323f466f5b4f6f7f778f91efbb5fc6bfe10006d01c5020e042205400656072b08fd08c909630a030b9d0be00bed0bc30b2d0b670a92098108620753062205f9030003f901f6000700e1fe94fd4afcd9fa64f924f8e8f6baf5bff4b8f3a8f2b2f19cf072ef64ee45ed2eec59eb9dea0fead4e9afe9a6e9cae9d0e9bce9a7e94fe9d5e868e8dae756e700e791e620e6c4e52de582e4e4e308e31ce240e12ee020df41de4add6adcbadbe0da0ada5bd985d8bdd722d75fd6afd538d5b6d471d483d49bd4e9d467d5b5d503d653d655d64ed64dd618d607d62cd64bd6b4d65fd7fcd7d1d8c7d988da5edb31dcb5dc47dddedd43dedcdea3df59e053e173e267e373e477e52ee6f2e6bfe76ae84be94dea34eb39ec34ede7ed88eef3ee01efeaeea5ee31eed6ed8aed52ed54ed5ded5eed69ed49ed0eeddaec87ec43ec37ec33ec72ec13edcfedd3ee20f04ff18ff2edf31cf580f646f82bfa8dfc77ff7d02e1059809220dbb10511470176a1a531de81fa32299257328822b9f2e4c31c633e035443760382f398c39013a7c3ac33a443bc43bfa3b493c673c133cc13b343b523ab2392339893860384538ff37f537ca3757371637bb3639361f3637368f36a9372d39f43a393d733f71416f430f455e46ba47e8480e4a724bb74cde4df64e884fa44f684f844e414dcd4be349db47d1456e430141823e803b4038b93484300f2c682741221c1d0d18c712ca0d200969040e0006fce4f709f474f0cdec80e999e6c9e373e194dfd5dd7bdc79db80dad1d96dd91ed923d971d9ccd955daf4da74dbf7db74dcd0dc27dd6cdd8add96dd8cdd6cdd4fdd31dd14ddfbdcdddcc0dc9fdc77dc4adcffdb91db0edb65dab1d916d985d81dd8fdd7ffd747d8f3d8c9d9e9da6fdc18de0de073e2fde4d2e706eb34ee80f102f555f8a5fb14ff44027205d008110c720f1a13a216311ae01d5421bb243328602b5e2e39319f33b835a2372a39803ab93ba53c6a3d0f3e693e993e963e443ec33d0d3d203c243b053ac2387a370d368d342433b3315a30372f0e2ef42cfa2bd92ab229a428762760268525a224e22350239422d9212a213f20561f851e841d961cc31bbf1ac219c618761713169214b512d010e00ea50c6e0a2a08990511038500bcfd0bfb52f859f579f2a7efc2ec2beac8e763e536e311e1c6de9edc80da57d86bd69fd4e9d28cd16fd090cf1dcfe0cec8cee5cefcce0dcf2dcf27cf15cf18cf0acf21cf78cfe0cf81d056d11cd201d3ffd3d8d4c2d5b9d687d77ad893d99ddad5db11ddfbddc9de65dfa9df00e066e0aee020e196e1d4e12fe299e2eae27be32fe4cce4a1e591e669e779e8a0e9a0eabfebdfeccbedd1eed7efa9f098f199f284f3b4f41ef686f721f9c8fa2dfc81fdb0fe7eff2c00bc00fe003c0183019501a2019b0132019600dbffd4fec8fdd2fcb3fb8ffa73f916f89bf61cf55bf383f1c5effaed5bec18ebf6e903e94de883e7b8e60de649e589e4f6e35ce3e3e2bae2abe2d2e241e3a0e300e47ce4cfe41ee586e5b5e5c8e5dfe5b7e58ce58fe56be540e51be597e4e2e32de330e22be147e02cdf12de25dd19dc32db91dad0d91dd985d8a6d7c4d6fdd503d524d474d3a0d2fdd199d125d1f7d011d11cd166d1ead14ad2d7d283d3f9d39ad46cd52ed644d7a5d8f5d973dbf9dc30de68df9ce09be1c8e21ee46be5f3e68fe8f6e94beb5aece9ec30ed1fedb7ec4cecd6eb59eb0aebb9ea58eaffe974e9b8e8f0e7eee6dbe5eee404e45ae328e338e3bee3c6e4f0e54fe7dee83feab8eb7aed55efb7f1c9f432f827fc9200e3043f09930d72113515fa187c1c27200b24c527a02b7d2fe032fe35ac38813ad73baf3ce53c0b3d2b3d173d363d4e3d053db13c083ccc3a7539d537de353834ca328b310c31f230f7307531f5313932bb322c337a333d343935603632384e3a803c143f9141c7430346e7476c49f24a3d4c6c4ddf4e4b50b15128532b54aa54b954fd53b7522b511f4fe94cbc4a3e48ad450f43eb3f743cb4384d34ab2ffe2a01262021791caa171013be0e520a290652026cfed4fa9ff776f4b2f15def1aed31ebb4e959e86ee700e7b8e6bde602e735e78ae70be87ee80ee9b3e930eaaaea29eb8aebf0eb4aec66ec4aeceeeb42eb6aea71e949e801e797e50fe489e21be1cfdfa4de8cdd75dc53db34da2bd940d894d73cd72ed78bd75dd873d9d3da68dcefdd8edf68e162e3c7e5b6e8e0eb65ef45f319f7fffafffead023406b609e90c1b108313c916161a771d80205623152668287a2a5b2cbf2dd72ec92f6f300c31b6313e32cf326233cc333334803488346c3415347933dc3230327231d33020304e2f8e2eb92dd92c252c692bab2a1a2a8229f728a92858280d28e727a52767275b274a274f277a27752750271f27a7261e26ad252025a3244324ab23f4221722c520301f761d6d1b681980177a1584138d11490fe40c5e0a820792049d0178fe70fb95f8bbf522f3c2f063ee35ec36ea3be87de6ffe49de38ae2c7e13fe11ce153e1c0e166e222e3d1e37fe421e5bbe567e61be7e8e7dbe8dde9fcea2bec37ed24eee1ee45ef7def97ef7def67ef58ef2aef0eeffdeec7ee96ee5ceee6ed69edf0ec69ec1eec18ec2fec83ecf2ec39ed78eda0ed94ed94eda6edb1edebed46ee9bee14efa4ef24f0c6f080f126f2e7f2b5f35cf40cf5c0f54ff6f3f6b5f76bf844f93dfa13fbe2fbaafc2bfd91fdf5fd26fe51fe8dfe9bfe92fe7dfe14fe6ffda4fc7cfb24fac3f82bf784f5ebf328f261f0bcee0ded89eb51ea2ae92be85de774e68be5bae4cde3f3e256e2c3e168e161e168e194e1ece11ee24be28ce2b7e20be3b3e37ce48ce5dee614e834e930eab5eaefeaf9eaa8ea44eaece962e9d3e845e86ae77ae692e57be47ae3a4e2aae1bee0e7dfdcdee3dd17dd39dc8ddb21dba6da5dda50da35da51daa9daedda61db04dc86dc27dddedd53decade46df84dfe4df74e0f0e0a6e188e23de303e4cee44ee5cee553e6a0e604e783e7d7e72fe873e85ce819e8b1e713e78ee63ce613e640e6a4e60ee770e786e72be772e654e509e4e9e2fde173e162e17de1bce119e24be27ce2dde24de319e47de54be7b6e9d4ec43f005f408f8dcfb86ff0203ff05bc08740b100ef8105b14f717e51bfc1fb92324271f2a622c392ebd2fcf30d631df32b6339b345b3593356d35bf346433e6316830fb2e262ec92da02ddd2d212e1b2e132ecc2d2a2dac2c3e2cf42b5a2c4a2da52ea430cb32c934cd368138e339663be13c693e554057425c4488466548d749ec4a404be54a164aa348db460745f642ec40063fe43cb03a62388b356332f92e0c2b0f273723511fc31b8b183415ea118e0eb20aae06a3026bfe8afa32f72ff4d1f10bf06fee17ede0eb76ea1ae9e4e7bee6fee5b2e5a5e5f3e576e6e3e64fe7aae7d5e702e83ae86ae8bae81be969e9b2e9dde9c8e97be9e9e800e8d4e675e5f6e374e208e1b4df68de20ddd6db7bda2bd903d8f5d619d682d511d5e7d430d5ced5d7d65bd808dad8dbe0ddecdf25e2cee4bae700ebc2eea0f290f6a2fa78fe2002d3055f09f20ccd10a6147918471c981f542290240a26ee268727be27c227c12783270d276c2671253524df226221e61f841e2e1dfd1bfb1a1a1a6719cc182e189517f2165216e01591156d157f159a15c9152a16ab166c177c18a219d71a0e1c121df91dc71e4d1f9c1faa1f4d1fb61ef81d001d021cf81aba197c184217f215bd148213f3112310f40d4f0b9908f4055d031301f5feb8fc76fa14f86ff5cdf23af0b0ed75eb98e905e8e5e61ee67ce506e59ee42fe4e2e3c0e3d1e33ce4efe4e1e513e74ee877e990ea76eb32ece5ec7eed14eebfee5ceff9efa3f032f1aff117f232f20af2a5f1e4f0f3efedeeb6ed79ec43ebf5e9c2e8b6e7aee6cfe513e549e4a3e32ee3cde2bbe2f1e232e39ee324e496e433e509e6f8e636e8bbe94deb0eede7ee9ff057f2fff369f5c9f624f861f9b9fa2afc80fdccfee9ff9000d300a900f4ffedfeb1fd35fcb8fa52f9e7f79bf66cf527f4dff29bf13ff0f9eeefed09ed61ecfbeb9feb53eb1eebdaea9fea7fea54ea2eea1dea05ea09ea48eaaaea4aeb26ec07edf5ede9eeb4ef7bf04bf104f2ccf2a4f34ff4e4f45bf579f569f53bf5c8f447f4d5f344f3c6f26ff204f2a4f152f1c4f018f063ef74ee79ed92ec86eb73ea69e928e8d1e681e50be4a9e28fe1a5e027e02fe06fe0e2e065e18ee176e13be1c5e075e083e0c4e06de184e2abe3fae462e67be769e83ae9b6e93dea04ebd2ebe1ec28ee36ef21f0e0f015f1ecf072f062ef02ee81ecceea45e913e8fee61de64fe53ee4f9e27fe1bbdfefdd3ddcb0da89d9c8d85ad841d83ed82cd812d8d2d794d79ad7e2d7a4d803dac7dbfedda1e050e315e6f5e8a6eb68ee6af171f4b4f73ffba3fefa014a053508f90aba0d2a108e120b155417b219361c7f1eb520cb225b24a725ba265b27e6276a28ad28052965298129a529ae2956290729b8284c2848289428f328c529c42aa22bc02cdd2dbb2ed02fed30f2316e333e353b37cc39903c313fed415b44464617489949d14a3b4ca14dfa4e8b50df51cd527d538853ff523e521051b14f704efd4c744bf1490148b9452a43e93f323c3a38c5333e2fe12a6f264e229c1eff1ac217dc14d211df0e050cf7083006e003ca0145003eff32fe4efd82fc71fb6bfa7bf956f84af76ff695f509f5d3f49af46df42cf488f3adf2b1f17bf03beffeedaaec69eb49ea32e92be81ce7d6e559e4b5e2fde060dffbddcedcdadb1bdb8bda29dafcd9f5d9f7d902da21da5bdae1dacadbf0dc47deb6dffde036e287e3dfe473e666e87beac7ec61effff1b3f48df736fac2fc5cffcb013c04e9068509190cbc0e1a1145136d155c172c19071bb21c431ee21f6121d52250249825b526a8274828b028ec28ee28e928e928e128ef28f628c7286828ad278d264d25fa23b722cd212121ab2085207420622067204020e81f881ffb1e5e1eef1d8b1d421d411d4c1d701dcb1d181e591ea61ebd1eb71ec71eba1ea01e821e0d1e451d411cd81a3c19a317e31520147412af10f60e670dcd0b490aed08830737061e050004fb0210020301f3ffecfebffd8ffc67fb21faedf8edf70ef780f64ef649f678f6ccf61ef781f7f3f754f8b3f803f933f956f961f94cf924f9d2f855f8cbf72bf78ef616f6acf55df539f51af508f509f5e1f493f425f46ff39cf2ddf11ef185f01ef0aaef35efcbee43eecfed8fed58ed42ed52ed47ed40ed5ded6bed8dedc9eddeede9edf9ede0edcbedd2edbeedaaeda1ed64ed15edc5ec42ecb7eb47ebc8ea6aea47ea22ea0aeaffe9b7e951e9e6e847e8a7e720e776e6cae527e555e486e3d7e21ae287e136e1e1e0afe0a8e086e078e096e0a2e0d5e041e1a4e12ae2dae264e3f6e3a0e426e5c7e5a2e679e77be89de985ea4febfbeb54eca4ec0bed54edaced07ee10eef0eda6edf4ec1cec2bebe9e99fe866e712e6f6e425e460e3dce29be255e243e26ce285e2bde215e33ce366e3a7e3c4e3fae357e49ae4f5e473e5cfe53de6c6e628e79ee737e8bfe873e950ea05ebbceb68ecc5ec19ed72ed99edceed09eef9edd0ed8aedefec46eca1ebd1ea1cea8fe9f9e893e85de814e8cce771e7d4e617e640e53ce42fe315e2e6e0c8dfc0dee4dd5add06dde7dc04dd31dd89dd35de13df3fe0bee136e3b3e446e6bce758e94ceb54ed90ef0df275f4fcf6c9f99efcbcff2f0392060a0a960dd9100b143217fc19aa1c431f7e21b023d62598273c29ad2a962b532ce12cff2c1a2d2b2df32ce12ce32cb72cc62ce92cd22ce42cf92cd62cf32c2f2d592de52dae2e872fe5309a327734cd363c39783bc53dd13f8a4168433c450b473649614b5e4d5b4fd750b0512952f1512d514550fd4e824d1f4c784aa848e146bb445a42e73fef3caf396a36dc32662f462c22293b26a023d7201b1e7a1b861886159112510f300c6109a60660049e02f900a2ff95fe74fd84fcd9fb30fbc9faa2fa70fa5dfa5cfa29faeef99df9fff841f855f718f6cef485f337f227f14af078efbaeee4edc6ec7feb0eea71e8d5e637e586e3d4e113e03ede76dcc0da22d9b3d77fd68ed5e7d491d48cd4c5d438d5edd5ddd61ed8c7d9afdbbfddeddf02e2fde30de621e83bea73ec92ee90f09ef2b0f4eaf687f955fc3bff4a023505e5077c0ab80c7d0ef10fed108811151294121413b9133f147c1484142f147f13b712e4112311ab107c109810051194111e129812e6120313fe12dc12a0124412d0114b11b11015108a0ff50e500e9f0dc70ce30b1f0b8c0a500a860a040ba60b400c8c0c7a0c030c170bec09a30846070d060b053f04ca03a903bc0303045a049904c604cf04b104a1049f04a604c704d504a60436045903fe014f004ffe1dfc07fa24f887f65cf598f42df423f44ff497f4f2f427f51bf5d2f42ef440f335f20cf1e0efdeee08ee74ed3aed38ed58ed8aeda0eda4edb9ede9ed4eeef1eea9ef67f01df1a1f105f255f265f247f2fdf164f1aff0f8ef3befa1ee3deef9edf9ed49eebfee5eeff8ef3bf03af006f09bef42ef13efe2eec8eeb3ee72ee44ee41ee41ee6deebceef2ee43efc1ef49f013f113f2f6f2d0f391f4f7f434f555f51bf5b0f424f443f34cf263f166f084efd2ee1cee87ed29edd4ecafecd4ec19ed97ed54ee11efcdef74f0c2f0c4f085f0ebef20ef46ee52ed79ecd7eb55eb1deb25eb34eb57eb6deb3aebfceacfeaa5ead2ea5debf0eba2ec5aedbdedf4ed0deec4ed56ede4ec40ecc0eb96eb8eebe8ebbeecbded02ef86f0cef1d5f28ff398f318f34cf214f1bcef80ee32edfaebf4eaefe918e97ae8d8e767e72fe7f8e6fee64ce796e70be8a9e813e962e9c1e9b9e97de94de9c4e846e8fce79de767e76ae766e7a1e726e8b2e867e922ea86eabfead8eab2eaafeae9ea29eb8aebefeb0aecebeb8eebe0ea0fea24e91ce81de723e633e56ae4b4e31ee3c9e297e29fe2efe24ce3b8e337e4a0e42ce509e617e791e884ea9becf4ee9af147f42cf758fa7cfdb800ff030007f009de0c950f5f124515fd17b91a631da81fc321a82324259226f3271b29652ab42bce2c082e392f1c300d31d9313432823298324132f831a3311d31ef30ed30db3028318d31c1313f32d3324d33353453356c36fc37b239433b0e3dab3ece3fea40ca416c427c43ca443d4645485f4a3b4c304ebf4fb9509151d05153519a50484f654d8b4b7149fd46a844fc41d13eae3b3b388c342531a22d212a242738247a21511f1e1dc41a7f18bb159312870f500c3209a40643042902a60048ff1afe4bfd69fc85fbd9fa1ffa91f970f969f98cf9ebf923fa47fa6efa49faf6f987f9c8f8f4f741f795f628f608f6ebf5d0f59ff513f53ff42df3bff11ff066ee8cecbeea14e98ce751e675e5e7e4a7e4a8e4bde4d2e4f8e442e5c3e59ee6dce758e9feeac6ec93ee79f094f2cef427f795f9dbfb02fe2500220218042a062508120a140cf70dc50fa2115c13f3148116d017dd18be19471a781a651aee1926192a180617e515d814da13fe12251241117f10cc0f100f5a0e730d4e0c2f0b1f0a4209e108d708fe0822090d09a808fe072c075106b80553052f05860537064107d408c20ad40cf30ed21046125613e9130a14df136613c01222128f111911cc1081103510f10fa40f5c0f2b0ff20ea80e3e0e890d820c2a0b76098b078905770376018cffadfdfefb8dfa49f942f86cf7a5f6f3f55bf5edf4cef4fcf46af511f6b4f62cf78cf7d8f725f8abf864f93cfa27fbf3fb91fc13fd6afd9cfdb8fda0fd5ffd0dfd99fc32fcfffbd8fbc2fbb3fb60fbc6fae1f974f8a6f6aaf476f263f0ccee9bede2ec91ec35ecb4eb12eb24ea32e979e8d2e75ae724e7ebe6c9e6dfe6f4e615e746e73be7f6e68fe6efe559e504e5dfe41be5c0e579e63de7ebe733e841e83de807e8e2e7f4e707e831e867e85ee841e82ae8dce775e703e763e6dbe589e53be51de52ce51de50de5fce4b3e459e4e2e319e34ae293e1dfe086e08de0a7e0f0e04ee188e1e8e17be217e3fee318e510e61ce739e821e91bea27ebf6ebbfec8eed28eed3eeaaef7af07bf1aef2c5f3dff4f0f5aaf635f79bf79ef769f700f727f60ef5bff313f254f09deec0ecfeea6be9d8e77ce671e594e426e422e43ae489e4fae435e560e584e56ae54de53de511e516e56de5ede5cbe607e856e9c5ea43ec8cedb6eeb1ef44f096f0b3f08af05ff045f01bf0f7efbeef3def99eee2ed12ed50ec96ebc1eae4e9fce813e858e7d6e69ae6b4e606e77de70ee897e824e9c9e96aea1eebf1ebbeeca2eda7eeaeeff8f0abf2a1f4f9f6a2f937fcb5fe10010503cd0488060b089c095b0b120df00e08111a134a159417b219c21bac1d251f50201a215b2176219121ad212222d22277233924e0244a25d9257426ea267d27e727ec27e927cd279d27d5274d28d428b129972a582b492c332df42dda2eac2f56302f310a32df32f83310351b36583783389c39e03af93bd53c943ddf3dbd3d623d8a3c583b0d3a67388e36bb34a8327730482ec12b042941263e234020811dbe1a2c18e815a3139311d50f150e8b0c500b0b0ae208da07990658053804f802e20116014c00aaff30ff80febdfd04fd2afc70fbf0fa6cfafcf99bf90af95ff8a6f7c6f6eaf518f539f476f3d1f22cf29cf112f17ff0faef7fef04ef9aee24ee88edd4ec05ec38ebaaea73ea99ea16ebbbeb5aecdbec30ed6ceda4ede1ed2aee6beea5eef2ee59eff7efe7f004f22af346f421f5b6f530f68df6edf695f781f8b8f955fb21fdf0feae000d02ee027303980375034a031803ed02f80225036903d5034b04b6041e0568058e05a805a80582054405dd045a04db035f03e902900247020f02fd010e0239028602ec025c03cb03250466049004a704ba04e1043905d905bf06d607fb08f209930adf0ad00a720aee095009a008e40710072a06500591040304b6038d0368033703e3026e02eb016401e0006500eeff78ff08ffa6fe62fe3dfe37fe5bfe9dfee7fe3cff92ffdcff1a00410055006c008c00bd0005014d0182019a017b012801b000090045ff6dfe70fd66fc71fb92faf1f9aaf999f9b0f9d4f9c0f96bf9e6f827f855f795f6cdf5faf424f427f323f250f1a4f030f00bf003f00ef035f04bf051f056f02df0d6ef68efd3ee3deec7ed54edfdecd8ecb8ecb3ecdfec0eed4bed8eed88ed41edd6ec34ec9feb4feb21eb2eeb77ebb2ebe5eb1aec1fec18ec22ec14ec0bec1fec2cec57eca8ece5ec1ded4eed41ed12edcfec5aecddeb71eb04ebc9ead6ea10eb98eb5fec2bed0eeef1ee92ef00f035f009f0b3ef58effbeedeee0fef68ef05f0e3f0e0f11cf386f4daf510f7fff777f8a5f8a2f86af832f8f6f793f733f7def686f666f687f6c4f631f7b2f70ef855f874f83df8d6f74bf79bf612f6d1f5d1f531f6d5f67cf72bf8dbf871f902fa7efab3faa8fa63faf6f9b0f9c1f934fa0cfb17fc0cfdc8fd25fe0bfe97fde2fc0bfc56fbe4fac0faf1fa58fbc0fb13fc3efc43fc42fc49fc49fc38fcfafb85fbe8fa40fab8f96ff96cf9a9f918fa9afa24fba6fb09fc54fc85fc92fc91fc83fc4dfc06fcb7fb5bfb2afb4dfbc7fbb8fc09fe66ffbd00ee01c1025503bd03e5030004200435047604ed047e05560665078208da095f0bde0c6b0ede0f03110a12e9128f134c141615c9159d167a172e18e5187419ac19cb19c7199f19b419fb19501ae31a7a1bdd1b471c9e1cce1c221d781db71d281eb11e411f232034215922c8233d258926cc27b72822294e291b299328172891270f27e226de26f6265d27cc27242885289f286028012856277a26b825df2404246223bc221d22b1211b215620861f651e1a1df71bd61ae3195719e8189e18951875183b18f4173c171416a214c012b110ca0ef50c650b500a850918091c0947099009ec090c0af009a60900091508fb069a052304c30271015e00a3ff16ffc4feb5feb3fec2fee1fedafeb4fe80fe29fecefd90fd56fd28fd12fdeffcc5fc9ffc62fc10fcb2fb29fb80fad7f931f9a9f85bf83ff856f8a9f826f9bef966fa09fb95fb0afc6dfcc6fc23fd8efd04fe83fe05ff83fff9ff6100b200e900110134015f01a30101026b02e1025603bd031b04640478044804c903eb02cd019d0073ff65fe7dfdadfcf7fb77fb3ffb62fbe7fbb7fcbdfdf2fe3a008201c202c7035e046f04df03b30227016dffb5fd35fcf6fa01fa6ef931f935f972f9cef938faadfa17fb7afbe4fb33fc5ffc6dfc3afcc9fb36fb6efa85f99bf89cf7a9f6f6f57ff563f5bff567f653f76ff86bf937fad0fafbfacffa67fa9bf992f877f720f6b3f458f3eef1a8f0bcef00ef8fee7fee86eeb1ee12ef60efa8efefefd9ef6befb7ee7fedfdeb79eacfe834e7d8e57be438e33be250e191e00fe082df09dfc8de91de91ded7de12df4edf81df61df1cdfc9de37dea1dd1edd81dc16dc03dc1edc98dc5fdd14dec8de63dfa8dfebdf40e07fe0f3e093e11be2cee29ce33ae4d6e44fe554e51be5b2e40be494e365e355e39ae312e470e4d9e438e563e5a5e5f9e53be6a8e62ce786e7d9e703e8d2e784e72ce7c3e695e6b2e619e701e858e9f8eaf6ec18ef12f1e3f25af460f529f6aff6f4f63ff78cf7ddf767f817f9cbf987fa15fb60fba1fbe3fb42fcfbfcf2fd07ff380047011002a802f102e402b602710224020502100234027002aa02d202f90220035303a30308047f0404058505f5054e067e06810660062a06f105c305ac05b005c505e80521066906bb061007430745072407ed06c106c206f1064607b5071b0860087d085f08fc075e078f06b005ee045304e3039a034603ce024902bf0143010401fd000e01360162018e01de015402e5029b035504f3048605fc054406790681064f061406e405cc050b069d065f0757085c094b0a3e0b200cd00c660dc90de40dd50d920d230dcd0c970c810cbb0c2b0db20d680e180f960f031048105910721088109210c610041130117b11c8110e12881209137913041469148514a014a0148114a81404157b1541161617cc179d185a19ec19a01a421bb71b431cb51cfa1c661dd91d481efe1ec01f66202621c7213122a522f7221a234a2358233e23412347235823ad230c246324cb24fe24f324cf2457249923d622f4211a2193203a200d201a20172002200220ec1fda1fe21fa01fff1e131ea91cf11a3f198517ed15a31475137712db1175114911591152112b11f3107510bf0feb0eca0d6b0cf60a6009e707c506e60555050e05c9047a041404650385029d01bc001700c1ff9effabffc7ffb7ff80ff18ff72feb3fdd7fcd0fbbffab2f9bcf80ff8b6f7b2f712f8b4f873f937fabbfad0fa6bfa74f90af883f60df5d7f306f379f212f2c3f162f1f8f0a3f05bf02ef027f023f029f049f063f07af097f09bf094f093f080f069f051f009f0a0ef37efcfee9eeec0ee0aef74efefef43f082f0bbf0d0f0dbf0e1f0bbf092f081f06ef080f0bdf0eef01ef14cf155f157f14ef114f1d2f094f03cf002f0ecefcfefd4ef00f027f069f0b7f0cbf0b4f063f0b8ef03ef77ee0fee06ee56eebaee45efe0ef4cf0b9f03cf1b3f14ff219f3d8f3a2f45ff5bcf5c3f577f5b7f4cbf3f1f22bf2c4f1d9f130f2caf28bf31cf47cf49cf442f492f3a1f256f101f0e6ee00ee8eeda3edf2ed6feee7eefbeeb7ee1eee0dedd1eba6ea88e9cce894e8b1e838e902eaa0ea1aeb6deb6beb5deb70eb8bebdaeb52eca7ecfbec5aed9bedf7ed78eee2ee5eefeeef4cf09ef0edf001f102f1edf088f0ffef60ef83eeabed04ed70ec26ec34ec5eecb7ec27ed64ed80ed76ed12ed83ece1eb19eb74ea12ead9e9fae970ea01ebbaeb80ec1bed9fedfced19ee36ee65ee9eee13efb3ef46f0ddf05df1aff10cf27ff202f3c4f3baf4c0f5e0f6f9f7ebf8c4f972faeafa53fbadfbf5fb4bfca1fcecfc3dfd85fdc0fd01fe3efe75febbfe0bff70fffbff9a004401ed017a02e3022603390334032a032403420394030f04ae045f05fe057906bb06c706cb06df061a07a20776088509c60a060c100dcc0d110ed90d5e0dce0c580c3d0c850c250d110e0c0fe30f8b10dd10ca106d10c40fd90ed50db70c920b9f0ae2096109390948096b099e09b909b509b409aa099f09b409cd09e109010a0c0afe09f709e509d109eb092d0a960a340bd40b5b0cda0c3a0d7e0dc70dfc0d0b0ef80d9d0dfd0c470c750ba10afc09750917091b096b09fc09df0acf0b9f0c5b0dd10df20df00db40d490df30c9e0c4e0c450c560c640c990cc40cda0c240d830dec0da50e7b0f481041112c12db128113e813f9130414f013c213d31302144314e314b1159116c4170919331a6d1b711c191da41de31dc91dac1d751d2d1d2f1d5c1d9f1d2b1ebe1e3d1fe21f7a20fb20a0212522682297227022e62148217f20a11f011f771efa1db71d711d261d101dfe1cfa1c3c1d811dc41d211e4c1e461e4a1e2e1e051e011ee91dc01da31d481db51c0d1c221b141a1a1915182b177516ae15d914fe13e812bf11ad108f0f890eac0dc20cdf0b100b2d0a5c09a908f50769071607db06d106de06bc066e06e005f604e403bd02850174008dffc3fe38fedffda1fd86fd5efd04fd82fcb0fb87fa30f998f7c9f505f453f2d2f0c5ef1cefcaeedfee22ef7cef01f081f0f0f067f1b3f1c1f1a6f136f173f083ef5aee20ed19ec41ebbaeaa2eac3ea0beb72ebb7ebceebb5eb3eeb80ea95e972e85ee78ce6eae5a1e5bae501e68be651e714e8dfe89ee906ea2bea12eaa5e931e9dde8a3e8c1e840e9eee9e1eaf5ebd6ec91ed12ee2fee2aee21eefeedf3ed02eefded09ee25ee33ee65eebeee0fef70efcdeff3ef01f0f9efc3ef96ef7eef6bef94effbef81f048f13ef227f312f4e4f46ef5cbf5eaf5adf543f5b8f40ff49af369f368f3c2f356f4e5f489f52bf699f6f9f63cf737f720f7f9f6abf673f656f636f643f679f6b9f630f7d8f782f846f90cfa99fafafa17fbc0fa15fa1ff9daf78df663f561f4b4f35bf32bf32ef34cf35cf370f382f378f36ef35cf31ff3caf254f2adf100f163f0d9ef94ef9cefd6ef53f001f1b1f168f212f38bf3e2f315f419f411f407f4f4f3fcf31df43cf472f4b7f4f1f42df561f574f573f54ff5f7f48af411f48af310f39bf211f280f1e8f04bf0d8efa6efb3ef03f073f0ddf036f16df174f168f15ef166f1a0f11bf2cbf29ff379f432f5bef522f66cf6bcf624f7a0f729f8aff820f980f9ddf944fac3fa5dfb03fca1fc27fd81fda4fd96fd63fd17fdcdfc97fc7dfc8efcd6fc51fdfafdcbfeacff87004b01d7011102f4017701a800baffdbfe39fe00fe2ffeadfe64ff2800d3006501d701270267029402a802b002af02a902b502df022b03a3033c04e904ab056c062607de0782080f0994090a0a780af40a6d0bd30b1e0c2f0c040cbb0b5f0b020bc30a8f0a5d0a450a3e0a480a780aad0ac40ab90a700aed096909f208900870088308b9082b09c309610a130bb60b300ca10c000d470d980dd70de40ddf0db80d7a0d720db00d350e1f0f3a1053117212671310148e14c614a7145b14d51320137c12df115511181110113511b0114d12e6128713f2130d140514bd133a13bb12221276110211bb10ab101411c711a112ae1390140f153f15ed1428145a139b121d123a12ce12ac13d314e915bb165f17a5178e175717ef1675164016451693164b172e181c19251afe1a901bea1bd41b4d1b8f1a8e1973188217a216df155015c4144114e4137d131113b2122e129211fb104a10940ff50e490e9a0df40c340c6d0bb40af0094009c50876087308c4084009e109840ae00ae80a8c0ab3097e080c076c05da0383027b01e600be00d900230166016d013001910088ff39feaffc03fb6ef9fff7c9f6ecf55af511f51df55bf5baf530f67bf67bf629f663f53ef4f4f292f14df05befabee4eee4dee6cee97eec6eec4ee98ee56eee1ed53edc5ec20ec8beb2eebf1eaf9ea55ebcdeb66ec20edc1ed4ceebceedaeeb7ee66eecfed26ed92ec05eca2eb76eb62eb7bebbfebf9eb30ec58ec47ec18ecdbeb7eeb33eb12eb0beb42ebb6eb3aecd6ec74edebed54eeb2eef1ee3aef8befc8ef14f075f0d9f064f10af29ef230f3b2f3fef33df47bf4acf401f57cf502f6abf664f7fcf783f8e9f819f946f981f9bdf927fab2fa30fbb1fb26fc70fcb5fcf3fc0ffd28fd30fd07fdcffc8ffc43fc1efc27fc4bfca3fc17fd76fdcffd0dfe10fef4fdbafd5afdfefcaafc4efc04fcc9fb90fb82fbb2fb1efcdafcc8fdb7fe9aff4d00ac00cf00be007b003100edffa4ff66ff27ffd5fe8dfe57fe37fe49fe84fecbfe17ff51ff5dff46ff07ff98fe10fe7afde4fc77fc3cfc2bfc42fc64fc78fc7efc75fc5dfc40fc1afce5fbb1fb84fb63fb5efb6efb85fba0fbb4fbc0fbcefbe2fbfdfb25fc5cfc9efcf0fc56fdcdfd4ffed5fe54ffc1ff15004a005e005c005000440043004e005b006400600045001600daff8cff37ffedfeb8feaafecefe1cff89ff06007800d40019013b013d012c010f01fd000c014501b20157022103fd03d6048d0519067f06bc06e2060d0747079d070d087d08d80810090c09d90896085608390855089708ef08440969095009fb086308a007da0625069f05630562059305e8053b068106bb06d506ca06a0064806cb054c05d9048b047f04a104e10439058f05da052306550668066c065d06460647065d068406c306020738077607b207e1070408ff07c60773070e07aa066b0648062b061206db057305ea043c047703c6023302d101c101ee013c02a302f40210030103bc024e02ec01a9019e01f2019102600350042b05ca052f064b062206de05890533050a050d053b05a3052406a0061c077907a807c207be07980770073c07f806c50699066f065b0647061c06ea059c052b05c2046804260429046704d0046c0512069806fe0624070007bb0660060a06ec0506065306e906a70772084709fe09790ac80adf0ac30aa40a8e0a920ad70a510bf30bc30c980d4d0edd0e210f0f0fc10e390e880ddc0c390cac0b510b170bf60afe0a150b340b630b800b770b3e0bb20ad309c908ac07ac060006a905ae050b0693062707b8071c0842083208e4076907e4065a06de05850544052105260542057605c1050e065a06a106ce06dd06cc068c062806a70508055b04a303df021b0257019500e2ff3aff90fee9fd36fd74fcb6fb00fb62faf6f9baf9a6f9b7f9ccf9cbf9b0f966f9f3f86ff8e4f767f719f7f1f6ebf608f723f72af71ef7eef6a1f650f6faf5b4f596f595f5b7f501f650f694f6c1f6b4f66df6fdf55ef5b0f417f497f351f359f398f309f49af418f571f59cf579f51bf593f4d9f30ef352f2a9f136f110f11cf15ff1cbf132f294f2f2f22ef35cf386f394f39bf3a4f39af398f3adf3c6f3f9f347f48ef4d8f41ff545f562f57ef58af59ef5c3f5dff500f624f62af61ff603f6c6f586f557f52df51ff52cf533f53ff54cf542f536f52bf505f5d7f4a4f45cf41df4f9f3e4f3f5f329f460f49ff4daf4f0f4f3f4e5f4b7f489f466f443f43bf44ff462f47ff49bf497f486f46df443f42ef438f455f498f4f3f445f593f5ccf5d4f5bef589f52cf5cff480f43ff432f459f4a2f418f5a9f532f6b7f622f757f762f741f7f2f69ef659f62cf637f678f6d5f654f7def759f8d1f83cf988f9c1f9def9cff9acf97bf93df90cf9e3f8b6f891f86ef847f835f836f845f870f8acf8eef845f9a6f907fa6ffaccfa11fb4dfb7afb9bfbc7fbfdfb40fca6fc2afdcdfd9dfe86ff780069013802ce022a033f031a03d80287023c020d02f201ea01fa0115023f027f02c30204033b0352034d033b0320030f03100310030703e802a0023e02db0187016a0196010602bb02a00391047f055206ec06540787078807770763074e074c0750074a0749074a0752078107d8074c08e3088209100a910af40a320b5d0b6c0b5d0b440b1a0bdd0aa50a680a260af709d309bb09c109d209df09ed09e109b909940970095a09690985099d09b509b709a709a1099d09a209c109e709170a670ac80a390bbf0b330c840cb20ca10c550ce80b520bac0a1b0aa4095a094e095f097809890969091709a8081c088d071507a5064006e5057905fd047c04eb035c03de026502f40193012f01d500950064004f005d007900a500e60028016d01b501ec0113022f023a024002520269028e02c602030342038103aa03b4039e035903e9025b02b20101016100d6ff6eff2fff08fff2fee9fee3fee5fef5fe0cff20ff2cff1efff8fecbfea5fe9cfec2fe15ff89ff1100950004015e019e01cb01f5011f024b028002b702e702150337034d0364037f03a403df0326046d04ad04d404e004dc04d004c404c504ce04da04ef040905270552058405bb05ff054a069906f0063f077a079f07a30788075a071907ca067b063006f705e605fe054006aa0622079a0704084e087108710850081d08ee07c507aa079b0789077107590744074107570778079a07a9078e074107c40618064f057c04a803e40233028f01fc0079000400abff6eff49ff3cff3bff38ff32ff1dfff5febcfe6dfe08fe99fd20fda5fc3bfce9fbbefbccfb13fc8bfc27fdc8fd55fec0fef9fefdfed1fe6bfed0fd0dfd2bfc44fb78fad3f967f939f938f957f984f99ef995f960f9faf878f8f6f782f734f713f713f730f765f7a2f7e9f73ff897f8f8f862f9c3f918fa56fa6afa5bfa31faf6f9c9f9bdf9d2f907fa4afa7dfa93fa85fa4dfa03fabbf97ff96df98ef9def95efaf9fa8bfb00fc40fc3efc0efcc5fb76fb3cfb20fb1ffb42fb8afbf1fb78fc0bfd8cfdf0fd2ffe4efe6dfe9efee7fe4dffc0ff2c008e00dc0008011101eb0095002000a6ff3dff03fffefe27ff77ffe1ff5200bf00170143013d01010199001c00a2ff39fff3fed5fedffe0fff5bffadfff3ff15000400bcff48ffb3fe10fe71fde4fc79fc3bfc2afc40fc73fcaffce7fc16fd37fd4dfd58fd4efd28fdebfc9ffc5cfc40fc5afcb0fc37fdd5fd6ffef3fe4eff7bff7eff58ff17ffd2fe96fe73fe70fe7cfe88fe8bfe7cfe63fe54fe54fe65fe85fea2feb3feb8feadfe8ffe63fe1ffec6fd63fd00fdaefc83fc81fcaafc01fd76fdfdfd8cfe0dff71ffb2ffc6ffb2ff8aff5bff38ff35ff4fff7bffa7ffb5ff92ff41ffc8fe3ffec4fd63fd1ffdfbfce7fcdafcd0fcbcfc92fc51fcf1fb7bfb0afbaffa84fa9afaedfa6ffb0efca9fc25fd73fd87fd6dfd40fd1afd16fd46fda2fd14fe89fee3fe16ff27ff1afffcfed9feb1fe83fe55fe28fe05fe01fe21fe68fed0fe42ffa7fff3ff15000e00e9ffaeff6bff32ff0bff03ff25ff6bffcfff4000a300e000ea00b8005700e7ff80ff42ff3bff61ffa1ffe1ff0200faffc8ff73ff10ffb9fe7bfe66fe7efeadfedffefbfee9feaffe60fe14fef1fd09fe5dfee3fe83ff18008a00c100ad005600caff1fff77fee3fd72fd2ffd18fd25fd56fd98fddbfd18fe3dfe42fe2efefafdaffd61fd1bfdf7fc0ffd63fde4fd7cfefbfe49ff60ff41ff04ffc7fe91fe70fe72fe8efec7fe19ff65ff9cffb3ff95ff52ff02ffabfe66fe41fe31fe3dfe5ffe7bfe8cfe86fe55fe0dfec5fd88fd77fd9efde5fd46fea8fee6fe05ff06ffeafed4fedefe0bff76ff1e00e700cd01b80283033504ca043b05a70515067a06e2063d077607a007c207e00721088308f9088809170a8a0aeb0a2a0b3d0b3d0b2b0b0a0bfc0a000b120b3e0b6f0b8f0ba30b9b0b6e0b360bf70ab90a9c0a980aa20ac30adf0aea0af50af70af30aff0a120b2d0b640baf0b0a0c7b0ce00c260d4c0d440d180de50ca80c620c170caf0b230b850ad5092a09a2083e080408f607f807f707e807b0074907bf0611064e058c04ca0310036402be01220197002100cdffacffbbfff5ff4e00a700ec000a01f500ae004300c1ff41ffddfea8feb0fef4fe64ffe7ff6000b600dd00d500a60061001000bfff71ff23ffd0fe71fefffd7ffdf4fc68fceafb7efb25fbddfa9afa4ffafbf99cf938f9e5f8aef89ff8c2f806f953f991f9a0f974f918f99ff82bf8e2f7d1f7fbf75bf8d8f85ef9e3f955faaffaf6fa29fb53fb8afbd3fb30fc9bfcf9fc39fd58fd55fd45fd45fd59fd88fdcffd22fe82fef7fe7eff1400b00033018b01b00197014901d300370084ffd1fe34fed2fdcbfd27fedefed2ffcb009a011c023902fe018701fb00870052006a00d4007f0146020803a6030b0439043c0425040704f103e403e503ec03f603fe03ff03f603e303c5039d036c032803d0026202e30166010101c200b900e1002f01960105026902b602db02cd0294024102f001c401cd0109026d02d7022d03640373035d0337030b03e602d802da02dc02d1029d023702b2012601bb009900c4002c01b30125025b024702e1013a017700acfff2fe67fe15fe0cfe59feecfeaaff7000000135010a018700d9ff37ffbcfe78fe6ffe90fed2fe37ffabff18005f004f00ceffe8febcfd8efcacfb44fb6efb21fc26fd40fe2fffafff98ffe6fea8fd1efca9faa2f95bf9fbf95bfb2afdfefe650024013801c40009004fffb4fe48fe0dfee7fdc1fd8dfd34fdbbfc3ffce2fbdafb4ffc3dfd77feb3ff9100c7003f0007ff62fdb1fb4cfa82f980f93ffa8dfb1ffd90fe88ffd5ff66ff5cfefffc97fb6ffac0f999f9f3f9b3faa3fb8dfc47fda1fd7dfddafcbffb4dfac1f851f732f68df564f5a8f542f60af7dcf7a1f836f984f984f935f9adf821f8bcf7aaf704f8b7f894f966faf5fa26fb08fbbafa69fa3efa40fa65faa2fae1fa1afb4cfb64fb4dfbf8fa5bfa87f9b0f807f8b4f7caf733f8cff885f93ffaf6faa8fb44fcb3fce6fcd7fc99fc56fc2dfc34fc6afcbafc0ffd6bfdd8fd6ffe3dff2800fb007301560197005cffeafd92fc91fbfffae2fa35fbf6fb21fda3fe3e009a01540227020a013aff26fd48fb0bfab3f960fa10fc9efec1010505d607a009fc09cf08630652035c0035fe56fde9fdc5ff7a026f05f80776098009fe073a05d801b2fe93fc01fc10fd5fff440202050007ef07c707b5060c052a0371014000dcff5c00a1014e03ed04130687064c069a05bb04e50332039c02130297013c01210164010402da02a3031204eb031d03c101110062fe01fd2afc00fc81fc82fdbefeddff8f00b0005500c1ff50ff3fff8dfffcff2a00c0ffabfe21fd8efb6ffa22fac4fa38fc32fe470007020c03ff02bc015fff46fc14f985f632f574f536f7faf90afda4ff2c016301640090fe76fcaafa98f984f975fa2cfc46fe4400a9012b02bf01950015ffacfda3fc20fc1efc78fc0ffdcefd99fe60ff05005f005800e9ff19ff12fe00fd0cfc63fb2cfb7bfb60fccefd8eff5201b90261031e03ff014f0098fe68fd26fd02fedbff4a02d8040d0788082009cd08a207e305e90321020801fa000d0210048106b4081a0a610a8b09f7072206770441038c023602220235026b02e002aa03d004510602089d09d30a440ba70afa087906a9034001d5ffb6ffd900d402170523079e085a09560990080e07f404810219003ffe55fd89fdc2fe9f00a3025d047505c1054405150464028000c5fe96fd48fdfbfd8cff9b01a0031a05b90568054f04bd0202016dff41feb5fdebfde0fe5700d901d502d702b901c6ff9cfdf4fb54fbe2fb54fd22ffbc00b601e50155013700d0fe75fd7cfc3bfce8fc7bfea500da027f042505ba048b0326022101d0003101f501a702e6028b02a0015a00fbfeb1fda9fc0bfcf7fb89fcc4fd79ff5601ef02d103af0374023c0069fd8efa4af834f7abf7a7f9c1fc46005a035305dd0501052203d30097fee6fc12fc40fc80fdadff650216051007ac079c060b0496003afdf6fa72fadffbd7fe7f02de0514088c0831076004d4008dfd81fb5afb47fdd7000f05c808000b290b61094806c102b7ffcefd47fd1afeecff3a02810445062f07240736069c04b002c6002eff2afed7fd27feeffee0ffb4004b01b0011202a60270034104c804b504ea0397021801d5ff18ffe8fe20ff90ff10009b003b01ee019502fb02e00230020e01caffc3fe36fe1ffe4bfe7afe8cfea0fef4feb8ffe4002402fa0209033b02d1004bff1afe79fd65fdaefd20feabfe4bff0700db00ab015902d2020b03ff02ab020002fe00c9ff9efecafd8cfde5fda4fe7eff28008b00c100ec00290173019d0188013c01da009d00a200c100ae001a00e2fe45fdbffbc3fa97fa28fb22fc42fd7cfeecffbd01d003980559067d05ee024fffbafb3bf974f85df95dfbc6fd19002402f6038d05ac06f9062c064404b80140ff82fde4fc5afd78fec5ffdf008d01d101b0011c011400a6fe0afdb4fb1ffb93fb0ffd2dff4201b602280388021c014cff7afdfffb11fbc2fa15fbe8fbeffcdefd70fe7cfe19fe7afddcfc7bfc7bfce2fcb0fdcafee9ffb700ce00edff2efe09fc2cfa44f9a8f931fb61fd93ff44014702b402b6027202e8010701deffadfed2fdb0fd6afebeff26010602f401f90086ff37fe99fdddfdd0fe0c0031010e02b7025003de033204fb03ee021a01f5fe3afdb4fcdbfd9b0058041a08d90ae10b000b8c084a051f02c3ff9ffeb4feb5ff4001fb029a04e805ad06a1069a059b03f20038fe1dfc1ffb60fb97fc29fe7dff2e0021007fff89fe69fd3bfc14fb17fa84f99ff97bfae9fb7bfdacfe24ffe2fe29fe61fdd9fc97fc78fc57fc2afc19fc5dfc05fde6fdaffe13ff07ffd2fed2fe4dff2f0009015001b30045ff85fd21fc8ffbe5fbd7fcddfd8dfec5fea5fe73fe70feabfe11ff89fff7ff52009500ab007200d8ffddfeabfd85fca1fb1dfb05fb5efb3cfcbffdd9ff2b020c04ae049603fb00c4fd3efb7dfac7fb6dfe2d01c502a3021a0110ff6dfda1fc74fc60fc0efc9ffba3fbb6fcf9fee5017f04c905440528032e0031fddefa80f924f9cff974fbeffdd6006a03d30488049302aefffffc8bfbcefb99fd2f00ac026404ff0479040b030101c6fee7fcf4fb5bfc30fe0401060455065307e90690050104e7029e021103e403a8040f05fd049304fe036c03ff02c502be02e7022e036f038203340366022401a5ff44fe66fd55fd1dfe8eff38018d020f037102b7004bfedefb3ffa1dfabcfbd3fe9702f005d307aa0785051f02a5fe45fcc0fb20fdb8ff660219043504ce028a0035fe5ffc29fb5dfabff964f9b3f91efbc0fd15010c048505de044d02d6feccfb3afa7efa37fc90feb7002a02c702bf026202f101a601a501f601870219035203e502bc01050033fec1fcf7fbd2fb01fc14fcbffbfbfa05fa4df938f9fcf994fbbbfd0100e701ff02f802d101d2ff81fd80fb57fa3cfa15fb8cfc33febafffc00e7017a02a80259028001220053fe41fc2afa59f831f715f738f88bfa9cfdb3001a0358044e043503640122ffb2fc5cfa88f8c0f770f89ffae0fd65014f04140698061506e20440034b0131ff45fdf5fb97fb22fc17fdc6fdaffddafcebfbc4fbfafc6eff470249047f04b10270ffdcfb14f9c5f70ef89cf9e8fb7cfefa000603490477047203760108ffc2fc18fb2cfacff9c4f9f0f961fa3efb8afcf8fd09ff45ff71febcfca5fab9f869f7eaf635f725f87ff9ebfa0afc8efc5dfcbdfb3cfb6afb8efc70fe5a007a014701c0ff71fd30fbb2f95df931fadefbfafd1400c101ab02a502ba014000c1feb9fd6cfdc8fd68fedefee5fe68fe8bfd76fc3ffbfcf9dff83bf87df8e3f93dfce6fe0501ea0179013900f3fe46fe47fe74fe24fe03fd4efbcaf942f909fad2fbe1fd74ff3d0070007f00c6004101900148013d0094febafc28fb2afae4f963faa7fba8fd3a00f4023f058d0680062205dc024100edfd5efcd9fb7efc44fee500eb03b806a7084d09aa081c074a05da03250323038303cf03c0035d03eb02c9023f0343048d05bb067907b1079507730795071408c208450940097608f206140568038502de0285042c07390ae10c740e900e2c0da60aa507d904d402e401ef0195025e03e003fe03ef03030479044c051d066d06f305bc043a0310029f01e3017d02ed02fb02e80237035c045b0698081f0a2e0a8f08d3050b033101b8007101b002d803be049a05d40696087b0abe0ba00bc8098d06d602a1ffa4fd1ffdcffd3afff900bd026004d405fd06be070308af07a906f704bd02620093fefdfd0bffa201f504d4072c096408b5051002a9fe94fc72fc3efe77014f05cf08130b8b0b0c0afa063403b8ff4ffd50fc74fc23fddefd70fe17ff51006b024a055e08c30aa90bb90a17086c04af00befd37fc5bfcf9fd91007f031206bc073c088707d4059003320138ff14fe01fef4fe9a004d0263038203c202c6017301630288041507c40883081806390251fed5fb84fb2ffd0000f8028b05c907010a460c240e9d0ec10c59081f02a8fbc3f6b1f4bcf547f91dfe000308079a09630a500984068c0265fe31fbddf9c4fa73fdef00270450062307c5068005a003790176ff23fe0ffe70ffec01b704d806ab073607fa059a04760377024f01e8ff92fef1fd8ffe5c009a023e047b044c037c0124000d00450118038804e9042704be026501a500a40042013c0253035c041b0545059704f2028a00e9fdc1fbaffa0ffbd9fcabffed02e305d7073e08db06d603ccffa3fb52f89bf6d5f6ddf835fc1f00cc038406c4074d074a05450206ff5dfcd8fa96fa49fb64fc57fdd9fdf8fdf5fd1efe95fe33ffa5ff97ffe6fec3fda7fc17fc6cfca4fd58ffee00df01ef01450149005cffb4fe4bfeeefd80fd19fdfbfc70fd96fe3900e201ff021c03160239001efe83fc08fce3fcc6fef8008f02d902ad0170ffe6fcd9fac5f9bdf98ffaeefb95fd45ffa5004801e4008affcffda9fce5fca1fe260128037903be01a7fe8cfbbef9caf93dfb11fd43fe62febafdf8fcb1fc1ffd0dfe08ffb0ffceff4eff51fe1efd21fce1fbaffc58fe26000e0137009ffd36fa6bf794f61cf84bfbcafe48011a0280013b00fefe30fed4fdbffdf1fd73fe10ff60ffc6fed5fcdef9e8f641f5f5f524f9e8fde702d806eb0803094f07fd0367ff22fa1ef5baf121f1aaf3b0f8a1fe91032206d4050903e3feb3fa95f76ef68ef77ffa3efe5c017a02260103fe79fa2df803f8a4f9fafbb6fd11fe4ffd3efc8afb7cfbbbfbb5fb55fb07fb62fbe2fc4bffa201d9023602aeff20fcbff88cf635f6a4f719faaafc69feaffe94fdb7fbe7f9f5f818f9d7f993fabbfa2bfa69f909f93af9cef92dfacdf9d8f8f2f7cdf7ddf8c6fa85fc38fd6cfc5ffafff730f65df59df59af6d8f71af91efa80fa05fa93f864f644f408f324f388f471f6cff710f830f7aef568f4edf34bf460f5daf65bf8b3f98afa61faf9f867f639f383f02aef6fef08f122f3eff44bf683f7e9f888fabbfb7efb4af96df519f114eea2ede5ef01f464f88cfbdcfc84fc2cfbb6f9a7f808f8b9f770f7e0f6fff5dbf4a0f3c6f2b8f29ff374f5c2f7d7f94cfb07fc32fc36fc3efc0efc53fbcaf97bf7fbf4f8f2e2f1e4f1b2f2c6f3e3f400f627f777f8d2f9d1fa2efbcefadbf9e1f869f8baf8e5f98efb0dfdd4fd7bfde0fb72f9e7f6fcf45bf426f5d6f699f87ff9e8f8fef68bf4acf284f291f46cf822fd66010e04a5045703b2007dfd51fa86f77af585f4e3f4baf6a2f9a5fcbefe34ff06fe2afceefa3efb3efd0e003e02b9022b011afea0fab3f7c3f5ecf416f53ff6a6f852fcb200b7040d07c206ef03afffa5fb4cf91ff96ffafefb97fcbdfb11fac6f8f4f811fb8ffe1e026c049e04ae0273ff10fc7bf93df832f8d1f899f936faaafa52fb7efc38fe3400c90141023a01cffea9fbc9f800f7b9f6e6f707fa81fce2fed6001a027602b901f5ffaffdb4fbdcfa89fb57fd4cff5d00f3ff57fe7afc4efb42fb05fcc7fceafc73fc08fc89fc5efe1601b3033905420556047c037f037904af050006bb040102befe3ffc68fb4ffc66fec0009b02c0035104830487045b04f20373031303f2020d030b0384027101200030ff51ffb300f4026d0569078208d4088e08c60776067a04fd01b6ff88fe2affc801920523093e0b280b0e09fc05230371015d019e0291049b061c08c208a708ff07260795066e069106cc06b6061806240522046f036503f903fc045106b8070d09490a1d0b330b740ae208e4064505a0044a052f078d097b0b5a0ccf0b200a2708a5062506da064808b909af0ac50a0d0a0909180880077707d6078908b009380b120d2a0f0c115212e712a7129911d30f1b0d5209d504540010fd72fc04ff4604ca0a6d109213ec133c120f10ea0e280f2510d6103810380ecd0b0d0abe09e90a7d0c420da00ca00a3708cf0633076e09df0c3e108412691317134112c011c2110b1233129d112810630ee90c590c000d4c0e5b0f7f0f4e0e350c5b0abc09fc0a1b0e0f1289158b176d175e154e121b0f970c550b380bf60b4b0db30ed70fa410e610b9108c109e10271140126113f413b413931221114d107b107e1197127c127310f00c34091c074108c20c64131e1a911e631fbc1cb2170912760db20ab609090ac40a530bb00be30b3f0c280d800e09108c11a21238139913df132e148e148814bb131b12a80fd90c730af308c4081c0a8c0c630fcc11ae127211660e780a480773067c08bd0ca3111c15ef1547143011270e3c0c490b8c0a5d098f07e5058705e5068909420c890db80c6a0ade077f0612071a097e0b290d480dd50b58095c0682037d01cc00e401d904d908990ccb0e870e130cbe08fe05dd047105b9068a073807c005dc037502e8012e0204030d043d05a206f507c5089e0839070405eb02be01d801d202a80384033c025300dcfecdfe59000f030e0657085409e008120756044e01b1fe4cfda7fd93ff39025204a904ee02e7ff0cfdf0fb5dfdd900fe0425081c09c107db049001eafe67fde6fc0bfd71fdd6fd3bfebbfe68ff58008401bf02bf031d047a03c9015cffe3fc3cfbf1faf4fba8fd19ff77ff8bfebbfcd6fab0f9a8f99ffa21fca4fdd6feb6ff5d00de0035013301b700dcffd2fed9fd1dfd85fce5fb21fb43faa2f9aaf97efaf3fb89fd7cfe3afea3fcfdf9f2f64ff4aaf268f2a5f30ef61ef91afc16fe6cfef5fc15fad5f677f4c4f3e9f44af7abf9f8faa4fac5f828f6d1f376f288f200f44cf6ccf8d5fab1fb0efb0df921f636f338f193f047f1c2f203f46bf4ddf3a5f297f170f151f2fbf3c4f5c1f687f621f5e1f27df09aee76ed48ed18eeb3ef22f243f57af824fb7bfcbcfbecf8bdf436f0adec02eb32ebcfec06efe6f023f2c5f2cef281f2eef1e4f09bef78eeceed1fee88ef82f180f3dbf4faf4f9f336f206f019eef6ecc7ecd7ed17f0dbf26ef5e4f65cf6dcf30bf0dceba1e819e71ee74fe805ea9beb2cedf9eef6f016f3daf476f5aef49af287ef40ec5de913e7cee5c7e5e6e641e971ec7fefb9f193f2dcf15cf00fef97ee66ef21f1c1f289f3dbf272f0eeec23e9d3e508e44de46ee6f4e9d0ed9bf098f191f0f2ed0aebffe84ee81de9cfea63ec75edf5ed05ee45ee00ef0bf059f1a4f28df31bf429f463f3d3f188efb9ec3eeac9e898e8d0e901ec5fee8ef059f29cf381f4d8f42df46ff2b9ef84ec00ea22e938ea22edf5f051f460f6bcf686f5abf312f242f1a1f1f6f296f405f6b9f646f6e5f4edf2c5f034efc6ee9cefc4f1d1f4eef770fab7fb65fbd3f988f707f501f3c0f11cf10ff171f1fef1c0f2a3f35ff4eff442f550f56ff5daf587f671f73cf860f8bcf75af672f4b4f2bef1d4f118f335f564f7fdf86bf95cf830f67af3c4f0adee66edb6ec90eceeecd6ed99ef50f29ff508f9cbfb23fddbfc0cfb09f88df43df191ee2bed6ded50ef9ff2a2f629fa3dfc34fcf4f945f649f209ef5aed59ed73ee05f05bf1f2f1e8f199f15af19cf17df2b8f304f5f7f533f6c1f5d3f4b4f3f3f2e7f292f3edf4a0f623f827f978f9fff802f8caf68df592f4e8f372f33af33bf36df3f7f3d5f4d5f5dbf6acf716f82df811f8caf765f7b6f686f5e1f3faf13ef052ef88efcaf0caf2f8f4ccf61df8f7f882f9f5f94cfa71fa6bfa42fa09fad8f97af99df817f7f0f49cf2f2f09ff0eaf18ef4b8f773fa0dfc43fc5ffb01fab9f801f825f81af9b4fab4fcb8fe68008701f001b7010601f7ffb6fe6bfd2bfc2afb8dfa49fa47fa5cfa68fa96fa3bfb9afcc9fe6a01cc035505a405cc046003e901ab00bfff08ff78fe65fe46ff770106055809630d2b10e410500ffb0bc407b603e900f9fff8009203df06d109b70b3b0ca60bc80a4c0a8b0a750b5b0c7c0c870b7c09d90682041d0303034f049d066b09520ccb0e7c1051111e11f10f300e2e0c5f0a60097209a10ad00c650fab1114131613a211430f9b0c7f0ab9095b0a040c1a0eab0f2310920f420ed70c000ce10b570c2d0df90d9f0e580f281015111812c412cd1240122011ad0f560e3c0d870c6a0cc10c700d5b0e010f0e0f870e7b0d5e0cdb0b250c280d930eaa0f0010a80fd40eff0da40dac0dd90df80dc00d5d0d530dd40de70e55106c11aa111411ea0fd40e7d0eee0eda0fc91012118f10b20fe30e880eca0e290f100f300e5e0cfc09d1075f060706fc06e5085b0b030e3e109e11fc112d11780f960d1f0c9b0b540cdc0d820fac10ce100010ed0e230e120ed90ee70f95109d10ec0fe20e1f0ec20d9f0d6c0dac0c580bff0924093a09670a1b0cae0dca0e380f330f430f7c0fb80fc80f4a0f3a0e0e0d260ce60b8d0cb50dd20e800f4c0f280e870cc50a5409ae08cd088c09cf0a340c800dbb0eb20f42106910df0f8e0ec70cd30a37099d082409950a800c000e640e980dce0bc10975085f088209870b880dda0e6d0f5d0f190f1a0f310fe70ee20dcd0bff087106f50420050807d109650cf80dff0dad0cd50a21091a08090899086f096d0a650b630c980dcb0eb90f3610fd0f2b0f430e940d670dea0dc70e9a0f2b101d10550ffb0d130cee0924081e074107c4082e0bc60de10fd7109210860f1e0ed10cf30b620b040bee0a1a0ba50b9a0c930d250e090e040d5c0bca09e4082a09cc0a540d11105312631308138411350fb10c8f0a0809320808084308b6084e09d909490aa80acb0a8d0ad7097e08a906db04b403f5031006a909cc0d3d11c81203127a0f450ca30952081f084508ec0791068704cc025402ac039b06110ac90ccb0db30cf0098506740390013f016302a1047d07580aa80cfb0df80da90c890a4608a3061b0691067a07220802081e07f9052e052b05ee05fd06d6073d0847085808c7088509210a0c0ad8089d06f603b701a7002401fe02a60564088d0aba0bd50bf70a5f0963075005750323029d010d0272038705d807df09250b7d0b0a0b140ae908b7077a061e05ab035d029a01b301b4024804cf059a064706e004db02e30098ff4cfffcff5301d3020104840449047d037602a4016501d401d102180455054506b9069306b8050a0488017ffe8cfb71f9dff820fadafc31000f0389043c0459027cff75fcf7f969f8e9f74cf82ef92dfaf3fa53fb74fbaffb50fc7dfd0fff97009e01d8013e011800b3fe36fdbbfb50fa0af937f82cf803f98ffa50fc9ffd0efe7cfd0cfc26fa3bf8a9f6dcf52cf6b6f75cfa85fd2e007601ec00bffedafb60f919f837f845f97cfa5dfbc8fbe9fb25fca1fc1efd55fd19fd65fc85fbc2fa2bfab5f93ff9b8f85df872f8fdf8d9f98cfa87faaaf940f8cef610f671f6d8f7eaf91ffcebfd08ff44ff72fea5fc13fa25f7a4f44cf36af3eaf42cf737f960fa6ffa99f97ff8abf741f72ff719f798f6a9f574f427f319f277f134f159f1e8f1c8f2f7f358f5a1f6a6f738f82cf89ff7b0f673f52df418f354f22ef2d5f227f4eff5baf7e4f80bf910f828f602f451f287f1e4f127f39ff4b6f5fcf530f59df3ccf143f094ef04f064f15ff361f5bef62ef7b3f67df518f402f36af27bf229f327f451f585f683f73ef8aff8bcf87af8e0f7bdf61df51ff3f7f04defcfeebbef06f219f5e9f7b0f908faf6f81ef72df57ff355f2a0f116f1b1f07df075f0dbf0e1f179f3a5f527f856fa98fb68fb83f968f6f3f2fdef52ee21eedceeedefcdf014f1eff0b6f092f0b6f020f18cf1f8f15bf28af2a2f2b1f29ff292f299f27af22af294f190f064ef70eedeede2ed56eebbeed9ee96eef6ed75ed6dedcfed98ee97ef6df022f1c7f137f26bf22bf21ef167ef58ed51eb03ead2e9a0ea54ec8ceeaaf063f269f35ef35bf2b0f0caee7eed61ed76ee79f09bf2cff3adf340f2f1efbced6fec4fec7ceda8ef28f288f440f6cbf628f68ff46ff2acf0e5ef21f031f168f2f7f2b4f2e8f112f1f4f0d5f15ef322f586f613f7f3f660f678f577f456f3f1f195f0a1ef61ef33f0fff136f459f6dff76ff839f877f756f62cf514f412f387f2b8f2adf35df54af7a6f8f0f8eff7e7f5b7f326f295f114f21af3e3f317f4abf3ddf247f247f2dff202f461f5a2f6aff767f8a7f878f8d2f7c2f6a8f5d6f47af4c7f48ff559f6cef6abf6daf5b3f499f3e5f2e8f294f39bf4c3f5c0f659f7aaf7cff7dcf7fbf72df850f85df833f8a5f7baf67cf511f4ddf23bf262f272f31ff5d3f60df865f8b9f76df61ef55af48ff4b5f563f71af95afadefaccfa68fae1f956f9a6f895f729f6a1f469f309f3bef352f552f723f943fa96fa31fa43f912f8cdf697f5c7f4a8f457f5bef671f8cff96dfa37fa77f9c3f884f8c1f83ff98ff95bf9bef816f8c4f717f8fdf810fae2fa1efba4faa7f976f860f7adf673f6a2f62bf7f0f7d6f8e0f908fb2dfc26fdb1fd93fdd5fcb8fbaafa25fa50fafafab8fb08fcaefbf1fa55fa61fa5cfbfcfc94fe71ff23ffccfd0afc95fafbf964fa70fb89fc37fd31fd86fc81fb6dfa98f93ef979f961faf4fbf8fd1500e001ed021a03870278015a008fff41ff85ff52007a01c402dc035f0423042d03b901540087ff90ff7200de014c035c04cd048c04dc030803500205024602f702fa030905d9056a06bf06d906d706aa062e068505ef04ca048e0541076c09780ba30c7d0c5f0bec09d908bc0881099e0a920be50b830be80a7f0a900a440b4a0c1f0d800d2b0d290cf50af1096e09bd09b80a030c6d0d9f0e700fff0f2810b90fb40efd0cc80ad708c107f4079e09260cb70ec210d511fb11be115b11e3106810a30f840e700d980c280c420c7e0c7b0c420cde0ba00b0e0c210d920e23104d11da1115121412fa11fd11d6116211db105210ff0f2d108f10ca10c11042108d0f450f910f57104d11ad110811b00f1f0e1f0d720ded0efe100f136114cb14c714931462144f14f0131e133612801171116412e4134c15301624165b1592142a145c142915e8151e16c815e214d11338133113b513ae1491150b162b16d215291594140b14911349130313c712e2123f13dc13be147015a4157215d7142314e1131414a814841528165e1659161316ac15641506157614dd1324136512e81183112011f010e61031112a12a0134115bb1666170217e9156014e8121812f0115312411365149215c31685177d17a616eb14b612f5103810dd10ef129715dd171719b218d0164b14e3115b104f10831172139615181788170d17c2150d1498129b114711da111213a3144a165d1771179f160d155a137612bd122b147416a418f219231a211951177315d613b312421242128e123313df136014bb14ab14261473139912c31146111e1158112012321350145515c41562155c14c112eb10750f930e710e3a0f9d104212dd13d414d014e0131712f70f4a0e6f0d9c0dce0e6a10db11cc12dc121712dc10590fd60da50cc10b430b5e0b020c310de80ea210d1110112b810090eb00a9007ad05b7057407250acb0c510e560e320d6f0bba098b08c4072f07ba0660066c06320794083b0aaa0b490cec0bc90a25096a07e70597048903e902d4027403d2049b065f08a7090f0a9b098f082c07c70595049103c2023e0210024f02e9028a03d3036a032402460063fe1afdf8fc14fe07002e02d1036704d6035f027700a6fe55fdc1fc09fd0ffe8fff3b01a1025b033d034802b700f4fe58fd2cfc91fb6ffb9afbe1fbfdfbc9fb43fb73fa90f9ddf879f871f8b7f810f94ef953f90af98bf803f88ff76bf7c3f783f891f9affa6cfb85fbe6fa99f9fbf77bf668f50df57af56af694f78cf8c6f815f891f686f4a3f294f199f1abf257f4d4f59df678f66bf5f2f389f263f1b7f08bf0a9f016f1d3f1aaf28af34ef4a8f49df44af4bef343f3f9f2b0f25df2e7f119f12ff076ef05ef17efafef6af012f16cf132f190f0beefd0ee20eeddede0ed37eeccee48efa3efd5efaeef5eef09ef98ee38eef9edaaed6ced47ed07edd0ecabec66ec3aec4eec7eece5ec6beda6ed7aedd4ec8eeb0ceaade894e732e7b5e7d5e87dea56ecb2ed55ee21eefaec6ceb0bea11e9e0e873e94fea46eb23ec8fecb7ecb3ec49eca6ebdceac3e9ace8dee755e75ae7f8e7d4e8dce9c2eaf4ea65ea1ae90ee7f0e467e3bae251e314e546e777e931ebf4ebfeeb95ebbdead3e9f8e808e86ee77fe730e8ade9a5eb35edf6edb4ed65ecccea8ee9c3e884e86ee8d6e7d6e6c2e5d7e4afe463e558e641e7cce7b0e769e75fe788e7fce772e856e8c3e7f2e605e69ae5f4e5c4e6fee75be958ea0aeb86eba9ebc2ebe7ebcfeb96eb2deb4cea40e945e859e7eae61ae794e74ee8ffe820e9bbe8eee7cee6f9e5d9e55fe6a0e741e986ea3feb55ebb0ead6e927e995e856e85fe866e89ee81ee9b4e97bea4eebc3ebf4ebf6ebb3eb81eb78eb4ceb16ebd8ea73ea3dea67eac3ea5bebf2eb15ecd9eb5deba8ea38ea50eac1ea90eb83ec25ed7eeda2ed8aed93eddfed2dee7eeeafee7cee1deeb5ed24ed92ecf6eb1aeb50eaf3e92aea3eeb05edd1ee2df0b5f037f037ef47eea1ed8cede8ed3cee7deeb7eeeaee60ef1df0cdf057f1a1f189f15bf148f13af148f161f156f158f186f1bbf102f23af21ff2caf159f1c4f02bf081ef9beec1ed56eda5ed0bef57f1bcf376f5e8f5e1f40ef361f196f028f1dcf2ebf4b5f6c3f7e7f77ff7f9f697f6acf63df70af8e3f876f96cf9c8f8b6f783f6b2f586f5e8f5b2f68af720f886f8def83bf9acf9fff9dbf927f9f7f7a1f6bcf5b6f5abf677f88cfa39fc0afdcefcbdfb7dfabaf9e8f922fbf8fcb7fecfff01008eff16ff1affbfffba0061012601f3ff33feb0fc2efcf6fcc5fee7008c023303d702cf01b100f8ffc4fffdff5b0090008b006800590099003201f0019902f002db0298027c02cb02ae03f304310621079807af07c8072408c7088909fd09c409e3088e07300667058905a506a8081d0b660d000f650f600e560ce109cc07ed06710701090e0bc60ca80dca0d660dd80c8b0c800c9e0cfd0c8c0d450e370f0e107a1081102c10d00ffd0fb910b1117a1272126111c90f400e6c0dd30d2f0ff110ae12e9138514dc14081519153a153215e81493142b14be138f1381138813c813061419140c14a113d712131280115e11031234139a140616fb1642170e175b164d154414391338128e1132114011101285137815d217f719631bf51b791b281ab9188717d916e81638175017121746162415521409145c144c15371691164b164a15ee130713e2129a132a15d91604188618311849177e16fa15ce1515166c16a8160d1788171a18dd1859193f19bf18ec172a171a179c174f18e018a7187b17ef1575149213c013a414bf15d9167d1792177217061748167a15841494132f135a13031426153216cd161d171717e316e016d61693163716a3150715f4146a154c1687178518eb18e1185e189117e8163d167415c714191489138313dd135814e114001596141414a31381130114c4146b15f0150f16d915bb159915541505156b1497130f13f21251133e141f157f156315b214c3135013841369140916c6171819c9196a19f517f215b913da110b114a115912ed133915bb158515971453136112e011d3114a12d1121c133c130813a3128112a2120913c1134a144114a6135a12ab10490f7e0e820e7a0feb106612c313a51409153c153215f714b91441148913d4122212a1119911d81121124612c9118310c10ec30c150b5f0aaf0ae50bbd0d880fd61091119b111e117110980fa80ed80d1d0d990c8c0cd60c5e0d170eb40e1f0f790fac0fb60f960ffd0ed70d610cdd0ad209c609af0a3a0cda0dc10e8a0e5b0d910bda09d808a8081d09dc09560a500ae5093f09b9089d08d4082a095909ff080608aa063f054c0442042905c6069b08f109560ab50941088a062905670449048a04a9045d04a403b90216021d02db0219045b050e06e705ed046803dc01bb0035004800b80038019701c401c901ce01e401fd01f7019501a70035ff77fdd6fbd6fac1fa99fb0bfd81fe6eff89ffd4feacfd92fce5fbd0fb4efc1bfdf2fd9bfee1feb2fe1afe28fd14fc1ffb66faf9f9d3f9cbf9daf916fa87fa3dfb1afcbffcd4fc29fcb8fae1f829f7e4f550f566f5d3f561f6e7f633f746f72af7d6f676f63ef63ff694f623f792f7b0f770f7e0f669f668f6e4f6c0f79cf8ecf87ef865f7d7f556f44cf3cbf2dcf250f3bdf3f1f3c9f31df323f226f14ff0ebef10f077f0f0f044f135f1f5f0cbf0d0f031f1def177f2e5f228f331f33bf355f336f3c5f2f8f1d3f0deef9bef1ef05bf1d3f2b5f3aef3c4f227f179ef23ee12ed41ec99ebfdead2ea76ebdcece9ee1af19af213f374f2cef0b9eebeec11eb18ea08eab9ea2eec21eeedef3bf1caf16df19bf0d3ef40ef1def44ef27efabeed9edc8ec0bec05ec99ecaaedccee4bef00eff7ed47ec90ea51e9a2e8c2e8a0e9ccea2bec89ed7eee0fef32efadeeb8ed7fecfaea8fe984e8dae7e5e7bfe81beae3ebc1ed16efc2efbaeff7eefced2fed8dec34ece9eb27ebf3e984e81be780e62fe7f5e883eb0bee76ef6def06eea5eb55e9dee75ee7e3e70ae92eea45eb5bec4eed42ee05ef07ef37eeafeca3eae0e800e814e832e9fbeab1ec04eea8ee48ee2aeda9eb09ea04e90ee911eaf1eb19ee98ef10f066efbaeddeeb88eaf6e96beaa7ebf8ec0aee94ee53eeabed06ed94ecbfec88ed78ee5cefedefdeef75efedee38ee7deda4ec6aeb1fea2de9e0e8b5e9a0ebeeed0ff061f16af184f037efe6ed26ed1fed8ded69ee87ef89f067f1f2f1d2f130f144f03defa5eeb3ee24efcaef3df008f053ef6bee8fed46edb7ed95eeabef95f0d9f086f0c6efc1eefbedbfedfaedb9eec3efaff071f1f5f117f207f2d6f168f1f4f09af060f08ef039f128f247f351f4dcf4e7f475f486f374f27ff1aff03ff034f05ef0c6f051f1c6f13af2adf205f360f3b0f3b4f365f3b3f29af182f0d3efc7ef9df028f2e1f367f564f6a5f671f60bf690f532f5f1f4b2f4a4f4e2f45ff517f6c7f60ef7e3f65ff6aef531f505f5fcf401f5f9f4e5f414f5b6f5b3f6daf7c1f800f99bf8c3f7bdf6eaf570f53bf54df59ff527f602f724f858f97cfa59fbc2fbc1fb66fbc8fa25faaef97bf9a4f90bfa6dfaaafaaffa95faa2fafdfa92fb28fc6cfc2cfc9bfb20fb21fbd9fb0dfd33fecdfe9afec5fddffc76fcd0fcd4fd02ffc2ffbdffeffeb2fd97fc13fc57fc4efda0feefff0501d201700202038303d003b5030b03e3018c006affdbfe06ffcaffdf00fb01ea02ae035a04f7047d05c2059905fe041504240383026502c9028e0374044105e6056006b406f1060607df06880610069c0565057805c7053a06a206e40618075107a5072b08c4084409950997094609c7082d088d071a07ea061b07da071609990a1d0c250d540da90c560bd209c0086508b80876091c0a580a4d0a3f0a8d0a760bb00cb00d0e0e870d5c0c410bb50af00ad30bc60c3e0d200d810cc00b5b0b6a0bd90b980c660d230edd0e630f890f520fab0ec20d060da30ca50c0c0d830dd50d1e0e5f0eaf0e2f0f9e0fbf0f940f080f460eb30d660d690dd30d6a0e020f9c0ffb0f0210d10f630fe30eae0ec40e140f950fef0ff90fe00fae0f860fa30fd50ff50f11100c10f90f1e106510b11006112011ea1098102410a30f540f220f0c0f390f760fa10fc60fb30f6b0f3f0f3b0f6f0ffd0f971002115111691165119611da110e1238121512a7114311f210cb10fe104c119111e7112012321247122d12d81181111a11bc10ad10c410e51021113d11301138113b1137115111501123110411e410df103f11dc1195126e130b1442144114f5138513531351137813d9131d141114d61347137e12d6114811e510e710211184113012e1126d13e113f0138c13f7122f126211ee10bb10bf1017118411fa11ae1276133b1408157d156b15f8141914021324127c110b11f510fb10161185112912f612f613b914f714b714d3137e1241114a10db0f3b1021113f126013fb13d91335132c121e118c1063107a10ba10c2108f108b10db10a211e7121114961450141d136311e40ff60ec90e6e0f6e106d115612dc12e6129412c01187105d0f790e280eb10ebe0fe410e01145120d129a11091189104510f90f810ffa0e530eb40d700d780dcb0d7b0e3e0fe50f65107010f40f2c0f2d0e410dcd0cc50c0f0d920df00d070efe0dd30da60daa0db80dc00dd70dd80dc50dba0d870d1a0d8c0ccf0b0d0b990a750aa70a300bbe0b1d0c480c180c970bfe0a4e0aa4093909050917098b09330ae60a840bb50b500b730a3409f0072007eb06550740083509e009270af2096909d5084608d5079f078e07a107de0716082d081c08cb074f07dc067906340618060506fb050f062d0649064f060a067705ca043e041e04930460052506840633064805240424039902a1020c03a1033704a804f10418050805b70427045f038b02e00172014d0164019301c801ff0130025c027d027f0262023002f601c3018d012d0180007aff43fe3afdcbfc39fd7afe1f0081011002830107002afe8afc9cfb84fb08fcd0fc9cfd4dfef5feacff5f00d800d4001d00c6fe27fda7fbaffa70fac7fa70fb18fc70fc63fcfffb5dfbb0fa27fad0f9baf9e0f91cfa5dfa99fab9fac9facefaa9fa54fac5f9edf8fff73cf7ccf6e1f67bf755f836f9e0f911fad0f93ef971f8acf71bf7b8f694f6a4f6b9f6d9f606f728f750f776f766f718f788f6a3f5a2f4b7f3e8f262f22cf223f258f2cbf253f3f2f389f4ccf4b7f44cf48ef3d4f266f249f295f21ef373f36bf3edf2f3f1e8f038f00bf090f099f195f234f332f367f236f109f013efa2eeb2eeeeee42ef96efbcefe6ef25f04df066f05af0eaef3def73ee8bedd8ec89ec8fec1bed20ee3def43f0d7f086f070efe3ed33ec18ebf4ea9febebec59ee3bef79ef1eef3cee4fed9eec15ecdcebe2ebe0ebeeeb08ecf8ebeaebe9ebcaebbeebcbebbaebafebb0eb8feb87ebaaebcaeb0eec6eeca0ecc0ecc2ec68ecddeb2feb44ea6fe9e1e88ae8aae836e9d1e973eae9eaddea81eafbe94ee9e1e8dbe80be988e932eab0ea20eb7beb84eb60eb08eb45ea67e9a8e816e813e8abe87fe978ea4eeb92eb69ebeaea0cea3ae9ade857e87ae80be9a8e94deacdead6eaa4ea56ead4e966e91be9c4e8a0e8c3e8fee879e917ea7fead0ea17eb35eb72ebccebebebdeeb9ceb06eb87ea54ea47ea82eae1ea1ceb6eebfbeb9bec68ed1dee37eebfedd1ec8eeb8cea0eeae5e916ea6bea92eac6ea27eb98eb3fecfbec6aeda6edb3ed72ed2eedfaecaeec8aec9eecc3ec26edaeed02ee38ee56ee46ee5ceea5eed2eedeeea1eeefed30edbdeca9ec31ed24eeffeea5eff2efbeef56efd8ee2aee88ed11edc2ecefeca5ed90ee8fef48f054f0ddef22ef53eef6ed3eee00ef33f084f16ff2d6f2a0f2c0f1aef0ceef46ef56efdaef5cf0bcf0e1f0c6f0d7f052f11bf223f30bf44df4def3d1f24df1e6ef06efd2ee82efeef098f227f421f519f52ff4b9f224f12df03df040f107f304f583f641f72af753f63af53df47df32af333f35ef3b0f31cf485f4fef477f5bef5dbf5d0f59bf580f5a3f5fdf598f645f7b5f7cef77af7aef6b0f5bdf402f4c3f313f4cff4e8f527f74cf849f906fa61fa5ffaf0f90cf9ebf7d5f618f617f6e8f655f806fa78fb3cfc38fc86fb67fa43f95ef8daf7d1f73df805f915fa3afb33fcd5fc06fdcefc66fc06fccefbcafbdffbebfbeefbfcfb3afcccfca4fd90fe51ffb2ffaeff72ff37ff29ff4fff7fff8aff56ffe6fe71fe36fe5ffefbfeecfff300d80168028b025402e9017f0151017a01f101a3025e03f7036a04ae04c704c504a10457040804c903b503ee036204eb047905f4055c06d9066407e40741084608e5075007b40643062d0657069b06f5064f07b4074d080b09cd09830af40a090be80a9b0a400a0c0aff091a0a7e0a130bc20b8c0c340d8d0da20d5f0ddc0c670c160c030c570ce70c890d340ea60ec50eb40e730e200e030e140e450e9f0ee10eea0ee20ec80ec00e180fbe0f951096116c12e3121013d4123b129311e51059104510a010571165125f13f1132214da134e13fb12f7124713f0137f14a2146314ad13b9121112da112b121c133c142115ad159315e31411144c13cf12ec126f1329141d15fb15a21639178f1798178f175617fb16c71698165c163216da154715c614541412145414e4149715721615175b1776174817e116971653161b162e1654167516bc16ee1607174f17a017e9174a18661814188d17c9160216bd15ed15821682176f18fd18411906196118c4173417d816fe165f17be1718180c1892171817b2169216fa168617e51720180318b717b717ee173e189f1899180e186317be166e16d816b0179d187e19da199519071934184e17b8164e1604160b1623163c169116e9162e17821793174817e0164e16c415b415021692165f17ea17f817be17321791164a163a1642166a165616f51593152215b81496148014631478149a14d4145f15ee154b167e163d169115db141d147a1336131b131c136513c01318148614b41480141c147913cc127e127612a3120b13551368137f1385138513a51395133313ac12f6114f111d1144119d110a121712a411fd104310c80fe40f5a10e6105b115311c7101010510fcb0ec50e020f530fa60fb30f790f3d0fff0edf0e040f2f0f360f170f970ec40deb0c1e0c990b9e0b080cae0c6a0dc80d920dde0cb80b7e0ab2097509ce099f0a640bc50bb10b160b340a6d09d30872084d082908f907db07c107bc07dd07f507f607ee07d207bb07c907d607c7078c0700073f068f051005e8041a055e057d055d05e8044e04d3038d038c03c003e503d7038f0305036502e50198019901ed016902ec024b034c03e302200224014200c9ffdfff88008a016e02d502810273010b00c5fefffdecfd5efeecfe39ff10ff7cfed0fd57fd33fd5efd99fda8fd7efd30fde8fcd9fcfdfc2cfd42fd19fdb7fc4efc00fcdcfbdbfbc2fb63fbc1faf1f93bf9f3f833f9e9f9dafa92fbc2fb57fb5ffa32f93df8b6f7b7f728f8acf8fef8f7f87ef8bef7fdf65ef607f605f621f63af63bf601f6aef57cf580f5e0f59df66bf70bf84bf8edf712f706f6fbf43ff4fcf302f437f47af490f485f474f449f414f4dbf373f3fbf29ff265f27ef2f2f276f3dcf3f8f390f3d6f21df291f180f1f9f1a4f246f3a1f36bf3d1f222f283f140f16af1aff1eaf1fef1b8f154f114f1f2f00ff15bf17ff175f146f1e1f08af06df061f070f084f053f0f3ef83effbeea1eea1eecdee2fefa9efdbefc9ef80eff1ee78ee5bee89ee17efdbef57f070f020f059ef8cee19eeffed5eee07ef79ef97ef57ef9ceec1ed09ed67ec0fec09ec16ec54ecc7ec31edaeed38ee8aeec2eee5eebfee7dee33eebaed48edf9eca2ec73ec78ec7deca9ec01ed44ed87edc0eda9ed70ed36ede5ecc9ecf9ec39ed97edf8ed06eedaed7fedd6ec31ecc5eb80eb9beb0cec75ecd0ec01edd1ec89ec64ec55ec97ec1eed89edd4edeaed96ed21edb9ec4fec23ec3fec61eca3ecfaec28ed55ed84ed7ced67ed4ded02edc2eca5ec80ec7eec91ec70ec3becffeba9eb92ebe6eb7aec5bed47eebbeea7ee09eee7ecd5eb40eb3cebf3eb22ed32eef4ee44ef02ef92ee34eed9edaced9fed6ded41ed29ed0aed19ed5bed98edf4ed65eeb2eef6ee21effceebdee82ee47ee52eea7eefbee47ef60ef0def92ee29eee9ed26eee4eed6efe4f0cbf134f237f2e4f135f17cf0e1ef5def2eef5fefc4ef6bf028f1a6f1e5f1d8f16ff1fbf0b1f097f0e3f084f12ff2d4f242f340f3f8f289f207f2c5f1dbf122f29cf216f349f345f314f3bcf28ef2aff216f3daf3ccf492f512f627f6bdf521f589f40cf4d8f3daf3e1f3fbf329f45ff4bff430f575f58ff57ef557f574f5f6f5bcf6a1f74bf864f8fdf73ff767f6dbf5c1f50bf6b4f68df756f8fcf859f94bf9f2f86df8e6f7aaf7d2f74af8fef8b4f934fa80fa9afa8afa75fa5bfa31fa0ffaf6f9ecf90afa47fa86fac2faecfa01fb28fb6ffbd5fb5afcdbfc34fd64fd65fd3ffd0efdd9fca7fc90fc97fcb9fcf8fc39fd68fd91fdc7fd2bfed9feb7ff7f00e5009e00a8ff4efefbfc23fc13fcc1fceffd46ff6600190158013101d400750034002a005900a700ff004f018401a001a70197017a015d01460146015b01680156011401aa005d007b0038019e025b04e305bc069c068f050c049b02ab017401d30171020a036d039503b103e4033404ab0428059105e905280647064f062f06dc0573050805b504a404d1042805aa053b06c9065b07d30711081108c2073207a5064606380698064107fb07a80816092f090f09bf085208f607b2078c07a207e6074a08d5086109cc09180a270af709b5096f093b0945097d09c809220a570a4a0a120ab309500934097009020ae20ac00b4f0c7e0c350c950bf90a840a4e0a6b0aa60ad30af50af30ad50ad00ade0a020b570bba0b150c740cb10cb70ca00c590cef0b9f0b6f0b720bc90b450cb80c140d220ddb0c770c070cb00ba80bda0b310cb60c3b0da60d030e240ef60d950dfc0c4d0cdb0bb40be00b6d0c0f0d8b0ddc0ddf0dab0d8b0d8d0db60d160e6a0e7f0e620efe0d6b0df90cb10c9f0ce20c490db10d260e770e9a0eb30eb00e960e8a0e6c0e300ef50da90d5e0d4e0d680d9b0dec0d200e200e1a0e090efb0d110e150ee50d950d220dbc0cc10c350d030e100fea0f451025107f0f860ea40df60c970ca50ceb0c3f0da50deb0d030e130e080ee90de60dec0df70d1b0e290e060ec80d5d0dda0c820c590c670cca0c510dd90d600eac0ea30e610edf0d410dd70ca80cb50c010d490d660d6f0d5f0d500d730da40dbd0dbb0d760df80c8a0c3e0c2e0c7c0cf60c6c0dd30def0dab0d2e0d7c0cbb0b350bef0aed0a440bc30b470cd40c380d5e0d590d180dae0c600c3a0c490c9e0cf60c1b0d060d9d0cfa0b6e0b0f0bed0a1c0b680bae0bf40b1a0c1b0c100cdf0b810b1c0bb20a5f0a550a7f0abf0a050b1a0bf00abb0a890a760aa00ada0afa0a000bd70a920a6c0a650a7b0ab40ae40af30af00ac80a7c0a2d0ad30976093b09160906091a0934094309550953093c092f092409250948096e0975095209e6083e089e073207220788073208e1087109b209a00961090109940842080a08f0070308200823080408aa072607b60676067806c2061b074e074b0700078c0632060e063506a6062c079007bb0795072f07b7064306e0059c055f052405030506053c05ae0534069c06ca069f062b06a5053205f104ef0403050205d8047804ff03a6038c03bd032d04a304ee04fd04c8046a040c04bf038b037a0381039e03d3030b0430043104fc0398032903c80291029302bc02fd0247038603b003bf03a7036503020387020d02ae01770170019401cc0102021f021502e801af017b015c01550158015e016c018e01d30139029a02c0027e02c801d000ecff72ff96ff45002c01e9012b02db0124015100acff62ff6bffa1ffdbfff7ffefffd1ffa5ff6fff33fff0feb6fea3fec9fe2bffaeff16003000e6ff43ff7dfee0fd9bfdc0fd40fee0fe6affb9ffafff54ffc7fe23fe8afd1cfdd5fcb3fcabfca3fc97fc8dfc85fc91fcc0fc07fd5dfdadfdcbfd9ffd27fd66fc8afbcefa57fa45fa9ffa3efbfefbbdfc46fd83fd6bfdeffc2dfc56fb8dfa05fadaf9f1f932fa7dfaabfabffad0fadbfaeefa05fbf7fab7fa44fa9bf9e5f854f8fff704f868f8faf898f91efa5bfa50fa0ffa98f90df98df81bf8d5f7d0f7f4f736f87cf88ff86cf82df8e1f7bef7def71ef85ef870f81ff87cf7bff60df6a9f5b5f50af689f60af750f761f74ff712f7c2f669f6e9f557f5d6f477f46cf4c8f453f5e7f552f65cf61ff6cff583f566f578f574f53ef5c9f410f45df3fbf200f382f362f43cf5d9f510f6baf507f535f45ef3bdf26df251f274f2d0f239f3abf311f42ff40af4aef31bf391f247f238f275f2e9f24ff399f3c0f3a9f379f349f307f3c9f298f255f222f213f213f235f273f29af2aef2b1f28bf262f24bf228f20df201f2e6f1dcf1f3f10ff23bf26df274f25ff240f208f2e2f1dff1dcf1e1f1e6f1c5f1a3f19ef1aef1f7f16ff2cff201f3eaf26ef2caf140f1e2f0dbf021f16df1b2f1ecf104f223f256f26ff26cf244f2dff179f141f134f169f1c7f10af22ef236f215f201f217f23bf279f2bdf2caf2a3f24cf2bdf13df105f11df1a9f18ef270f320f46df426f47bf3a7f2cdf13cf115f136f1a3f13df2caf24ff3c4f304f41ef40ef4b9f348f3e0f28df286f2d3f23df3b4f312f42af41bf405f4ecf3f5f320f43df451f454f433f416f419f42cf466f4bdf401f537f556f547f52af510f5e9f4d1f4cef4caf4e1f419f554f59ff5ebf512f627f635f635f642f65cf661f658f63ef609f6e4f5e6f508f65df6dbf655f7c7f71ff83cf82ff801f8b1f76cf749f740f765f7aaf7ebf728f857f867f86ff87df888f8a9f8daf8fdf80ff907f9d7f8a4f889f891f8d6f84ff9d2f955fac1fa00fb20fb28fb0cfbdefaa3fa58fa21fa12fa31fa8ffa19fba6fb20fc69fc65fc2cfcd8fb85fb5ffb76fbbafb23fc8efcd7fcf9fcf5fcd6fcbefcc2fce2fc20fd63fd8afd8ffd74fd48fd35fd50fd9efd1cfeaafe26ff7fffa9ffa0ff74ff31ffe5feadfe94fea4fee0fe35ff8effe0ff1b003b00450038001400e8ffbeffacffcaff17008900060169019a019601680131011101160147019901ee01320258025c024f02440245025f028f02c402fa02250339033e0334031c030703fd02ff0217033e036a039f03d80310044b047c0490048a046c04490449047d04da045005ad05c6059c053e05cd0485047c04b3042705b4053906ad06fa0615070d07df0693064c061306f40506063b067f06ce060e072c0737072d0714070d0710071407230728071a07170725075507bf074b08d1083d095d091e09aa081a08990761077007b5072b08a108fb0845097309840998099b097f0958091409ba08790858085e08a108fa0843097f0995098c099709b109d5090a0a260a160afe09e309dc090c0a540a900abe0aba0a880a5c0a3b0a280a380a440a380a320a2e0a3b0a850af10a600bca0bfb0bdd0b970b2e0bbf0a820a700a7d0ab50aeb0a090b240b250b120b1d0b3b0b6a0bc10b130c410c580c3f0c050ce70be60b010c450c750c670c2b0cb90b340bec0ae80a250ba60b240c720c990c860c4f0c320c2c0c350c5b0c6a0c500c350c140c010c290c660c960cb50c950c390ce10b990b7b0bb00b0d0c6d0cd00c030dfe0ce50cad0c620c340c110cf50bfb0bfe0bf10bf00be30bd00be40b0c0c400c940cda0cf80c010dd30c720c0e0ca30b460b260b2f0b550ba20be20bfe0b0f0c020ce20be00bea0bfa0b200c320c250c170cf50bc90bb80baa0b950b8e0b780b4d0b2e0b050bd40abc0aa30a880a8d0a9f0abe0a0a0b610bb50b0b0c320c170ccd0b440b940afe09910965099609f409550aac0ac40a9b0a620a210af209f709100a280a470a4b0a340a220aff09c6098e094509fa08d808d508ee0824093f092509ee089c08560854088b08e7085409910983094009c7083c08d8079a078707a907d707fd0723082c081b080708e307b6079a078307750788079c07a107970760070107a2064e061f062e0658068606b506ce06d606e606ed06e106c4067d061f06db05c205e3053d069106ab067906ed053605a2045a047204e3046a05cc05f105c7056d051f05f304f1041705350530050b05c304710434040704eb03e103d603cc03d503e503fd031c042c0429041b04ff03e303d203bc0399036f033403f402c902b402bc02d802e602d702ae026f023c02340257029702d802ed02c80276020d02b40184017501790179015e0132010c01fe0019015901a001d501e101b8016c011901d100a50094008c0086007e0072006d006e00650044000200a2ff43ff08ff0aff54ffcdff4900a300c100a2005a00feff9cff3dffddfe82fe3dfe1cfe2afe69fec6fe21ff63ff73ff51ff0bffa8fe3bfed7fd86fd58fd61fda0fd0bfe87fee1fef9fec3fe40fe97fdf8fc82fc49fc4efc77fcb1fcf1fc24fd4bfd6afd73fd66fd44fdfffca2fc3ffcddfb9afb8cfba7fbe1fb21fc3cfc2cfcfdfbbdfb94fb96fbaefbc9fbcafb8ffb25fbb1fa4bfa1dfa38fa7dfad5fa20fb2efb00fbaafa39fae0f9c0f9ccf901fa46fa6cfa71fa5efa35fa12fafff9dff9aff96bf902f996f849f825f843f89cf805f96df9bdf9ccf9a7f963f9fef89ef85bf82bf81ef836f852f874f88ff87df847f8fcf79cf755f747f760f79ff7e9f708f800f8def7a8f78cf79ff7bef7ddf7e2f7a3f73bf7cef66af642f666f6aaf6fff642f746f720f7e6f69bf666f654f640f633f630f622f629f64cf66bf68ef6a4f687f64ef610f6c7f599f591f593f5acf5d7f5eff503f610f6f6f5ccf599f54cf509f5e1f4c3f4cdf404f542f58bf5c9f5caf5a3f55ff5faf4acf491f495f4c6f40ff53bf553f554f528f5f8f4d9f4b9f4b8f4d1f4d6f4d0f4b7f474f438f425f437f48df40ff576f5aff5a4f53cf5b3f43df4e5f3d7f307f43bf46ef494f494f49bf4bcf4dff411f538f51ff5ddf48af42df408f431f481f4eff44ff564f541f5fbf495f44df439f43af45df491f4adf4c7f4e3f4e9f4f9f414f51cf529f538f523f500f5d2f489f453f447f459f4a2f412f56df5b3f5d1f5adf574f541f510f504f51cf530f54cf565f560f55df567f567f578f594f595f58ff589f576f57df5a6f5d0f507f63af641f638f62df615f615f62bf633f63bf63af61df60bf615f62ff674f6d9f634f788f7bdf7aef771f717f7a4f654f641f665f6d0f666f7eaf74ff87bf855f808f8b5f767f74ef773f7b7f71bf883f8c8f8f6f809f9f0f8caf8a0f86af84af850f86ff8b7f811f953f97ff98af96cf953f957f977f9c3f921fa62fa81fa75fa39fafef9def9d9f902fa43fa72fa91fa97fa81fa73fa7ffa9dfad9fa1ffb51fb7afb99fba5fbbafbd7fbe8fbf3fbe9fbbffb91fb71fb6afb98fbf9fb6cfce1fc34fd47fd25fdd8fc75fc2afc11fc2ffc8dfc15fda2fd21fe6ffe74fe3efedbfd67fd10fdf0fc09fd5cfdcafd2dfe76fe99fe9efea9fec9fe03ff54ff9cffb7ff96ff3bffc1fe5afe2ffe58fedafe8fff4000c7000a010601d80097005b0030000f00f2ffdeffd9fff2ff350099000c017701bb01cf01b7017f0140011001ff001c016701d0014302a602dd02e102b8027402360212020d02230241025502630276029d02e8025003b603fd030804ce036f031503ea020f037303eb0350047b0462042704ea03c603cf03f303190440045f047e04b7040705550592059f0573052f05f004d504f90442058405a80596055c0533053d0589050e068e06cb06b4064c06c10569056b05c905740620078d07a7076507e90678062e06180640068006b806ed0615073b078207d90727085f085908090899072307d106d5061e078c0709085b0864083c08ef07a3079207ba070e088408e1080009e9089a083208f007de07fc074b089808bf08c508a308700864087d08b10801093b09430931090a09ea08fb0827095109730966092809ea08bb08ac08d7081509440966095d093209150906090d0945098c09c709fe09110afa09d6099f095c0935091a090e0932097309c209270a6d0a770a560a000a9109500946097609df09410a6a0a5e0a0a0a8e093709150933099a09080a4a0a560a140aa1094d0931095a09d4095c0ab80adf0ab50a4e0ae909910952094109380928092a09340950099c09f909480a850a850a430ae9097f092109ff08060927096809a009bc09ce09be098d095e092609f108e108df08e308fe0812091e093e0966099109ce09f009df09a8093a09ac083a08ef07da0712086f08d3083a097a098a0985095c091509d10884083c081e081f083e088308c108db08d908a9085e0829080c080a082d084608430838081d080608180842087308a308a60872082708c80770074e0754077507b107e007f407fe07f107d507c807b7079f078c076a073c071d070407f70609071d072a0734072307fa06d306a80688068f06ab06d006ff0616070e07f706cd06a00691068c06880682065a061106c605820561058005c205100657066d064d061006c1057e0568056d0581059f05a705970585056b05570554054c0536051805e704b504a204a904cb04050536054f05520533050405da04ad04820463043f041a040504fa030304230442045a046e046e0462045a044b0436041b04eb03b0037f035f0363039203ce0304041d04fd03af034c03eb02ad02ab02d80226037703a2039b0366030e03b6027b0262026e029302b002b902ab0281024d021e02f401dc01d601d601dd01ea01f301fa01fe01f601e301c40193015d012b010001e800e400e800f50004010a010901fe00e900d200b9009900790056002a00feffdaffc3ffc4ffdafff6ff11001600feffd6ffa8ff7bff5aff3dff1bfff7fed3febdfecafefafe3dff80ff9aff74ff13ff89fe01feaafd98fdc8fd25fe7cfea7fe9bfe5bfe05fec4fda4fda8fdc5fdd5fdc2fd8dfd3cfdeafcb6fca3fcb3fcdffc06fd1cfd22fd11fdf3fcd6fcb1fc87fc5ffc30fc07fcf2fbecfbfafb1bfc34fc3bfc30fc01fcbafb6dfb1ffbe5facffad3faf2fa24fb44fb49fb34fbfcfab5fa77fa43fa2afa32fa43fa59fa70fa70fa5ffa44fa11fad6f99ff965f93bf92bf92af942f972f999f9b5f9bff99ff961f915f9bcf872f847f82ff833f855f876f898f8b9f8c0f8b4f898f859f80cf8c6f77ff753f74bf750f768f78df7a6f7c2f7e7f7f7f7f9f7e7f7a7f74cf7edf68ef659f65df67df6b9f6fef622f72af71af7e4f6a8f679f64bf634f634f629f621f61cf606f6fcf508f60df616f61ef606f6e0f5bcf58df573f571f568f564f566f550f53ef53bf532f53cf559f568f574f577f550f51cf5e6f4a0f46ff460f455f462f481f490f4a4f4bcf4baf4b8f4b6f497f474f453f421f4fdf3f1f3e1f3e8f304f410f41cf428f419f40cf406f4eef3def3d8f3c1f3b9f3c5f3c9f3d9f3edf3e2f3cdf3b4f385f36af370f377f397f3c3f3cdf3c5f3a9f366f327f304f3eef209f34bf384f3b8f3ddf3d0f3b2f392f35cf335f320f303f3fbf208f30ef327f351f368f386f3a7f3a7f3a1f397f36ff34af32df302f3eaf2e5f2d8f2e2f207f32af360f39bf3b0f3b1f39ef363f32ef30ef3f0f2f6f21cf33cf36af39cf3aef3b9f3bdf39ff382f36cf349f33af340f343f35ef38bf3a8f3caf3ecf3f2f3fcf30cf409f40ff41af40ff40bf40ff402f403f40ef40af40ff420f42af448f479f49ef4cff402f518f529f535f527f51cf516f504f506f51df532f55cf591f5b3f5d7f5f8f5fff509f61af61ef62ef647f652f668f688f6a3f6d2f60df734f755f767f75cf752f755f75cf77ff7b2f7d6f7f7f712f81df837f863f88ef8c3f8f5f809f910f914f912f927f952f97ff9b2f9dbf9e8f9f1f9fdf90dfa39fa7bfabdfa01fb34fb43fb3efb2afb0cfb03fb15fb3bfb80fbd8fb2bfc77fcb1fcd0fce2fce6fcddfcdcfce3fcedfc0cfd3dfd7afdc6fd14fe57fe91feb5febdfebbfeb2feabfeb6fed2fefbfe32ff6cffa7ffe7ff250060009a00c700e300f200f300f100fc0014013f017901b301e70112022d024102580271029502c602f90232036e03a403d603fc030c0410040b040304110439047104bd040b05460572058a058d058f0594059c05ba05e605150653069506cc0602072a073c074807450732072c07310740076f07b007f1073b0878089d08ba08c308b708b608b908c408f0082b0960099609b409b409bb09c309d309050a400a690a900a9f0a910a8f0a900a970abf0aef0a150b480b710b880bac0bc70bd20be60bee0be50bef0bff0b0e0c3c0c6b0c8c0cb60ccb0ccc0ce10cf70c050d2b0d4c0d5d0d7e0d920d900d9d0d9f0d930da50dc00ddd0d1c0e560e750e950e940e720e630e540e4a0e6f0e9b0ebc0ef00e110f160f2a0f360f330f490f540f4b0f570f5d0f5c0f800fa50fba0fe20ff20fe60fea0fe50fd70fed0ffd0ffd0f1810271024103d10501052106c107410661075107d107b109c10b610ba10ce10cb10b010b110ac109d10b110c010be10d910ed10f61020113e11481163116311411131111211e910ec10f81006113e116e118511a811a91187117611551127112311251127114f116c11741193119c119011a011a311901192118011561149113a112e1153117a119111b311ad117e115e1135110d111a11311141116911721158114d1130110411fb10ec10d110d310cb10ba10c810cb10be10ca10c0109d108b106710351026101b1016103b10591061106d1050100a10ca0f800f3a0f2b0f2c0f360f630f800f7e0f7a0f540f140fe70eaf0e730e5d0e480e330e3f0e420e360e380e210ef60ddd0dba0d910d860d750d5a0d510d340d090df00ccd0c9f0c870c690c460c3c0c2d0c1d0c1f0c0e0ce80bc70b8f0b4a0b1d0bf30ad20acf0ac40aac0a9b0a760a480a300a180a040a010aea09ba0983093409de08a4087b086d0886089f08aa08ac0886083f08f2079a0747071107e606cb06c806c606be06b606970667063306ee05a6056e0538050f05f804e304d304c804ab047e044b040a04c803940369034f0341032b030e03ed02bc02820249021102e201bf019c017e01640146012a010d01e800bf008f0054001900dcffa0ff6dff3fff16fffdfef1feecfef1feedfed2fe9ffe50fef1fd9cfd55fd26fd18fd17fd19fd1cfd0ffdf2fccefc9dfc66fc34fcf7fbb6fb7cfb44fb1ffb16fb15fb19fb1dfb03fbd2fa96fa49fa01fad4f9acf990f985f96ef953f93ef91af9f3f8d7f8b2f890f876f84df822f803f8d9f7baf7aff79bf786f772f743f70bf7dbf69ef66ef659f643f63af642f630f614f6f3f5b4f576f54cf51cf5fff4fbf4eaf4dbf4d5f4b7f49af488f45ff436f415f4dbf3a6f387f361f34ff35af356f354f357f335f309f3e4f2a8f276f25ff23df22bf22ff21ff215f214f2f3f1cff1b0f176f14af13ef129f129f141f13bf12df11cf1dff0a1f077f03ef020f028f026f033f051f04ff04bf04af021f0f7efd5ef93ef60ef4cef2def29ef48ef50ef5cef6bef4def27ef08efceeea7ee9fee86ee81ee90ee80ee75ee7bee65ee5eee6dee5dee53ee4eee1deeeeedceed9bed8beda7edb6edd6ed01eef6edd8edb7ed75ed50ed57ed5aed79eda9eda5ed90ed79ed3ced12ed0eed04ed16ed3ded3ced38ed3aed17ed06ed10ed04ed0aed1fed0aedfbecfeecebecf1ec13ed1bed2ced44ed30ed1fed19edf5ece7ecf4ece9ecf3ec12ed13ed23ed45ed49ed59ed73ed62ed51ed4bed28ed1aed29ed2ced4aed7ced8bed9eedb7edaaeda3edaaed97ed9aedb5edb7edcbedededebedf1ed06eeffed0aee29ee30ee46ee6cee70ee7cee93ee8cee91eea3ee9aeea3eec0eec6eedeee0bef21ef3fef62ef5def59ef5bef47ef51ef77ef8defb0efdeefecef03f024f030f04ef079f085f096f0aaf09ff09ef0aff0b4f0d3f007f128f158f18df1a1f1b8f1d3f1d1f1dcf1f7f101f21bf246f261f288f2b6f2caf2e0f2faf201f31bf346f361f38bf3bdf3d8f3f7f315f41cf432f453f465f489f4baf4d9f402f531f54bf56df595f5adf5cff5f5f508f623f644f653f66ef695f6b2f6e0f618f743f776f7a7f7c1f7d8f7ecf7f1f7fff718f82ef859f893f8caf809f946f96df98ff9a6f9a9f9b0f9bff9d0f9f8f92dfa5efa95fac9faebfa0dfb2efb4afb73fb9ffbc0fbe1fbf9fb00fc0cfc23fc43fc7afcbdfcfefc37fd5ffd70fd7bfd85fd98fdc2fdf7fd2cfe5efe7cfe85fe8bfe96feb5fef2fe44ff99ffe6ff140022001c000b000200120038007000b000e8001a0149016f019901c601eb01090221022e023a024d026a029a02d1020403380361037b039703b703d303f90321044204670485049804b604d804f904260556057c05a405c205d405ee050a0623064c067a06a206ce06ec06f60601070b0716073c077107ab07f3072b084308530852084408490858086e08a208dc080d094b097c099309aa09b509b009bb09c709d109f509180a320a5f0a850a9c0ac30ae40af90a1c0b360b3e0b530b610b630b790b8f0b9d0bbf0bda0bec0b140c380c520c7d0c980c990ca50ca50c9b0cb00ccd0ce70c1c0d440d530d6a0d6f0d630d770d910da70dd60dfa0d060e180e130efc0dfe0d020e050e2e0e590e770ea70ec40ec50ed10ecd0eba0ec40ecd0ece0eeb0eff0e030f1f0f330f390f590f6c0f6a0f790f780f670f700f740f6f0f8a0fa00fa30fbb0fc50fbf0fd30fdc0fd40fe90ff30fe70ff00ff00fdf0fe60fe50fda0fed0ff90ff80f1310231020102e102910111011100810f50f00100310f80f08100f1006101c102910231032102e1012100810f30fd60fda0fd90fce0fdf0fe30fd60fe10fe50fdb0fea0feb0fd40fcd0fb20f850f750f670f580f6c0f7b0f7b0f8c0f880f6b0f5e0f440f240f240f1f0f0d0f130f090fea0edf0ecb0eae0eb00eac0e9c0ea10e960e770e6c0e570e380e380e310e190e140e030ee20dd70dc30da60da00d910d730d690d550d360d300d240d0d0d080df30cce0cbc0ca30c820c7f0c780c660c650c540c2f0c150ced0bbc0ba60b900b740b700b660b550b560b490b2c0b1a0bf80ac80aac0a8d0a690a5d0a500a390a2d0a160af209dc09c0099f099209800967095e09470923090809df08af0896087e08680869086408520842082008ef07c907a007770765075107370728071407f706e606d006b506a5068b06640643061806eb05d005b8059f059205800565055105340515050105e804c804af048f0469044d04310417040604f103d603be039c0375035503350316030203ed02d602c402ae0292027c02620245022c021202f301d601b801980179015a01410130011e010b01fa00e100c000a1008200680054004100310021000a00ecffcbffa8ff87ff6bff54ff44ff37ff2aff1aff05ffecfed1feb2fe92fe78fe64fe51fe3efe29fe14fefffde5fdcbfdb9fda8fd99fd8afd75fd5efd48fd2dfd14fd03fdf1fcdefccffcbbfca7fc93fc7cfc6afc5efc4cfc37fc25fc0dfcf2fbd9fbc0fbaffba8fb9efb96fb8efb7efb6cfb56fb37fb1efb11fb03fbfcfaf9faebfadafac6faa6fa8afa7dfa71fa6efa74fa6ffa65fa56fa38fa1dfa0dfafef9faf900fafaf9eff9e4f9cdf9b9f9aef99cf992f993f98af980f979f96af960f95cf952f94cf94cf942f939f935f926f921f926f922f920f921f910f900f9f5f8e1f8d7f8dcf8def8e7f8f4f8edf8e3f8dbf8c6f8b8f8bbf8bdf8c6f8d3f8cef8c4f8bbf8a9f8a3f8acf8b0f8bbf8cbf8c8f8bff8b6f8a2f899f89bf897f8a0f8b5f8b8f8bbf8c2f8bef8bff8c6f8c0f8bbf8bbf8adf8a4f8a7f8a5f8b0f8c5f8ccf8d4f8ddf8d2f8c9f8c9f8c0f8bff8caf8cdf8d5f8e1f8ddf8dcf8e3f8e0f8e2f8eef8f2f8faf804f9fff8fef802f9fbf8fef80bf90cf913f921f91ef91ff928f926f92bf939f93af93df944f93cf93bf944f943f94bf95af95af95bf962f95ff965f975f97cf989f99cf99bf995f990f97ff978f982f98af9a0f9bef9cbf9d5f9d9f9cbf9c1f9c2f9bef9c5f9d6f9dcf9e8f9f5f9f4f9f6f9fef9f9f9f9f9fef9f8f9f9f904fa06fa10fa24fa2efa37fa3ffa35fa2cfa2cfa28fa2ffa44fa53fa64fa73fa71fa6cfa66fa56fa4ffa51fa52fa60fa79fa84fa90fa9dfa9bfa96fa96fa8efa90fa9bfaa0faa8fab2faaefaaafaadfaa9faacfab9fac1facffadefadefadffae4fadefadafae1fae4faebfafbfa05fb14fb23fb23fb20fb1dfb10fb08fb0dfb13fb22fb37fb44fb51fb59fb53fb4ffb50fb49fb4afb58fb63fb75fb8dfb9bfba5fba9fb9afb8afb82fb7cfb86fba0fbbafbd6fbeefbf1fbe6fbdbfbd0fbcffbdcfbecfb03fc18fc1dfc1dfc20fc1bfc1ffc2dfc39fc46fc55fc59fc5afc5afc55fc59fc66fc73fc83fc97fca1fca7fcaefcadfcaffcb7fcbcfcc2fccafccefcd8fce8fcf0fcfbfc0efd1afd1ffd24fd23fd22fd25fd2dfd3cfd51fd5ffd6bfd72fd6bfd60fd5bfd5afd63fd79fd93fdaffdc7fdcffdd0fdcffdc7fdc2fdc7fdd0fdddfdedfdf8fd04fe13fe1bfe22fe29fe2afe29fe2cfe31fe3efe53fe65fe75fe83fe89fe87fe86fe86fe8bfe97fea6feb6fec5fecafecafecbfeccfed0fedafee9fef8fe06ff11ff18ff1eff21ff26ff30ff3bff49ff57ff60ff65ff6eff76ff7bff82ff87ff89ff8cff8fff95ffa5ffbaffccffdeffeaffeaffe1ffd9ffd9ffe2fff4ff0d002a003e0045004100360029002200270036004e0066007a00890094009700960097009b00a300ab00b300bc00c500c900d000da00e100e800f300fc0005010f01180122012d01330138014101460149014f015401590163016d017801830189018a018f0192019801a501b401c301d401e001e601e801e501e301e701ef01fb010a02160222022d022c022702280229022d023c024d02600276028202850285027f0277027b0283029002a202b002b802c002c002bc02c002c502cc02db02e902f40202030c030f03150319031c03220325032a0334033a0340034d03540356035c035e035e0366036e037703880393039a03a703aa03a403a603a803aa03b603c303ce03de03e503e103df03d803d203dd03ed03ff031a042c043004310427041704120413041d0430043c0441044b044c0447044d04540456045f04650467046f047304770486048d048e04950495048c048a048604830490049c04a404b204b704b304b204ad04a704b104bd04c704d604dd04da04d604cc04c004c004c004c104cd04d204d104d904db04d804df04e204e004e504e304db04de04df04dc04e204e404e404ea04e804e104e504e404df04e404e504dd04da04d604d104d704d804d804e204e604de04dd04d704ca04c704c104b904bd04bf04bf04c804cb04c704c904c104af04a704a2049e04a904af04af04b304ab0497048c0483047a047f0483048204870485047a0476046f04640462045f04570454044e0448044b0449044104400439042c04240417040a040b040b0408040e0412040d040704f903e903e403df03da03e003e103d903cf03bc03a303990391038c039603a103a103a003950380036e035f0356035d03640365036903630353034403320321031d031a0316031a0318030f030a030103f502f302ef02e702e402dd02d002cc02c702c002c202c102b902b202a50293028702810280028a029302950290027f026602530244023f024c025a02620266025d02470232021f02130216021e022302290228021f0214020502f901f701f701f601f701f401ed01ea01e201d501d001cd01c901cb01cb01c501c001b901b401b501b501b501b801b601ae01a7019f0198019601940195019901950188017a016d01650167016f017d0191019b019501860171015a014c0147014b015b016c01760175016a01570146013a0135013c01490155015b0157014d01410135013101380143014a014d014a013d012b011e0118011c0124012d0133013101290122011d011c0121012601280126011c010e0104010101010106010f011801190111010601fc00f400f400fb000601100111010701f800e500d300cc00d200de00ec00f600f700ec00d900c600bc00ba00bd00c900d600dc00da00d200c500b800b000af00af00af00b100b100ab00a00095008c0088008b0091009600950091008c00860080007e007e007c00790076006d00620059005300500054005a005b0057004e00410035002c0028002f003a004000400037002a001e0012000b000c000e00120015000e000100f4ffe8ffdfffdeffe2ffe9ffeffff1ffedffe5ffd8ffc8ffbaffb0ffacffb0ffb4ffb5ffb4ffacffa2ff9aff95ff94ff98ff99ff96ff8fff86ff7aff6fff69ff67ff67ff65ff61ff59ff4dff45ff41ff3fff42ff47ff49ff45ff3cff2fff22ff19ff0fff0dff12ff13ff11ff11ff0afffdfeeffee3fedcfedcfedefee2fee4fedffed4fec7febafeb4feb6febcfec4fecafec6febcfeacfe97fe86fe7ffe7bfe7dfe85fe88fe87fe82fe77fe6efe67fe60fe5dfe5dfe57fe53fe52fe4bfe45fe41fe3bfe37fe35fe2ffe29fe26fe1ffe18fe14fe0ffe09fe09fe06fefffdf8fdeffdeafde8fde5fde5fde8fde5fdddfdd4fdc4fdb4fdabfda5fda6fdadfdb0fdb0fdaffda6fd98fd8dfd83fd7bfd7afd7afd7bfd7afd70fd63fd57fd48fd40fd40fd41fd47fd50fd4ffd47fd3efd2cfd1cfd14fd0dfd0dfd14fd14fd0ffd0afdfdfcf0fce8fce0fcdcfcdcfcd7fcd2fccefcc3fcbefcbffcbcfcbbfcbdfcb4fcabfca2fc92fc89fc8bfc8afc8cfc93fc8dfc7ffc72fc60fc50fc4efc4ffc54fc5cfc5dfc59fc53fc44fc37fc30fc27fc24fc27fc23fc20fc1efc12fc06fc00fcf7fbf5fbfafbf6fbf4fbf6fbedfbe1fbd7fbc9fbc3fbc5fbc0fbc1fbc7fbc3fbbefbbdfbaffba2fb9cfb93fb8dfb8cfb86fb86fb89fb82fb7efb7ffb77fb70fb6dfb60fb54fb4ffb46fb46fb4cfb49fb49fb4afb3cfb30fb2bfb1ffb17fb1cfb1cfb23fb2efb2afb21fb16fbfffaeefaebfae8faebfaf6faf8faf8faf6fae6fad9fad4faccfacdfad8fad8fad4fad2fac7fabefabdfab4fab5fac0fabefabafabafaaffaa5faa2fa9afa99fa9ffa9efaa1faa8faa3faa1faa3fa9bfa98fa9efa98fa93fa95fa8efa8bfa90fa8efa8ffa96fa95fa93fa93fa88fa82fa86fa86fa8dfa9afa9efaa1faa2fa95fa8bfa8afa83fa85fa93fa9afaa2faadfaadfaaafaa9faa2faa2faabfaacfab0fabafab9fabafac0fabefac2facdfacefad1fad8fad5fad3fad8fad7fadefaedfaf0faf6fa00fbfffafffa06fb08fb11fb1efb20fb23fb29fb27fb29fb32fb35fb3efb4bfb4ffb56fb5ffb5efb63fb70fb73fb7bfb8bfb91fb98fba1fba3fba7fbaefbabfbacfbb6fbc0fbcffbe0fbe8fbf2fbfdfbfbfbfafbfdfbfffb09fc19fc26fc35fc46fc4bfc4efc56fc58fc5dfc66fc6cfc75fc80fc84fc8dfc9bfca5fcb3fcc4fccafccefcd6fcdafce1fcebfceefcf8fc07fd0dfd12fd1bfd20fd27fd37fd45fd53fd62fd6afd71fd77fd79fd80fd8bfd92fd9cfda9fdb2fdbafdc4fdcafdd4fddffde5fdeffdfcfd04fe0cfe18fe22fe2dfe3afe42fe49fe50fe54fe59fe63fe6dfe79fe89fe94fe9afe9dfe9ffea5feb0febbfec7fed6fee4fef1fefcfefffe00ff06ff10ff1cff29ff32ff39ff40ff46ff4cff53ff5eff69ff71ff78ff80ff89ff90ff9affa7ffb2ffbaffc2ffc6ffc9ffceffd5ffddffe7fff4ff000008000e00120016001d0025002c0038004600500058005e00610066006a006c00760084008f009a00a300a500a400a500a900b100bb00c600d500e200eb00f200f400f200f400fa00ff0006010e0113011a0121012c013b01450148014c01510153015801610169017101780182018a018b018c01910193019601a101ac01b501c201ca01ca01ca01cb01cd01d501df01e801f601010204020802080204020802100219022602320236023a023a0239023d0242024902580265026d02760279027502770278027802800287028b0295029e02a002a602ab02ac02b102ba02c002c502c702ca02cf02d102d602e202eb02ed02ef02ee02ec02ed02ee02f40202030c0313031b031a0312031103110313031d032a033403400341033803350332032c0330033b0344034f035503520350034b034903500359035e0369036d036903680364035e0364036b036d03720372036d036d036e036f0377037c037d0383038203790377037603730377037e0380038603860381037f037b03750377037b03800388038a0383037f03790370036f03720374037e0386038403800379036c036503640365036c03730375037603710365035e035c035d0364036703640362035d0352034a034603440347034b034d0352035003470341033b033503350335033403360333032b0326032203200326032703240323031a030d030403fc02f902010308030d0313030e030203fb02f202e902eb02f002f202f502f302eb02e302d802cf02d002d102d202d902dd02d702d102cc02c402c302c402c302c602c702c202be02b602ad02ab02ab02ac02b202b702b602b402ab029e029a02990299029c029e029d029e029902930290028d028e02940292028d028e028b0282027d027b027b0283028702860285027f0275026f026b026c027202750277027b0276026d02690263025f02640269026d0272026f026602600257024e025002530254025a025d025902570253024d024c024d024c024b024a02480245023e0239023c023f0240024302450240023b0232022c022c022b0229022c022d02290224021e02170217021c0222022602260224022002130205020002fe01000209020f020f020a02ff01f601f001e901ea01f401fa01fb01f601ed01e201d601cc01cc01d301d801dc01de01d801cd01c301b901b501b601b501b401b401ad01a301a0019d0199019b019d019d019b01920186017c017401700170017101740175016d0163015c0152014c014d014c014a01480140013601310128011f011b011a011a011c011b0115010d010101f600ee00e700e500e600e500e000d900d100ca00c400bd00ba00ba00b600af00a7009c00920087007e007d007e007d007c0078006f00630057004f004b004800450043003b002f002300180010000f00110010000e000a000000f4ffe8ffdeffdaffdaffd6ffd3ffceffc3ffb6ffacffa5ffa2ffa2ffa1ff9fff9dff94ff88ff7dff72ff68ff61ff61ff61ff5eff5bff57ff4eff43ff3bff33ff2dff2cff2aff25ff21ff19ff0dff03fffefefffe00fffefefffefcfeeffee1fed7fecdfec9fec9fec7fec6fec4febcfeb5feb1fea9fea7feaafea7fea4fea3fe99fe8dfe87fe7ffe77fe76fe77fe77fe78fe75fe6efe69fe62fe5bfe59fe59fe58fe56fe50fe48fe40fe37fe32fe34fe37fe3afe3ffe3efe35fe2cfe22fe18fe14fe11fe11fe15fe16fe13fe0ffe08fe02fe01fe00fe02fe07fe07fe01fefafdf2fdeafde4fddffde3fdeafdecfdebfdeafde5fde0fdd9fdd2fdd3fdd8fdd6fdd5fdd6fdcefdc5fdc2fdc1fdc3fdc9fdcdfdcffdcefdc8fdc1fdbbfdb6fdb7fdbafdb9fdbcfdbefdb9fdb6fdb7fdb6fdb7fdbbfdbdfdbefdbefdb6fdaffdabfda7fda8fdb0fdb5fdb8fdbdfdbefdbdfdbbfdb8fdb6fdb7fdb7fdbafdbcfdb7fdb3fdb5fdb4fdb4fdb8fdbdfdc6fdcffdd0fdd0fdd0fdc9fdc4fdc7fdc8fdccfdd5fddbfddefde0fdddfddcfddcfdddfde6fdedfdeffdf4fdf8fdf4fdf2fdf3fdf3fdf8fd03fe0cfe14fe18fe16fe17fe1afe1bfe1ffe25fe29fe2ffe31fe2ffe32fe36fe3afe42fe4dfe56fe60fe65fe63fe63fe65fe63fe66fe70fe7afe84fe8efe91fe91fe94fe96fe9bfea6feaefeb5febdfebefebcfebffec2fec7fed1fedefeebfef5fef9fefdfe02ff02ff03ff0aff12ff1bff26ff2dff2fff33ff37ff3cff44ff51ff5eff6bff74ff7bff7dff7dff7dff80ff85ff8eff9affa7ffaeffb2ffb8ffc1ffc8ffd2ffe0ffeafff2fff8fff9fff9fff9fffdff0600130020002e0039003f004200450049004d00560062006c00730078007c00800086008f009a00a800b300bb00c000c000bf00c200c700cf00d900e200ec00f600fc00000106010d0114011e012a0131013301360138013801390140014a0155015e016701700173017401760178017b0183018e019401970198019a019e01a201a801b501c001c501c701c701c701c701c701c801cf01d901e001e601e901eb01ed01f101f701fc01fd01000203020102fe01fd01fc01fc0102020b0214021b021d021e021f021e021b021b021d021f02210223022302240221021e021d022102290231023302320231022c022702260228022b022f0230022f022e022b0227022802290228022902260222021e02190217021802180217021d0220021e021d021b02160212020d020b02090204020002ff01fa01f501f401f501f701f801f401f201f001e801df01dc01d801d401d401d201ce01cd01c901bf01b901b601b301b101af01ab01a601a1019a0193018c018501820180017f017f017e017b017301690160015a0153014c014b0147013f01380134012f012d012f012e01290122011a0110010701ff00f700ee00e900e600e200e100df00da00d500d200ce00c900c300ba00b300ad00a5009f009a0093008c008a00880084007e0075006d00650060005d005b00590057005100490041003b003800360033002d00270021001a0013000c000500fffffafff8fff6fff2fff1ffefffebffe9ffe7ffe1ffd8ffd0ffc9ffc5ffc0ffbaffb7ffb4ffafffadffabffa6ffa1ffa0ff9bff96ff93ff8fff89ff86ff82ff7cff77ff76ff74ff71ff6dff6aff67ff63ff5cff58ff54ff51ff4eff4aff44ff40ff3cff3aff3bff3bff3aff38ff31ff27ff23ff21ff1fff1cff1aff19ff16ff0fff0bff0aff08ff09ff0bff0cff0aff06ff00fffcfef7feeffeebfeecfeeefeeffeeffeecfee9fee7fee5fee5fee2fedefedffee0fedffedcfed8fed4fed3fed5fed6fed7fed7fed5fed4fed2fecdfecafecbfeccfecbfecbfec8fec7fec9fecafec9fecbfecefecffecffecefecefecbfec5fec6fec8fec5fec6fecbfecbfecafecbfecafecafec9fec8fecffed6fed5fed4fed4fecffeccfec9fec8fecdfed4fed6fed8fedafed7fed5fed3fed1fed2fed5fed7fed9fedcfedbfedbfedafed5fed6feddfee1fee2fee2fedffedcfedbfed7fed6fedbfee1fee7feeafee6fee2fee3fee3fee3fee4fee6feeafeebfee5fee2fee2fedffeddfee1fee5fee7fee9fee9fee9fee6fee2fee2fee4fee3fee6feebfeeafee9fee8fee2fee0fee3fee5fee7fee9feeafee9fee4fedffedefedffedefee3fee9feeafee9fee7fee3fee1fee3fee3fee3fee2fee4fee5fee3fedffedefedffedffee0fee3fee4fee3fee3fee3fee3fee1fedffee3fee7fee8fee9fee9fee5fee1fedffee0fee4fee8feebfeeefeedfee9fee9feecfeebfeeafeecfeeefef0feeffeeffef1feeffeebfeedfef0fef0fef5fefafef9fef9fef8fef5fef3fef5fef9fe00ff06ff06ff06ff05ff00fffbfefbfefffe05ff08ff09ff09ff08ff06ff06ff06ff09ff10ff15ff13ff12ff14ff14ff13ff13ff13ff14ff17ff18ff18ff18ff15ff15ff14ff13ff17ff1fff22ff23ff23ff20ff1dff1dff1dff1fff22ff27ff2cff2bff25ff22ff20ff1fff22ff28ff2bff2dff2fff2bff29ff2aff2aff2aff2fff31ff33ff37ff37ff34ff34ff35ff34ff35ff36ff37ff3aff3dff3bff39ff39ff3aff3cff41ff46ff48ff4aff4bff46ff41ff42ff45ff48ff4dff53ff53ff51ff51ff52ff53ff55ff58ff5bff5fff64ff64ff63ff66ff68ff66ff67ff6cff6fff70ff73ff74ff72ff73ff76ff77ff79ff7eff83ff8aff8eff8cff8bff8cff8cff90ff98ff9cff9effa0ffa2ff9fff9cff9effa3ffa8ffacffb1ffb3ffb4ffb6ffb8ffbcffc2ffc7ffc9ffcdffcfffcfffcfffd1ffd3ffd8ffdcffe0ffe4ffe7ffeaffebffebffedfff0fff2fff8ff0100060009000a0009000a000d00130018001d002200270028002600280028002a00300038003e004300470049004b004d005000550059005e006400670068006a006e007100730076007b00830089008e009300970098009b009d009e00a300aa00ae00b000b200b400b800be00c100c700ce00d100d500da00dc00dd00e100e900f100f500f900fe0000010201060109010c011201160119011e012101240129012d0132013b01430149014e0150015101540152015201560159015f0168016d0172017801780176017c0185018b018f0192019501980199019b01a001a401a701ad01b201b401b801bb01bc01c101c601c801cc01d001d201d601d801d901de01e201e401eb01ef01ef01f201f301f201f501f801f901fd01020206020a020a020a020e021002120219021c021b021d021d021d021f021f021d022002230227022b022b022c02300231022e022e0230023302360238023802380237023402350237023b023e023e023c023d023b0237023602370238023d0240023d023d023e023d023c023a0238023b023b023502320230022d022c022b022b0230023102320232022d02270226022402220224022302220223021f021602120210020f020f020e020d020d0208020202ff01fd01fb01fb01f901f701f601f201ed01e801e301df01de01db01d801d701d201ce01cd01c801c301c101bf01bd01be01bb01b501b101ab01a501a1019a019601970193018c01880181017a017a017b017a017a01750170016c0160015601550152014b014901450140013c0133012d012c012701240125012101190115010e0106010201fe00fc00fa00f500ee00e900e200da00d300ce00ca00c600c100bc00b800b100a800a2009f009f009d009a0095008d00850080007a00740070006b0064005e0056004c00460043003e003b003900350030002a0023001e0017000f000d000b0007000300fbfff2ffecffe5ffdcffd6ffd1ffceffcdffc9ffc2ffbeffb9ffafffaaffa8ffa2ff9dff9aff94ff8eff88ff80ff7aff75ff70ff6bff66ff5fff5aff56ff51ff4fff4cff47ff42ff39ff32ff2fff29ff21ff1cff18ff13ff12ff0fff0aff04fffefefafef7fef0feeafee8fee3feddfed7fed2fecffec9fec1febefebdfeb7feb3feb1feacfea7fea2fe9bfe96fe96fe93fe8efe8bfe86fe81fe7efe78fe74fe73fe6ffe69fe68fe63fe5dfe5afe57fe50fe4bfe49fe48fe46fe43fe42fe43fe3efe38fe35fe31fe2dfe2bfe26fe23fe23fe1ffe1bfe1bfe16fe12fe12fe0efe0bfe0cfe07fe04fe05fe06fe07fe05fe00fefdfdfbfdf5fdf4fdf4fdf1fdf0fdeffdeafde9fde9fde4fde4fde6fde1fddffde4fde3fde0fde1fde2fde2fde3fde1fddefddefdddfdddfdddfddafdd8fdd7fdd6fdd6fdd6fdd6fdd9fddcfddafddafddefddafdd7fddbfddbfdd9fddafdd9fddafddefddefddcfddefdddfdddfde1fde0fde1fde6fde5fde6fdeafde8fde9fdeefdeefdf1fdf6fdf3fdf3fdf9fdf8fdf8fdfdfdfcfdfcfd01fe01fe04fe0afe0bfe0dfe12fe14fe17fe1afe18fe19fe1cfe1efe22fe26fe25fe26fe2bfe2ffe35fe3cfe3ffe41fe46fe48fe4afe50fe54fe59fe5efe5ffe64fe69fe68fe68fe6cfe6ffe76fe7ffe80fe84fe89fe89fe8efe99fe9cfea1fea9fea9feaefeb9febafebbfec2fec6fecbfed3fed5fedbfee1fee0fee4feeffef1fef4fefefe04ff09ff11ff16ff1bff21ff24ff2bff31ff35ff39ff3eff40ff42ff49ff50ff56ff5cff62ff69ff6eff73ff7aff7fff84ff8bff91ff95ff98ff9dffa3ffa8ffaeffb3ffb9ffbcffc1ffc8ffceffd0ffd4ffd8ffdbffe1ffe7ffecfff4fffbfffdff030009000b000f0016001a001e002300230025002b00300035003a003d0043004b005000530057005b0060006300620065006b006e00700076007c007f00800085008a008f00930097009a009b009c009f00a300a700a900ad00b200b600b900bc00bf00c100c500c900cb00cc00cf00d200d500da00de00e000e300e600e800ec00ef00f000f100f300f300f400f700fb00ff00010105010a010c010b010d0110011101140118011a011c012001220123012501240125012901290129012d012f012e01310135013601360139013b013c013d013f0141014301450148014601450148014a0148014801480149014c014f014f01500151014f01510152015101540156015501550156015401520152015301550156015601550151014f01500150014f01500151015101530151014c014a014b014a014901470146014701470144014301430141013e013c013b013a0138013401310130012e012d012c01290128012801240120011e011c011b011b01190117011501110110010e010a0109010901050102010001fc00fb00fa00f600f600f400ef00ed00eb00e700e600e300df00de00da00d500d500d500d200d100ce00cb00ca00c700c500c300bf00bc00bc00b700b200b100b100af00b000af00ac00aa00a600a2009e009a0099009a009a009700960093008e008d008c008700850082007f00800080007a00780077007400740074006f006e006d006900660062005c005d005e005a0058005700550053004d004a004b004a004700460043003f003d003900360035003300320030002e002d002c002a002b0029002400210021001e001b0016001300150014001000100010000d000c000a000700030002000100ffffffff00000000fdfffbfff8fff6fff6fff7fff7fff5fff4fff5fff1ffebffebffecffe9ffe6ffe6ffe9ffecffebffebffedffecffe8ffe7ffe9ffe9ffe8ffe8ffe7ffe4ffe1ffe1ffe0ffe0ffe4ffe5ffe4ffe6ffe5ffe0ffe2ffe6ffe6ffe9ffebffecffedffebffe6ffe6ffebffebffe8ffe9ffedffefffeeffefffefffeefff1fff3fff3fff4fff4fff3fff5fff8fffafff8fff7fff8fffafffcfffefffffffdfffeff0000020004000600060005000500060009000c000c000a000e00130013001100120012000f0011001300120015001900190019001b001d001f0020001f00200022002400230023002300240023002400280029002a002e0030002c002b002c002c002e003200330034003600340033003300320033003800390037003700380037003600370039003b003c003e003e003c003d003e003d003f0042004100400040003f00400041003f0040004400460047004700470049004a00480046004600460049004900450044004500430044004a004d004c004c004b004b004d004e004c004c004c004c004c004d004e004d004a004b004c004c004d004a0048004a004c004b004c004c0049004a004b004b004b004a0048004600440044004600460047004900480047004600440042004100410041004100400040004100420041003e003c003c003c003b003a00380038003800370036003700360033003200340032002d002d0030002e002b002b00290028002900290029002800250023002500250021001f00200020002000210020001a00170017001500140014001200110012001400150012000f000f000e000f000f000c000b000c000800060005000000fdfffefffafff8fffbfffafff7fff7fff7fff8fff6fff2fff3fff5fff2ffefffeeffedffecffe9ffe4ffe3ffe3ffe1ffdeffdbffd8ffd7ffd6ffd5ffd2ffceffd0ffd2ffd2ffcfffccffcaffc8ffc6ffc3ffc2ffc0ffbbffb6ffb6ffb5ffb0ffadffaeffadffaaffa9ffa6ffa4ffa5ffa4ffa1ffa1ffa1ff9fff9eff99ff93ff91ff90ff91ff92ff90ff8cff8aff88ff86ff83ff81ff80ff7fff7dff7cff7cff7bff7aff79ff7aff7aff76ff74ff74ff71ff6fff6fff6bff69ff6bff6aff69ff6aff68ff66ff65ff63ff64ff67ff69ff68ff65ff65ff65ff63ff5fff5dff5cff5cff5cff5aff5aff5cff5dff5cff5bff5cff5dff5fff61ff61ff5fff5eff5fff5eff5eff60ff5eff58ff58ff5cff5eff5eff5cff5aff5cff5eff5dff5dff5fff5fff5fff61ff61ff60ff61ff61ff5fff5eff5dff5cff5dff5eff5fff61ff61ff60ff60ff60ff62ff65ff63ff60ff62ff64ff65ff65ff66ff65ff63ff62ff65ff67ff65ff65ff68ff6cff6eff6eff6dff6eff6dff6cff70ff71ff6fff70ff74ff74ff76ff76ff74ff76ff7cff7dff7bff7cff7eff80ff82ff83ff86ff8aff8aff8aff8eff91ff8fff8fff93ff94ff93ff94ff95ff98ff9cffa0ffa4ffa7ffa8ffaaffadffafffafffb1ffb5ffb9ffbaffbbffbbffbcffbdffc0ffc4ffc7ffc9ffceffd3ffd6ffdaffdbffdbffdeffe0ffe2ffe5ffe6ffe5ffe8ffecffedffeffff4fff8fffafffdfffeffffff00000300050007000a000e00110013001300150018001b001c001c001d001d001e001e001f00220026002a002b002a002b002f0030003200360037003600340033003200350039003800350038003d003e003e003d003d00400040003e003e003e003c003d004100430043004300450045004400440042003e004000430040003f0040003f0041004300420045004a004a00470045004200410041003f003e003f004000410040003f003e003d003d00410044004500430040003f003e004000420043004400450046004700470045004500460044004300430041004000400040004400470048004b004d004e0050004e004a004c004e004d004d004d004d004f0050004f005000520051005100530053005400560055005300540055005500560057005600570056005500540053005200550055005300530052005300560057005900590057005700580053004f004d004c004d0050004e004e004e004a00480049004700450044004300430040003b0039003a003a003a0038003600390039003600340031002f0030002d002600240022001d001b001a00180019001b001b001a001900150010000c00070006000800060003000300030001000000fdfffbfffcfffcfffcfffcfff8fff4fff0ffecffecffecffebffeaffeaffe7ffe5ffe5ffe7ffeaffebffe9ffe9ffe7ffe3ffe2ffdeffd6ffd6ffd8ffdaffddffe0ffddffdcffdeffdeffddffdbffd8ffd8ffdaffd8ffd6ffd4ffd2ffd2ffd8ffdcffd9ffd6ffd6ffd5ffd4ffd4ffd4ffd4ffd5ffd4ffd5ffd3ffceffcdffd1ffd3ffd3ffd3ffd4ffd6ffd6ffd3ffd2ffd3ffd1ffd0ffd0ffceffceffceffceffcfffceffccffccffceffcdffcbffc9ffc7ffc6ffc6ffc4ffc2ffc2ffc4ffc5ffc6ffc7ffc7ffc7ffc5ffc2ffc2ffc2ffc2ffc2ffc2ffc2ffbfffbbffb9ffb5ffb1ffb0ffb1ffb0ffb1ffb4ffb5ffb7ffb6ffb4ffb5ffb5ffb4ffb4ffb4ffb1ffb0ffb1ffb0ffb1ffb2ffafffabffaaffa9ffa7ffa6ffa6ffa8ffaaffaaffaaffacffabffaaffaaffaaffa9ffaaffabffabffaaffaaffacffacffacffb0ffb3ffb2ffb1ffb3ffb3ffb3ffb3ffb2ffb3ffb2ffb0ffb1ffb1ffafffb1ffb4ffb3ffb3ffb6ffb8ffbaffbcffbeffc0ffc2ffc1ffc3ffc4ffc2ffc3ffc9ffccffcbffcbffcdffccffcaffc8ffc8ffc9ffcaffcdffd3ffd6ffd6ffd9ffdbffdbffdcffdcffdbffdcffdaffdaffdeffdeffdfffe4ffe7ffe8ffedffedffe9ffeaffeaffe8ffe9ffe9ffeaffeefff0ffeffff0fff1fff1fff3fff4fff4fff3fff3fff4fff5fff5fff7fff8fff8fffafffdfffcfffbfffcfffdfffbfffcfffdfffefffdfffcfffcfffefffffffdffffff03000600080008000700070006000300030005000600090008000700080006000000ffff000002000600070008000c00100013001500120011001200100010000f000c000d001000110015001b001b001b001e001e001e0020001d001b001c001c001c001d001e001e001f00200022002200240028002c00300032003200340038003b003a003b003e003f003d003c003b003d003f003e003e00420043004100420042004300470049004d0053005600570059005a005a005b005c005e005f005d005b005d005f00620064006300640068006a0069006700660065006400650068006800680069006b006d007000720077007a007800760077007400720071006f006f00700072007400760076007700770076007600760074007300740074007400730072007400740071007000730074007100710073007300740074007100700070007000700071006f006d006c006c006b006b006b00690069006a00690069006c006e006c006d006f0070006f006d006900680068006600660064005f005e0060006100610062006400660067006600660066006600650065006600670068006a006a00680067006500620061005f005c005d006000600060005f005d005c005d005f0060005f005e005f006300640060005f005f005e005c005d005f00610062006400660066006500650063005e005a00570053004f004d004d004e005000520056005a005c005e00610061005f005c005b005900550050004d004c004b004a004a0049004a004d004c004c0050005300510050004d004a00470043004000400040003e003c003c003d003a0038003700340034003800380037003a003900330030002d0029002900290029002b002d002e002e002c00270021001d001c001b00180018001a001a001a001a001800150011000c000800060004000300050006000500040006000700070006000500060004000100fffffbfffafffafff8fff5fff6fff4fff0fff1ffefffe9ffe7ffe5ffe4ffe6ffe8ffe9ffebffedffecffecffebffe9ffe6ffe1ffdfffdeffdbffdaffdaffd8ffd8ffdaffd9ffd9ffdcffdcffdcffdcffd8ffd4ffd1ffcdffcaffc9ffcaffccffcdffcfffd2ffd3ffd3ffd1ffcfffcbffc9ffc8ffc7ffc7ffc7ffc7ffc5ffc5ffc3ffc1ffc0ffc0ffbfffc1ffc3ffc4ffc3ffc1ffbfffbcffb8ffb6ffb6ffb5ffb7ffb8ffb8ffbcffbfffbcffbbffbcffb9ffb6ffb5ffb2ffafffaeffacffaaffa8ffa8ffaaffacffaeffb2ffb3ffb2ffb3ffb2ffafffb0ffadffaaffabffabffa9ffaaffaaffa6ffa4ffa2ffa0ff9eff9cff9aff99ff99ff9aff99ff9aff9dffa1ffa3ffa5ffa7ffa7ffa6ffa4ffa2ffa0ff9dff9aff99ff99ff9aff9bff9dff9fff9dff98ff95ff93ff91ff8fff8eff8fff91ff94ff97ff97ff95ff95ff94ff93ff96ff98ff99ff9effa1ffa1ffa1ffa1ff9eff9bff9aff97ff97ff9aff9dff9eff9eff9fff9eff9bff99ff96ff94ff94ff94ff93ff97ff9bff9effa3ffa9ffafffb4ffb9ffbcffbeffbfffbdffb7ffafffaaffa6ffa4ffa3ffa5ffabffb0ffb6ffbdffc2ffc6ffc8ffc9ffc8ffc6ffc2ffc0ffc0ffc0ffc1ffc5ffcaffceffd4ffdaffddffdfffdfffdfffdcffd6ffd1ffceffcaffc6ffc8ffcfffd7ffdeffe3ffe7ffecfff0fff1fff2fff2fff0ffefffefffedffeaffe8ffe6ffe5ffe8ffecfff0fff6fffafffcfffcfff9fff3ffebffe4ffe0ffdeffdfffe4ffecfff6ffffff05000c00110011000d0008000100fafff6fff3fff2fff3fff5fffaff010005000600070006000100fcfff8fff3fff1fff0fff2fff5fffcff030009000f00150018001b001e001c00180014000f000a0007000300fdfffcfffeff010006000f00190023002b002f002f002d0025001c0014000e0009000a000d0013001b0023002b003100350036003500320030002f002e002f0034003a004100460049004a0047003f0036002d0024001d001b001e0024002f003e0050005f006a007100730072006d00630058004c0042003b0036003300350038003c0044004d00560060006a0072007b0080007f007e007b00720067005d0054004e004a0048004b00520057005c00610064006500630060005f00600064006a0072007c0087008f00930093008e0083007500640051004100370033003900470058006d00830092009b009c00930085007400630058005300510054005b0062006b00720074007500730070006e006c006a006c006f007100730072006e006900610059005300520054005b0063006c0075007900780074006e0067005f00580054005300540056005c006200660069006a0066005e0056004d00470048004f005b006a00790085008900840076005f00430029001400080007001100240040005c0076008c009a009c00960087006f0054003a00230013000a0008000d0014001d0028003100380040004900510058005c005d0058004f00430037002b002000190017001400120010000e000a0006000100fbfff4ffeeffecfff1fffaff0b002500400059006b006f00630047001e00eeffbeff95ff78ff6dff70ff82ffa0ffc4ffe9ff090021002d002d0022000e00f7ffdfffccffc0ffbaffbbffbfffc1ffc1ffbbffafffa1ff91ff84ff7fff80ff88ff95ffa6ffb7ffc5ffcfffd1ffceffc6ffbaffabff9dff8fff84ff7bff74ff70ff6eff6bff67ff64ff61ff61ff66ff71ff81ff95ffaaffbbffc3ffbeffaeff92ff6eff49ff29ff12ff09ff0dff1fff3aff5bff7bff95ffa5ffa8ff9dff85ff64ff41ff23ff0fff07ff0eff22ff3eff5bff72ff80ff82ff76ff62ff4bff32ff1cff0fff0aff0dff15ff1fff2bff36ff3cff3bff37ff31ff2aff26ff25ff2aff33ff3dff47ff4eff4bff40ff30ff1cff06fff3fee5fedefedffee8fef5fe03ff10ff18ff1dff20ff1eff1cff1bff1cff22ff2eff3aff46ff50ff52ff4aff38ff1cfff7fed1feb0fe98fe90fe98feaffed1fef8fe1dff3bff4eff54ff50ff45ff39ff30ff2eff34ff40ff4bff51ff4cff3aff1affeffebffe92fe73fe67fe73fe98fecffe13ff59ff96ffc2ffd8ffd4ffbcff94ff63ff31ff08ffe8fed2fecafecbfed1fedcfee8fef4fe03ff15ff2aff42ff5dff79ff93ffa7ffb1ffaeff9fff84ff61ff3aff17fffdfeeefeeefefcfe14ff32ff50ff68ff78ff7eff7aff71ff68ff62ff64ff6eff7fff95ffabffbbffc3ffbfffadff92ff70ff4dff2fff1aff12ff18ff2cff4bff72ff9bffc2ffe3fffcff080009000000edffd4ffb9ffa0ff8bff7fff7bff7fff8bff9cffafffc2ffd0ffdaffe0ffe1ffddffd7ffd0ffc9ffc5ffc3ffc5ffccffd9ffeaff02001d003b0058006f007c007c006a0049001c00e7ffb5ff8dff76ff76ff8fffbcfff8ff380073009f00b600b700a3008000590037002200210036005c008d00be00e200f300e900c5008a004200f9ffbdff96ff8effa7ffdeff2c008700e0002f016b018c0192017f0159012501ec00b3007d004f002b0011000100fdff06001d0040007200af00f3003a017a01ae01d001d801c401960155010701b80071003b001c0017002b0052008600bf00f50020013e014e0153015201500150015701640174018201870181016a0144011301dd00aa0082006900640074009500c500fd0037016d019b01bd01d301dc01db01d201c001a8018901630137010701d700ab008b007b0080009d00cf0011015b01a501e4011102260221020402d40198015a012201f600da00cf00d400e400fc001601300149015f01740188019a01ab01b901c101c101b701a40187016501430124010f0106010a01190130014901600171017a017a0172016501560147013b013201300135014001500163017701880196019e01a0019b01910181016e0155013a011c01ff00e500d100c400bf00c300cd00dd00f000070121013d015c017c019901b101c101c601bf01ac018f016b0140011101e000ae007d0051002c0012000500090020004a008600d20027017e01ce010e02320236021502d3017401040190002500cfff97ff82ff8fffbafffaff46009200d50009012a013801340123010a01ec00cc00ae0092007900630050003e002d001f0013000c000c001500280045006a009200b900db00f30000010001f100d400a9006f002800d8ff87ff3bfffefedafed5fef1fe2fff8afff9ff7200e9005201a201d001d401ae015f01f0006c00e3ff64fffbfeb3fe8efe8efeacfee2fe26ff6fffb6fff2ff1e00390043003e00310024001b001c0029003f0058006d0076006d0050001e00dbff91ff47ff07ffd9fec2fec4feddfe08ff3dff74ffa4ffc7ffd8ffd5ffc3ffa5ff83ff66ff54ff56ff6cff97ffd0ff0f0049007200840077004d000900b0ff4effeafe8efe45fe14fe02fe0ffe3afe7efed2fe2bff80ffc7fffbff1900220019000300e4ffc2ffa0ff84ff70ff65ff64ff6aff73ff78ff74ff62ff41ff13ffdcfea5fe76fe55fe49fe52fe71fea2fee1fe28ff71ffb4ffebff0f001a000b00e4ffacff6bff2efffefee5fee6fe02ff35ff75ffb7fff0ff12001500f2ffaaff42ffc6fe42fecafd6cfd37fd34fd67fdcefd60fe0fffc8ff78000c017301a4019a015901e8005600b4ff12ff82fe11fecafdb0fdc2fdf9fd49fea3fef9fe3eff6cff7fff7cff68ff4cff2eff14ff04ff01ff0cff27ff50ff84ffbdfff4ff2200400049003d001f00f1ffb9ff7dff3fff05ffd2fea7fe87fe74fe6efe75fe84fe99feb0fec5fed7fee8fefafe0fff2cff51ff7effb4ffeeff2b0067009d00c900e700ef00dd00ae005f00f3ff6fffdcfe43feb0fd31fdd0fc98fc91fcbffc23fdb7fd74fe4bff2c000401bf014b029902a3026702eb013d016f0096ffc8fe18fe94fd46fd31fd52fd9ffd0afe82fef5fe52ff8fffa5ff98ff71ff3cff0dfff1fef8fe27ff7ffff8ff83000e018401d101e601ba014c01a500d6fff7fe21fe70fdf8fcc9fce7fc49fde1fd95fe4efff2ff6f00b800cb00ab00630003009cff43ff08fff6fe15ff62ffd4ff5900dd004a018c0197016601fb006300adfff0fe42feb7fd60fd45fd69fdc4fd49fee4fe7fff08006f00ad00bf00ad00820049001100e6ffd1ffd7fff7ff2d007100b600f2001b0128011501e0008d002000a1ff18ff90fe13feadfd65fd44fd4efd86fde9fd75fe21ffe4ffb00076012802b4020d032a030603a202070243016a0090ffcbfe2bfebdfd86fd86fdb4fd08fe73fee7fe54ffaeffecff0b000d00fcffe5ffd7ffe0ff09005400bd003901b70123026a027c024e02db012901450045ff46fe63fdb8fc5afc54fca7fc4bfd2dfe34ff41003801fd017c02ab02890220028301cb00120074ff04ffd2fee4fe34ffb4ff4e00e7006101a501a0014c01ae00d8ffe4fef1fd22fd94fc5dfc89fc19fdfffd25ff6a00a801bc028503ed03e8037b03b702b7019e008fffaafe07feb7fdbafd08fe8ffe34ffdbff6700c400e100bc005a00cbff26ff85fe04febbfdb9fd07fea0fe75ff6e0070015c0216038703a1035d03bf02d801c00099ff85fea6fd19fdebfc20fdabfd74fe5bff3b00f200660188015701de0035007bffd2fe57fe1ffe38fe9efe45ff1800f900cc017702e4020a03e3027702d2010601290051ff91fef9fd96fd6efd82fdcdfd45fedcfe81ff2200ae0015014f0158013501f1009b0046000200ddffddff03004800a000fc004b017d0185015901fa006f00c7ff17ff77fefdfdb7fdaefde0fd46fed2fe76ff2200c9006001de013f027f029b029102600208028a01ec00350073ffb4fe0afe86fd39fd2ffd6efdf3fdb2fe96ff83005b0100025e026a022902a90104015b00cdff75ff63ff99ff0e00aa005101e2013d024b02fd0153015c0035ff06fefbfc3ffcf3fb2afce4fc0dfe83ff17019702d203a304f004b004eb03bc024901c0ff54fe33fd81fc54fcb0fc87fdbafe1f008601c102a7031e04170492039e025901e8ff7afe3dfd5efcfcfb29fce1fc0bfe7dff020160026403ec03e8035c0362022301d0ff9efebafd49fd5dfdf6fdfffe5300c30118031f04af04ad041104e802540184ffb3fd1dfcf5fa63fa79fa35fb7ffc2ffe1300f2019403cd047a058f050d050d04b2022b01a7ff55fe5bfdd3fcc8fc37fd0cfe25ff5a007b015d02dd02e402700292016e0036ff1ffe5bfd0ffd49fd01fe1aff6600b101c6027f03c0038503d902d601a20066ff49fe6efdeefcd3fc1efdc2fda7feafffba00ab016b02ed022b032903ee028302f5014f019d00eaff41ffaefe39feeafdc7fdd0fd07fe67fee7fe7dff1700a600190164018201750147010801c7009400770074008800ab00d400f8000d010b01ec00af005700ecff79ff0affabfe66fe43fe47fe75fecdfe4dffecff9f005301f6017202b602b7027102e80125013b0040ff4dfe7afde2fc99fcb0fc2efd0efe40ffa400110258034d04ce04c70438043403da015800dcfe94fda8fc31fc3afcbafc98fdadfecbffc6007b01d501ce017301dc002b0083ff02ffc0fec6fe14ff9dff4e000d01c1015002a902c002920224028301c000eeff20ff68fed7fd7bfd5dfd83fde9fd85fe45ff1200d2006c01cf01ed01c5015f01cd00280089ff0cffc4febdfef8fe6afffeff9a0023018201a90195014e01e2006500ebff85ff40ff26ff38ff74ffcfff37009700dc00f400da008f002000a0ff23ffbcfe77fe5bfe65fe90fed4fe29ff89fff1ff5e00ce003d01a501ff014202680269024302f3017a01dd00270065ffabfe0dfe9afd60fd63fd9ffd0cfe9cfe3effe2ff7800f3004b017e018d017b014e010d01bf0068001100beff78ff43ff25ff23ff3dff71ffbaff0f006300ac00de00f300e700bf0080003700eeffb1ff89ff7eff8fffb7ffebff1d003e0044002a00f3ffaaff5cff15ffe1fec4febefecffef4fe2dff79ffdaff4c00c6003d019f01e001f501de01a1014b01e80083002200caff7bff37ff00ffdafec8feccfee4fe0dff3eff70ff98ffafffb1ff9dff78ff4bff22ff0bff11ff40ff9bff2200cc0086013a02cc0223032a03d90231024201290006fffffd39fdcefccdfc36fdf7fdf5fe0a000f01e20166028d025202be01e700ecfff1fe1cfe89fd4afd63fdc9fd67fe24ffeaffa7005101e3015902b102e402e802b6024902a701e0000c0046ffa7fe41fe18fe27fe61feb5fe10ff65ffa9ffd7ffecffe7ffceffa9ff85ff6eff73ff9efff1ff6800f600860105025c027d025e02fe0162019800b4ffd1fe0cfe81fd49fd6ffdf6fdccfed8fff300f801c00232033f03e70237024901390028ff30fe66fddafc93fc97fce5fc79fd4afe48ff5e007001640220039003ac037303f10238025e017c00a7fff1fe6bfe1ffe13fe4bfebdfe59ff0600a50019014c013401d700440094ffe2fe47fed8fda5fdb8fd15feb6fe90ff8c008e017602250380037a0310034f025001320019ff27fe75fd16fd15fd72fd25fe1bff3a005e015f021603650337038d0278011b00a3fe45fd2ffc89fb68fbd3fbbcfc07fe8bff17017c028c0327043c04ca03e702b501620021ff20fe84fd60fdb7fd74fe73ff86007a0125026a023b02a101b1008cff57fe3bfd5dfcdcfbcffb40fc27fd6dfeeeff7701d802e3037804870414042f03f301840007ffa4fd81fcc1fb82fbd4fbb2fc04fe9cff3f01ae02b503310419047b0377023501e3ffaafeaefd07fdc3fce2fc54fd01fec6fe81ff1100630070004000e5ff7bff20ffedfef4fe3affbbff69002d01f0019802100346032f03ca021b022e011800f0fed1fdd3fc0efc91fb69fb97fb17fcdcfcd4fdecfe0d0024011d02e5026a039e037703f1021602fa00bfff8efe8ffde4fca2fccdfc58fd2dfe2bff33002601ec016e029e027502f701330144004bff6afebefd57fd34fd4bfd8afde0fd3ffea0fe01ff64ffc9ff2e008e00e30026015101620158013201f2009a002f00baff47ffe7fea8fe94feadfee9fe39ff87ffc1ffdcffd4ffadff73ff37ff09fff6fe07ff3cff8effecff43007d008b0064000a008bfff9fe6bfef9fdb6fdb0fdeffd72fe2fff12000201de018602dc02cd02550280016d0044ff30fe5afddcfcc2fc07fd9bfd66fe4cff3100f9008901cd01b6014001770072ff58fe50fd85fc14fc12fc83fc5dfd8afeecff5e01b702cd037c04a60443045b030f028e000fffc7fdddfc64fc5cfcb1fc44fdf2fd9bfe27ff86ffb4ffb4ff92ff5fff2cff0dff13ff47ffacff3700d7007401f20138023502e4014c018200a1ffcdfe26fec7fdbdfd06fe92fe43fff5ff8a00ea000a01ee009d0028009cff09ff7ffe10fecdfdc4fdfefd78fe24ffeaffaf005901d40116021b02e6017f01f1004a009cfffafe7cfe31fe22fe4dfea5fe12ff80ffdbff1c0044005b006a007700810085007d00670045001e00faffdeffccffbdffa9ff87ff54ff13ffcefe95fe78fe85fec5fe37ffd1ff81003101c7012d0254023702de015701b9001b0090ff26ffe2fec1febffed2fef4fe1eff4eff81ffb6ffedff25005a008900af00c600cc00bc00950059000d00b9ff6cff32ff18ff27ff5fffbaff2c00a50016017301b501d901db01bc017d012101b1003700c3ff61ff17ffe4fec3feaafe94fe80fe76fe81feaefe04ff83ff2300d300810118028702bf02ba02790203026a01c3002500a6ff56ff39ff4bff81ffc8ff0b00390048003100f8ffaaff57ff13fff3fe06ff52ffd4ff7c003301dc015a02970289023202a001e70023006effe0fe8bfe7bfeb3fe2cffd5ff93004701cf0114020902b20126018400eeff83ff52ff61ffa4ff09007a00e30035016601720157011801bb004a00d4ff69ff1cfffbfe0aff47ffa8ff1e009b0014018101dc01210249024e022902d9016501d8004200b5ff3effe8feb7feb1fed6fe27ff9fff3400d5006d01e10120021c02d8015d01c200210093ff31ff0aff25ff7dff0400a1003601a901e601e801b50160010001a800650038001a000000e3ffc3ffa5ff93ff97ffb5ffeaff2c006e00a600cc00e000e300dc00cf00bf00b100a500a100a900bc00d700f100fa00e400a7004200c2ff3cffc8fe7efe6efe9efe0fffb4ff80005d013102df024f03690325038702a201940080ff8afecdfd59fd35fd5afdbdfd4bfef0fe9aff3900c1002d018101c001f2011a023802440235020302ac013601ad002400aaff49ff02ffcffea7fe83fe63fe4bfe47fe60fe9afef5fe69ffeaff6d00e9005a01be0110024b02650256021602a30106014d008effe2fe5afe06feeafd04fe4cfeb5fe32ffb3ff2b008c00cf00ef00f200e100ca00b900b400b800b900a6006f000c0080ffdffe44fed0fd9dfdbcfd2ffee7fecbffbb009301370292029a025302ce0123016c00bfff2effc0fe76fe50fe4afe61fe8efecafe06ff34ff4bff48ff33ff20ff24ff54ffb8ff4a00f600a001270271026d0219027e01b100cbffe7fe1ffe85fd27fd08fd26fd75fde7fd6bfef3fe77fff2ff6600d60040019f01e4010102e6018b01f60037006cffb2fe26fed8fdcbfdf4fd40fe98fee8fe24ff45ff4dff42ff2bff0efff6feecfefdfe34ff9bff3300f600d001a6025303b303a403130300027f00bbfeedfc57fb30faa1f9b7f965fa89fbf5fc78feeaff3001390200038103bd03b5036c03e802350263018300a3ffd1fe17fe7efd10fdd6fcd5fc0dfd75fdfcfd8bfe11ff82ffdcff230060009500c000d700d100a80061000700b0ff6fff52ff5cff85ffbbffe9fffbffe7ffb0ff65ff1bffe9fee3fe0cff5dffc3ff240067007c005f001600b3ff4bfff2feb5fe99fe9bfeb3fedcfe12ff57ffafff1b00970015018201c701d00192010c014b0066ff78fea1fdfefca8fcadfc14fdd3fdd3feeffffe00d501570279024202d0014301be0055000f00e1ffb9ff86ff3bffd9fe68fefafd9ffd67fd5bfd7ffdd5fd5afe0bffdfffc800ae017402fa022303e00235023c01200017ff52fef6fd11fe96fe60ff3d00f5005d015701e300130011ff0efe3bfdc1fcb6fc20fdedfd00ff300050013902cc02f802bd022d0263018300afff02ff8ffe5bfe64fea3fe10ffa2ff51000d01c201510299027c02e601de0081ff04fea9fcacfb3afb61fb15fc32fd8afef1ff460173026b0324049504b3047204d303e002b10169002fff24fe5ffde9fcc1fcdafc27fd97fd1bfea4fe2bffa7ff15007700d00024017701cb011e026c02aa02cd02c7028d021d027901af00d6ff04ff4dfec1fd67fd41fd4dfd89fdf4fd8afe42ff0f00da008901060240023402f4019a014a01230134017901d801290244020d027f01aa00b3ffc5fe03fe82fd45fd44fd6cfdaffd04fe6cfeebfe83ff3300f200b0015b02e6024a0386039c038e035803f30259028d01990097ffa6fee2fd5ffd22fd25fd5afdb4fd27feadfe43ffe4ff88002201a201fc01290229020502cc018a014e011c01f200ca009e006c0036000800eefff5ff1d005f00a800e000ed00c1005c00cdff31ffa6fe48fe23fe37fe74fecafe2bff92ff04008d003201ed01ae025603c703e803ad031b0348024e014a0053ff7bfeccfd52fd13fd17fd60fde8fd9bfe61ff1800a500f7000e01fa00d600bb00bc00e10020016b01b401f1011f023f0250024b022202c6012b0153004bff32fe2ffd67fcf7fbeefb46fceefccbfdc2febdffb100950167022203bd032a045c044704eb0353038c02aa01c100ddff01ff31fe6dfdbbfc27fcc6fbb0fbf8fba5fcacfdf4fe5400a201bb028503f8031804ed038303e6021c0234013d004fff86fefcfdbffdd2fd2afeacfe40ffcfff4b00af00fc002c013a011e01cf004e00abff02ff75fe25fe26fe78fe0bffbfff73000d017f01cc01fd011e0235023e022a02e8017101c300edff08ff31fe83fd13fde7fcfcfc4cfdc7fd62fe11ffccff8c004701f2018002e70218030b03c20242029801d5000a0042ff88fee3fd5ffd08fdeefc1efd9efd62fe53ff50003501e301490263023702d20140019000d1ff12ff65fee5fda9fdc4fd3dfe08ff090018010402a902ee02cf025902a701d200efff0fff3afe79fdd8fc69fc41fc73fc06fdf0fd18ff58008501790218035b034803f1026b02ce012a018a00f5ff6efff8fe94fe41fe00fed2fdb7fdb3fdccfd07fe68fef0fe94ff4300e9006b01b701c30192013701cb006900250008000a0018001d000400c5ff66fffbfe9ffe6dfe77febdfe32ffbcff3e009f00ce00c80095004000d7ff68fffffeaafe7afe7ffec4fe48fff8ffb8006001cc01e301a00114015c009efffffe96fe6efe82fec3fe1bff75ffbdffe8ffefffd6ffa5ff6cff3cff2bff48ff9bff1b00b4004201a201b7017501e400210051ff9dfe22feeefd01fe4cfebafe36ffb1ff1e007800be00ed000201f700c7007100f8ff69ffd9fe63fe20fe25fe79fe12ffd9ffaa005d01cf01e901a5010d013f005dff8efef3fda3fdaafd03fe9efe63ff3200ea0069019e01830120018e00edff5ffffdfed0fed5fe01ff41ff84ffbdffe6fffeff0300f7ffe0ffc4ffb3ffb6ffd9ff1c007300c90002010301c0003b0089ffcafe27fec2fdb2fdfcfd92fe5fff3e000d01ae010b021802d6015301a500edff43ffbefe6afe47fe4efe73feaefef6fe48ffa2ffffff5a00aa00e60008011001fc00d3009d005f002200eaffb9ff91ff6fff51ff32ff11ffedfeccfeb5feb2fed1fe1bff8fff2400c9006601df011d021302c00131017600aaffe9fe48fedafda8fdb4fdfdfd78fe12ffbaff5f00f0006301b201d801da01b6016c0101017c00e6ff4dffc2fe53fe0efef7fd0ffe50feb3fe2affadff3000ab0017016c01a301b801a80171011701a5002600a5ff2dffc6fe78fe48fe39fe52fe95fefffe88ff2400c4005501c901120227020602ac011d0164008fffb3feebfd50fd00fd0ffd7efd43fe47ff63006d014302cb02fd02dd027902e50137018100d1ff35ffb6fe5bfe2bfe24fe45fe85fedafe35ff8cffd6ff1100400068009400ca000c0151018c01af01a901710106017100c8ff1eff90fe34fe1afe48febafe5dff1800cc005801a501a7015e01dc003b009aff1affcffec1fee9fe38ff96fff1ff40007f00b400e60016014301630169014c010801a1002400a4ff30ffd8fea3fe8ffe97feb6fee8fe2aff7cffdeff4a00ba001f017201ab01c901ce01bc0192014f01f1007600e5ff4dffc0fe51fe12fe0ffe49feb9fe50fff9ffa0002c018801ab0190013f01c6003e00beff5eff2fff3eff8aff07009f003701ac01e201ca016401c100fdff3dffa3fe4afe39fe6cfecffe48ffbbff1800560078008b009900a900bf00d600e600ee00ea00dd00ca00b4009d00840069004d0033001c000600eeffcfff9fff5eff11ffc4fe89fe73fe92feeffe84ff3f000701bd014302880284023e02c70135019a0008008bff29ffe6fec2febefed8fe0fff5dffbcff24008800df001f01410144012b01f700ab004a00d8ff5cffe2fe7cfe41fe43fe8afe17ffdcffbe009e015d02e40224031a03ca023d028201a300b2ffc4feecfd43fddefcc9fc08fd93fd56fe3bff27000101b7013c028a029e027a022402a70112017600eeff8eff61ff69ff9cffe2ff20003f003000f4ff98ff32ffe0feb6febffefafe5effd6ff4e00b600040132013e012a01fc00c0007c003f001200fcfffbff0d00270040004f004d003d0025000d00fffffdff02000500f7ffccff80ff1fffbbfe6dfe51fe75fedffe85ff53002c01f8019f0213034a033e03f1026802a501b400a6ff8dfe81fd99fceefb95fb9bfb05fcd2fcf6fd5bffe4007102d903f3049c05b50536052804ab02ee0029ff93fd55fc8efb46fb79fb17fc06fd26fe5aff810083014e02d4020e030103b20230028c01d800260087ff00ff96fe4dfe23fe1afe35fe74fed6fe52ffdfff6c00ec0050018d01a301930162011c01ca0072001700baff5eff05ffb5fe75fe51fe52fe77fec2fe2affa5ff25009d00000146016901660142010701bf0079004200200011000f000b00f8ffc8ff77ff0cff9afe37fefefd07fe56fee2fe98ff580003017e01ba01b7017f011f01ab003800d1ff84ff55ff46ff56ff80ffb8fff5ff2b0051005e004f002400e3ff97ff46ff00ffcdfeb5febcfee6fe2fff95ff0f008e0003015f019101920164010a0196001a00a4ff41fffcfed2febffebefec8fedcfef9fe21ff59ffa1fff1ff42008e00cd00fe002201360138012401ed008e00090066ffb5fe10fe93fd57fd6afdcdfd77fe52ff3c001501c301350263024f0201028901f3004d00a8ff16ffa2fe56fe36fe39fe57fe88febffef9fe36ff75ffb6fff5ff2b0058007b009700b000d300010137016c01910193016101ee00400069ff86feb8fd23fddcfcebfc4afde5fda5fe75ff3c00e7006e01cb01fd010b02fa01d0018f013501c1003900a5ff0eff85fe16fecafdaafdb7fdf3fd5cfeeafe8cff3400cd0044018c01a2018a0154010b01bb0070002900e2ff97ff47fff6feb0fe7cfe65fe71fe9dfee1fe38ff9bff06007800e70048019001b1019f015901e8005e00cdff48ffdefe9dfe84fe8bfeaefee1fe1bff57ff94ffd3ff1b006800b500fd003101460138010101a7003700bcff47ffebfeb6feaefed5fe1fff7dffdfff3100680081007e0064003f001c0006000300150035005a00740075005c002c00eeffafff7bff57ff45ff42ff48ff5aff75ff97ffc6ff02004a009b00ea0029014b0144010e01af003300acff30ffccfe8bfe7afe9bfee9fe60fff3ff900020018a01c001ba017501fa005f00bcff29ffbbfe82fe7ffeadfefcfe5cffbdff15005e009800c300e100f200f800f200e500d400c000a700850052000a00adff47ffeafea9fe93feb1fefdfe66ffd9ff4700a000e00004010e010201e300b700850051001f00f1ffc7ffa6ff92ff92ffa8ffd6ff120050008300a100a50093006e003c000300caff98ff75ff66ff72ff97ffcfff0c0043006b007d007400540029000000e7ffecff15005b00ac00f3001f0127010701cc007f002600c7ff66ff0affbbfe87fe7dfea4fefafe73ff00008e0009016601a101b901b20192015b010f01b0004000c7ff51ffeefeadfe96fea7fed9fe23ff78ffd2ff2e008b00e6003a017d01a501ad018f014e01ef007b0000008bff25ffddfebafebbfedbfe12ff57ffa3fff1ff3c008600ce000d013e015e01660155012f01f600b60073002a00dcff8dff3dfff6fec7febdfeddfe20ff7affddff3e009000d700150144015f015f013e01fe00a3003900cfff73ff2aff00fffafe15ff4cff99ffedff3f008a00cb0001012b0144014a0136010301b90062000600acff5cff1bffeafecbfebefec7fee7fe19ff60ffbdff3000b5004101c101250258024c020402900100016900dbff61ff04ffc9feaffeb8fee0fe17ff52ff85ffa9ffbfffcfffe0ffffff32007900ce0025016c019301910163011501b8005600fdffb3ff74ff42ff21ff13ff1aff3aff6cffadfff8ff43008b00c600e800f100e100bc0090006b0050003b0025000700e1ffb2ff7fff58ff46ff46ff57ff7dffafffe7ff23006400ac00fc0048018901b201af017b011b019a000c0080ff00ff92fe3dfe07fefffd30fe9afe37fff2ffab004801b601ed01f201d20196014f010601b70067001500bbff59fff3fe93fe49fe27fe38fe85fe0bffb6ff71002501b8011c0249023b02f5018401f2005200b7ff2cffc0fe7bfe5ffe6cfe9ffeeafe45ffa4fffbff46008a00c400f4001801270124010f01ea00c00099007400510031000f00eaffbeff8bff55ff25ff07ff09ff2dff66ffa6ffddff000015002b004e007d00a900bf00b800950060002e0012000b001200220034004a0060006e006a004e001300c8ff80ff4dff38ff41ff60ff89ffb7ffe4ff0f00300040003b0028000c00f4ffebfff2ff05001e003b005b007c0092009600810052001800e7ffd0ffd5ffe9fff7fff0ffd2ffa9ff8bff83ff90ffa7ffb7ffb7ffabffa0ffa2ffb6ffd7ffffff27004c0071009600b300c000b7009b006f003f001300ebffbfff8dff59ff2dff10ff09ff18ff38ff60ff8dffbffff7ff30006300880096008f00770054002a00fdffd4ffb4ffa3ffa6ffbaffd8ffeffff4ffe5ffc9ffa7ff88ff74ff6eff77ff8bffa8ffccffedff02000800060001000000030007000400f2ffd6ffbeffb6ffc0ffd8ffeffff4ffe1ffbbff8eff66ff49ff36ff2dff2eff3fff6affaefffeff4c0086009f0098007e005c0037001000e5ffb8ff8aff5eff3eff2bff1fff1aff1dff27ff3aff53ff6bff81ff93ffa6ffbeffdbfff7ff0d001a00220035005e009100bd00c40093002e00a9ff26ffc5fe93fe86fe94feb3fedcfe13ff56ff9bffd9ff020010000b00fcffe9ffd8ffc9ffb9ffb0ffb0ffb9ffccffddffe3ffdfffd0ffb9ffa1ff8bff70ff57ff44ff3eff4cff69ff8cffabffbbffb8ffacff9dff88ff72ff5aff3fff29ff20ff2bff4aff70ff92ffafffc6ffd9fff5ff1b00410061006e0061003a00fbffa5ff44ffe1fe8afe56fe4ffe6ffeb1fefdfe3dff6fff97ffc1fff5ff2e005c00730069003c000000c2ff85ff49ff0cffccfe9afe83fe93fed2fe37ffaeff2b009f00f7002b012e01f5008600ebff39ff8dfefafd8cfd51fd4ffd86fdf6fd91fe3effe7ff7700e3003201600167014301ef007000e2ff61ff01ffc7fea4fe81fe57fe2cfe19fe3bfe96fe19ffafff39009c00d500e600d00096003b00c6ff4dffe2fe90fe63fe56fe63fe8bfecefe24ff86ffe7ff3200620079008000810073004800feff94ff1cffbbfe87fe83fea6fedbfe18ff5effb0ff09005c00880072002000aeff44ff09ff06ff29ff5aff83ffa0ffc1ffeeff1a0035002500e4ff86ff28ffe3fec7feccfee6fe19ff6affdcff6a00f10041014001ec005e00c4ff3effd9fe90fe52fe20fe11fe38fe98fe23ffb7ff32008400b200cf00ea00ff00fd00d7008d002d00d1ff8cff61ff4bff3bff29ff1cff1aff26ff39ff47ff49ff43ff3cff41ff5cff89ffbefff6ff2f0068009c00be00c200a20067002500fbfff2ffffff0a00f8ffbfff6eff21fff3feeffe07ff29ff46ff5fff81ffc0ff1e008d00f9004d01790176014401ed007900f1ff6afffbfeb2fe91fe96febcfe00ff5cffc7ff35009500d000da00c1009a0076005d004e0044003c003a0049006a008b00950079003800ecffb4ffa3ffb1ffc4ffc4ffabff88ff75ff8affc6ff150060009d00ce00f9001c012d012001f000a9006c00500056006d0077005f002a00edffbfffb0ffb7ffbfffbcffadffa3ffb4ffe7ff35008f00e2001e0145015b0163015c0145012201fc00d200a600770043000900d5ffb4ffb3ffd3ff06003b006e009800bd00e4000d012e01420141012f011501f400c50085002c00c4ff6cff3fff4dff9aff0d008700f00041018501cd011702590283027d023c02cb013e01a8001c00a2ff48ff19ff14ff39ff84ffe5ff5100c8004401bb011d024f024402ff0195012501d0009500680041001c000c002e008a000f019c0103022a021802e10199014601db005300c4ff50ff23ff5affe5ff99004901ce0123025c028202970291026002060298012501bc0066001c00e0ffc3ffd3ff18008700fe005d019c01bf01d501ee010202fa01c8016a01fc00aa0089009c00d50013014301670184019c01ab019d016e012901df00ab00a000b500da000b0144018901da012702560254021902bc016901370128013101340124010f01050112012e013a011d01dd00900066007e00cf00300179018d01780163016c019d01e901290246024602360225021602f401ad014501ca005b001600fbff000022005e00c10055010302a20205030703ae02240295012101cf008a0046000c00f4ff1a00860015019801eb010102f101e001e001ee01f801e301b0017a015901520156014001fb008c001900d6ffe7ff4500ca004d01a901d901f001ff010d0215020602dc01a20162012d010701e300bc0096007700690073009100bb00e900150142017501a301c301cb01b00173011e01bd0060001800edffe5ff000035007b00d2003701aa0126029802e502f602bd024302a401fa005b00d3ff63ff0cffd7feccfef3fe49ffbfff4400cc004d01c50131028202a8029e025f02f5017101e2005500d5ff6bff28ff15ff2fff69ffb2fff5ff31006e00b40009016501b001d801d501af018001570132010501bc004e00c6ff48fff8feeefe23ff7affd6ff24006500ac0007016801b401c4018001f000380084fff9fea6fe8afea3feeffe6cff1700d4007b01e401f601b7014301bc003d00d3ff7eff3eff1aff12ff25ff48ff6bff82ff94ffa8ffc6fff1ff1a0031003800370041005e0083009a0090005d001100c7ff8dff61ff37fffcfeb0fe69fe3dfe3dfe6bfeb5fe0dff6bffc7ff21007300a400a800830045000700d6ffabff73ff23ffbffe68fe46fe68fec1fe2fff82ffa4ff9eff81ff5eff39ff07ffc8fe8cfe71fe95fefefe88ff020044003900f0ff89ff16ffa1fe2bfeb3fd50fd22fd37fd8efd0bfe85feeafe3dff8bffdfff3700700073003a00d5ff67ff0affb9fe66fe01fe8afd23fdf7fc18fd7cfdfbfd60fe95fea2fea3feb7fee9fe1fff3cff2efff9feb9fe8bfe75fe71fe6ffe5afe39fe22fe1dfe2afe36fe26fef5fdb4fd7dfd71fd99fddffd28fe60fe77fe7bfe7afe6ffe57fe2ffefbfdd5fdd4fdfefd4bfe9efed2fedffed3feb8fe9bfe74fe34fed8fd6efd0dfdd4fccdfce3fcfcfc09fd08fd13fd3ffd8cfdf4fd61febefe07ff3eff5eff60ff3affe6fe75fefffd93fd38fde4fc83fc1cfcc6fb9afbb9fb27fccbfc87fd3dfed9fe5bffc1ff03001a00fbff99ff04ff52fe9afdf8fc7efc2cfc01fcf4fbfafb1afc59fcb2fc21fd92fde9fd1dfe2dfe26fe23fe2efe3dfe46fe44fe3dfe40fe54fe6efe7bfe61fe12fea5fd3afde4fca9fc81fc61fc54fc6afcaffc21fd9ffdfcfd2cfe3bfe4afe7dfecffe12ff1affd0fe46feb6fd56fd35fd43fd51fd3efd13fdeffcedfc16fd4ffd6afd56fd21fdf4fc00fd59fde7fd7ffef3fe29ff29ff06ffd1fe97fe4ffeeefd82fd1efdd5fcbefcdafc15fd58fd8dfdaffdc8fde1fd00fe2afe56fe78fe91fea5feb3fec2fec9feb9fe8efe4afefafdb2fd79fd4efd2cfd05fdd6fcb7fcc3fc09fd8efd38fedafe50ff89ff8cff73ff55ff35ff07ffb6fe40fec1fd5cfd2cfd41fd85fdcffd04fe24fe40fe6dfeaffef5fe29ff35ff1bfff2fecefeacfe86fe50fe0afed2fdc4fdecfd3cfe91fec7fed7fed3fed5feebfe03fffcfec9fe75fe25fe0dfe42fea7fe0dff4dff5bff52ff53ff6fff94ff95ff53ffd7fe51fefbfd01fe5dfee1fe58ffa0ffb6ffb1ffa7ff9cff83ff4afff6fea2fe6ffe73feb2fe14ff77ffc8ffffff17000f00e6ffa0ff49fffefed7fedbfef9fe16ff27ff38ff60ffb6ff3300a900e900e0009e004e001400ecffb0ff3cff97fefcfdbafd00febefeadff7a00ff0052019e01f001280203025701400021ff62fe33fe74fed3fe13ff36ff7aff1c000f01f4015602f001e500b3ffe2feacfef1fe60ffb5fff2ff4e00fc00ed01c9022403cf02ec01d900fbff7fff4bff2bff05ffedfe18ffa4ff77004f01e1010d02ee01c001b101c201c901920111016d00deff99ffafffffff59009c00c800f8004301a201fa011f02f0017d01fb009f008b00b600f30017011301ff000f016301e801650295025302c0012801cc00ca00050135012e01fa00c900d40028019a01e601e1019101360114014101a70112024f025d025a0260026e0268022702a6010c018e005a007300b100ec0017013a017501db015402b602e502d702a80283027d029502b302b10284023502ce0166010d01c3008d0074007700a000f4006e010602ae024603af03d803b7036103f90290023402ea01a1015901210104010a01300161019101bd01e4010d023f026c028e02a802b702c302cd02c702aa028002520236023f0263029002b302b6029d0273023502e80193013b01f500dc00f6003c01a00106026802ca02250370039c0391034d03ea0286024002240219020502e001ab0186018f01c5010e0241023d020702cd01bd01f6016f02e90224030803aa0253024a029c0219036f034d03ad02d8012f01f9003901a701f001f401c601ad01e6016802f5024a033c03e0027a023b0234024b02510232020402e501ea01160249026e0287029b02b102c502b5026a02f3017a0134014701a50120028902bc02c102bf02c902e002f302e2029f023c02d9019b019d01d10116024c02560236020b02f201fd0129024e0245020a02b2016c016b01b8013602b402040326033a0358037f038f034c03970292018700cfffa2fff1ff80000f017d01dc015802ff02b30333043d04c203fd024102d001b901cb01bf017e012a010d015d010102a602e7028d02c001f0007e008400d1000d010b01f2001a01c701e6020904a9048804cd03f5027402620275024a02a401a400bbff49ff65ffd8ff4e009c00d7003801e701d202a4030f04fa038803f80286023a02fa01b1016001270129016901c90117022602e8017601f40089005300530072009800b300c500ed004e01f901d802ab032c043604d3034003c40275022e02b201df00d3ffe6fe6ffe8ffe22ffd8ff79000601a801820287036504bc045f0463031402d100d6ff31ffddfeddfe46ff26005c019f029403ec039803ce02dc01fd004800b0ff26ffb8fe93fee3feb1ffc700cb016a02860250021e022f027c02c502ad020602f900ecff42ff1eff52ff8fffa0ff91ffadff38002c013502e402ee0263029a01f600a3008c007c004f001700feff22007300b800c20091004f002e003f0057003700c5ff2fffd5fe13fff9ff3e016402ff02f5028102fc019f015d01f700350025ff1bfe86fda8fd67fe5cff1200530048004a00a0003c01c501d6014e016e00acff5cff7affb4ffaaff4fff06ff5bff8a002c025a034703d401b8ff0afe76fdc1fdf8fd3cfd8efbf9f9ecf921fcfbffc603d0058905d40353021f02f7027603380209ff32fba8f8aff8eefabafd4fff16fffffdabfd0fffa401b803b3034f01defd5cfb10fbb4fccbfed6ff6aff6dfe3efe84ff9f011903ce02ce0054fed5fce6fcd6fd49fe60fd72fbd9f9e3f9ccfb8afe8c00e700fcff1aff66ffe9007b02ac02eb000cfebffb51fbc0fcb9fea0ffc7feeefcacfb30fc4ffe9b006b011c0080fd47fbbefae5fb89fd40fe88fd2bfc96fbb9fc3cffb701b702cc01ccff2bfed8fd94fe35ff9dfea6fc4cfaf3f861f92ffb20fd13fed1fd20fd15fd2dfee9ff30013301f8ff4cfe22fdd6fcf7fcbdfcc2fb68fa95f906faaefbbcfd26ff60ffb2feeffdb9fd0efe50fed4fd85fc08fb47fac8fa3cfca9fd26fe7ffd53fca2fb0ffc5bfd9ffef4fe14fe8cfc52fb07fb99fb5ffc9afc1dfc63fb1efbb5fbedfc0bfe6ffe01fe37fdbbfce4fc67fdabfd3dfd24fcf4fa57fa85fa3afbe5fb13fcd0fb8efbb0fb49fcfbfc42fdf0fc4ffcd9fbf6fb94fc2cfd40fdb5fce4fb71fbc7fbbcfcc0fd3afee5fd0cfd39fcc1fba7fb90fb12fb27fa2ff9a2f8d8f8c5f905fb3dfc40fd12feddfe9eff1000f0ff21ffc3fd44fc0dfb45fae3f9baf9a0f9a4f9e9f977fa3cfbf7fb5efc6efc55fc4bfc83fcf6fc56fd61fdf5fc2dfc66fbf8fa02fb74fb0cfc8efcf7fc58fdabfde3fdd7fd5dfd84fc7efb80fab7f930f9e1f8e1f847f919fa4dfba3fcb5fd49fe5cfe1efedafdacfd78fd18fd77fcb3fb27fb19fb7ffb16fc71fc47fcb6fb1ffbd9fa0cfb84fbddfbe2fb9afb4efb5efbdefb91fc24fd5afd36fd09fd1cfd82fd0cfe5bfe20fe63fd64fc77fbe4faaefaaefac6faecfa30fbb7fb81fc63fd23fe84fe69fee9fd28fd58fcb1fb56fb52fbacfb50fc1afde6fd8efef4fe12ffdffe5bfe9bfdbdfcedfb60fb2ffb4dfba2fb0bfc71fce8fc88fd54fe26ffb2ffb8ff2fff46fe56fdb7fc7dfc7bfc73fc41fc05fc12fca9fcc9fd21ff2900780002000fff15fe76fd3efd36fd23fdf1fcc3fce0fc72fd66fe64ff05001500a5fff7fe55feebfdabfd72fd2dfdeafcd0fc0bfda2fd75fe4dfffbff6c00a500ad008c004000c0ff12ff59febffd63fd50fd7bfdd2fd3efeb1fe2cffa6ff09003d003300ebff86ff2bfff8fef9fe25ff65ffabfff5ff4700a000e800ff00cf006100d8ff67ff33ff3cff5eff6eff5fff4fff67ffc0ff4800c500f600c7005d000100f8ff4c00ca002f014a012401f600eb000f0147015b012e01e200b400ce002b018f01b3017201e3005000070022008300f6004c017f01ad01e6012702590259021f02cf0193018b01bc01090253029302c302e402ec02bd0243029301df0062004b008d00fa006001a901ee015b02fc02b70354048c045004ce034003d902af02a002800245020202d901ee014702c9025403c203080423040804b30331038e02e801710140015801b7014d021603130428052706d406e40640061d05cc03a702f001a0018e019c01c5012a02f20208042405eb050d068e05cb042c04f6032e0483049b045a04e2037e037503c10330048e04b504b804d2041f058905e105e4058405ef045104d20391037c038003ae030b0490042d05b105f6050206eb05d705de05e405c20577050805a2048304ac04f604320533050705f2042205a8057106290784077207f8063d067c05c304180495034b035203c603930490059706700701085708660824089707bd06b705ce042d04f8033a04ba044305ca053d06a0060507490751072407c60658060d06e405c00590054a0515052f05a1055b062a07b007cd07b30791078b07a5079707200747063c05670429047f042a05d805390657067806c0063d07d6072e080f089107de063a06e105c805d405ef05fd050a063e069a061807a7070f0832080d089407e4062e068005fa04c404d6043005d30590064007cc070f080008bc074907c2064906e0059d059c05d1053106ab060b0738073c071d07f706e106be067e062506ba05650556057d05bb05f3050106fe05290694062e07c407ff07c007340792061b06e705c10579050f05aa049c0421050d060607a907ac0726077106cb055305fa048c040904b303c7036f049805d306b5070a08cf074507b6062f06a5050b055b04c1037f03a7032c04de047005bf05d705c505a5058e0568052a05e804a9047904610449042204f003c603d7034304ec04a5053b066a0622069505e0041a045903a3020202a101a901360236035c045605e605ed058e0509057604dd0341039102e201790183010b02ef02d8037404a40470040b04b303790350032603da026d02fe01a3016f017301a401f5015802b202f10210030603dc02a6025e02fe018d011001a5008000bf0061013d020703800397035503e1026702e7014a0186009effbefe29fe0dfe79fe57ff71008b017e022c0389038d032e03790290018f0099ffcffe38fecefd97fda7fd10fed8fee0fff800df0153023c02b301dd00e0ffe2fef9fd36fdb1fc87fcd1fc92fdabfee5ffff00be01ff01ba01fe00efffbbfe90fd98fceffba1fbb0fb10fcaefc7afd5efe30ffc4fff7ffb6ff0dff31fe64fdd7fc96fc93fcaefcbffcc2fccffcf4fc38fd91fdddfdf5fdcafd5afdbbfc10fc79fb18fb03fb34fb9ffb29fcabfc11fd55fd72fd6ffd4bfdf7fc79fce4fb51fbe0faa8fa95fa8ffa85fa78fa8ffaebfa7bfb13fc75fc68fcf8fb6bfbf9fac6fabefaa2fa5afa01facff9fbf980fafefa22fbcdfa27faa5f9a8f928facafa08fb93faa8f9d0f877f8d2f89ff947fa78fa44faf7f9f3f94dfaacfaadfa17fafff8e6f747f73bf7a3f72ef886f8b0f8e2f833f9a8f912fa23facbf92cf973f8e6f797f75df733f71ff722f767f7ecf76af8b9f8caf89df875f883f8a8f8b5f86ff8aff7b8f6f2f59cf5d9f575f607f76bf7aaf7d5f723f885f89bf838f863f75af6acf5b2f546f613f796f76ff7d9f649f602f626f675f677f619f69cf555f5a9f58df67ef70ff807f875f7d5f679f647f615f6a4f5d5f40ef4cdf33af44df59cf695f70ff81af8d6f786f72bf78bf6b1f5caf40cf4d9f341f4ebf495f504f616f611f62ef65af688f68ff642f6d5f57df54af553f577f577f566f564f57af5c9f52ef656f63bf6eef587f559f57bf5aef5c7f59df525f5c1f4c3f430f5f4f5b9f60cf7e6f672f6ebf5a4f5a5f5a2f57cf52bf5c4f4a2f4faf4aef58ff63af753f7f3f651f699f51bf5ebf4e0f4f9f42bf55cf5a0f5fbf54ff6aaf606f746f769f752f7ddf62ff67ef5f7f4e7f451f5ebf584f6e9f6fcf6f6f6fdf603f704f7dbf66df6f6f5bcf5dcf56ff634f7bbf7e1f7adf745f701f709f735f75ff75af714f7cff6c2f6ecf645f795f799f76af73bf735f785f70cf875f895f863f8fef7c2f7def738f8a6f8e0f8b8f863f82bf83af8a6f83af995f98ef928f98bf811f8e5f7f6f737f885f8c5f814f988f918fab3fa2cfb5bfb45fbf3fa7cfa0efab4f963f929f9fff8d9f8d0f8f1f83ef9c9f984fa45fbf1fb61fc7efc68fc34fcecfba7fb5afbf8faa0fa74fa8cfaf6fa85fbf6fb30fc3afc36fc64fccdfc3bfd75fd47fdb1fc03fc92fb80fbc3fb22fc69fc98fccffc32fdd7fd90fe13ff37fffcfe8afe26feeffdd2fdb7fd84fd3ffd12fd22fd80fd1ffecafe55ffb7ffecfff9ffe9ffb9ff6fff26fff5fef9fe44ffbcff3a00a500ec00120127012e011a01dc006800d8ff5dff22ff4bffdbffa300710117027c02b102c902ca02b80289023202ce0186017501b1012b02b6022803680372036703610363036e036b0347030d03d602c102f0025f03f403a3044505b805fc050b06e10596052d05ad043a04e303b003bd030f0497044e051006b406290752073407f906a9064f060c06d605a1058d05a005e2056e062807db076a08ae089f086a082508e807d107c407ae07a907b107c407fc073d0866087c0878086d088c08d20829098e09d609ec09f109e709d509d009bd0994097c0974098009b709f009090a140a0c0a090a3d0a8e0ad90a170b240b090bfe0a0a0b2e0b720b990b8b0b6b0b430b2e0b590ba20be60b1f0c1e0ced0bc70ba80b960bb30be20b0e0c4f0c8d0cc40c080d350d360d1e0dd20c600c080cd40bd30b200c870ce50c3d0d750d980dd20d040e1b0e1a0ed80d5f0dfa0cb70ca70cda0c0d0d1a0d200d190d210d760df00d5c0eac0eb70e8b0e740e7a0e9b0ed10ecc0e6b0ed80d290d960c6b0c890cc90c2e0d940dfc0d990e4e0ff00f61104d10a40fb20eaa0dcd0c600c400c500c9b0c080da30d8b0e810f4210b0108e10e40f0d0f2f0e620dc40c300cac0b770b9c0b2e0c360d580e4b0f031059105e104310e80f380f4f0e260df60b280bd00aec0a770b290ce70cc50d9d0e530fd80fdb0f440f540e320d260c840b350b200b490b8b0be90b8e0c4e0d010e8e0eaf0e570ec00df90c2c0c960b2a0be50add0aeb0a050b480b8d0bc70b080c2c0c2c0c260c080cdf0bd30bc60bad0b960b630b150bd90aa60a7d0a670a3f0a0c0af309e509ec091b0a3a0a320a1d0a000af6091d0a4d0a680a680a310ad8098f0950091a09ef08ab085c08360835085a08a308d608da08be08800840081a08f407c607a1076d073c07320738073f0752075807500751074f0746073e071d07de0695063c06db058905470516050105fd040d0536056c05af05f40517060c06d4056c05f6049a04570428040304d503a003750365037d03aa03c603c2039b0358031c03fb02e702d502b5027c0245022202130215021a0212020502fc01fc010b0219020502cb016f01fa008b002c00ddffa4ff81ff78ff9affe3ff3d009500cd00d600bb0081002e00d5ff71ff01ff9efe5bfe3ffe4ffe72fe8afe84fe54fe09fec1fd88fd68fd67fd73fd85fda5fdc5fde1fdf0fdd7fd93fd3afdd8fc87fc5afc3efc26fc08fcd5fba1fb8bfb8afb9ffbc2fbd3fbcdfbbdfb97fb6cfb4afb1bfbdffaa3fa5cfa18faecf9d3f9d6f9fcf92cfa61fa91fa94fa6efa36fae6f996f958f910f9bff879f83ef828f847f876f89cf8a6f87af836f803f8e2f7ddf7edf7e7f7d1f7cef7e4f724f879f89bf86ef8eff729f761f6d1f572f54cf54ff553f56bf5b4f521f6b5f653f7b0f7c1f78df70af767f6d0f53ef5c5f46df420f4f6f303f430f48df410f584f5e3f526f62cf607f6c6f554f5c7f437f49ff324f3e3f2d0f2fbf257f3aff306f45cf491f4b2f4b8f487f440f4faf3b4f392f38df370f33bf3f2f28ef251f25ef295f2edf23bf347f332f31af3f9f2eef2ecf2bdf276f233f2fcf103f24ef29ff2e8f216f315f317f32bf327f30cf3c8f23ef2a5f12ff1e2f0e1f017f14bf186f1caf1fef142f295f2c9f2e9f2eff2c0f289f25af21af2edf1d2f1a5f17ef158f110f1d1f0adf09cf0cef045f1c8f158f2dbf21cf339f334f3edf289f20ef265f1c8f05cf01bf030f097f016f1b0f14bf2b7f20ff34ef34bf32cf3f0f272f2e8f16cf1f1f0b1f0b1f0c4f0fff058f1a0f1f7f165f2c2f222f376f386f36cf331f3c6f262f21bf2d8f1bef1c8f1c6f1d6f1f9f107f224f254f273f2a1f2daf2f7f21bf34bf367f38cf3b4f3b3f3a8f398f369f342f327f3f2f2baf28af257f259f29af2f8f27bf3fef34bf47bf494f484f474f45ef425f4eef3c6f3a4f3bbf306f44df498f4d3f4e2f4eaf4ecf4d1f4b3f489f446f425f434f45cf4b3f41df564f5a7f5e8f511f647f67cf67af651f607f699f543f51af506f51ef55af59df508f698f622f79ff7edf7dff795f72bf7aef659f635f623f62ef651f67cf6cff647f7c7f751f8c3f8f3f8f9f8ddf89ef86ef85af845f832f81af8eef7ccf7bef7c1f7ecf737f885f8e0f843f9a0f904fa5dfa89fa8dfa6afa23fae9f9d4f9d6f9ebf9fcf9f4f9e4f9d9f9ddf90cfa5afaa5fae5fa0ffb1ffb38fb61fb8efbc4fbeffbfafbfcfbfffb02fc14fc2bfc32fc31fc2bfc23fc2cfc44fc5cfc78fc95fcb2fce8fc37fd87fdcefdfcfd09fe0dfe1bfe2ffe48fe55fe44fe1dfef3fdd9fde6fd15fe4ffe8efed0fe18ff73ffd7ff2c005f00660043000c00d6ffaeff96ff88ff86ff95ffbbff06007100e7005501ad01e401ff010402f301d301a9017b015f015b0167018e01c90103023a026e029702c002ed0213033a035e03730384039203a203c203ed030b0416040504d603a1037f038203bc031d048704ee043b0560057505800586059605ac05bb05cd05d605d305d805de05dc05e405eb05ea05f805110637067806bb06ef06270752076e079a07c907e9070208fb07d807bf07b207b007cf07ec07f107f907fa07fd0728086708a808f90834095209790994099b09b009b809a5099e098d0968095909540956098509c909070a510a890a9f0abd0ad70adf0aee0aea0ac70ab50ab10ab90ae40a0b0b150b200b230b260b550b900bb60bd90bdc0bc40bc90be10bfb0b280c400c350c2d0c220c160c220c1f0c000cf40bee0bf30b270c690ca20cea0c210d440d7a0d9e0d940d760d2e0dc50c7b0c500c450c760cb60cea0c2c0d5b0d6d0d870d8e0d7e0d840d910da50dde0d100e1b0e160eea0d9b0d620d360d110d160d210d290d560d900dc60d110e480e530e520e380e0e0e010efc0df70d0f0e230e260e320e240ef60dc90d8c0d4c0d3d0d470d600da50dea0d1f0e640e960eaa0ec30ec30ea20e830e4d0e030ecc0d8e0d4d0d3a0d3b0d480d7c0daf0dd10d020e210e2a0e430e510e480e4a0e380e0d0eeb0db60d6e0d420d220d0c0d250d4a0d6a0d9f0dc40dd30ded0df20ddc0dcc0daa0d750d570d360d110d090d000df30c030d0c0d010d000dee0cd00cd60ced0c0f0d4a0d6e0d6b0d5e0d350dfa0ccd0c940c510c260cff0be50bf80b0d0c170c290c230c120c220c380c500c7a0c8a0c7f0c7e0c670c3d0c1f0ce90b9a0b5b0b1e0bec0ae40ae30ae80a0e0b340b540b870ba20b910b760b450b0b0bef0adb0ac60abd0a9e0a700a590a450a340a3d0a3f0a310a260a0b0ae709d709c409b109b909c609d409ec09ec09cf09ac0971092f090809e608c508b30894087208670863086d089408b208c008ce08c408aa08990875083808f10793073407f906d406ca06e70602071007260738074b076d077c0768074107fa06a506650633060f060106ec05c6059f05700540052e052e053e05650589059d05a905a10584055f052f05f404b70477043e041904fa03e203d003b50395037b03630356035c0368037f03a603cd03ea03ed03c2036e03fc027802fc019b0154012e0130014e018e01e30133026c027f0266023102e60185012101bf005c000b00dcffcfffedff280067009f00c000bb0096005400fbffa3ff56ff18ffeffed5febffeb3feadfeacfeb8feccfedafedefecbfe9ffe64fe1afec5fd76fd37fd14fd13fd2cfd5efd99fdbefdccfdc2fd90fd44fdf2fc92fc31fce0fb9afb6dfb67fb7cfbabfbeefb25fc44fc49fc20fcd7fb8bfb42fb09fbe7fac8faaffa9efa89fa78fa72fa6afa65fa61fa4bfa2cfa10fae7f9c0f9a0f97af95df953f94cf94ff95ff969f975f982f97af964f93cf9f4f89ef84df8fcf7cbf7c1f7c5f7dcf701f81df83ff868f87bf880f873f83bf8eef79ef746f701f7d5f6abf693f695f69ff6c6f60af749f77ff7a2f792f76af739f7f0f6acf677f639f603f6ddf5b3f59df5a4f5adf5c9f5fcf528f657f687f697f68cf66af61ff6cef58ff557f540f54bf557f56ef58cf593f598f59df587f56bf553f52bf50ef504f5f2f4eef4fdf401f511f534f546f550f54ff528f5fcf4def4c0f4c1f4def4ecf4f4f4f8f4e1f4ccf4c6f4b3f4a8f4aaf49ef49cf4aaf4acf4b7f4ccf4c8f4c8f4d3f4c8f4c0f4c1f4a7f48ff48bf483f48ef4a7f4a7f4a8f4aff4a0f4a4f4c4f4d0f4d9f4e1f4c6f4a5f496f480f478f480f477f479f491f49ff4bcf4e9f4faf405f515f510f510f51cf50ff501f5f3f4caf4abf4a1f48af486f49af4a5f4c2f4f4f413f531f547f539f531f539f531f53af554f550f549f54df541f543f556f54ff544f539f512f5f3f4edf4e7f401f53bf56af5a5f5ebf511f62af63bf627f607f6e1f59ef561f535f506f5f9f416f53bf57af5cff515f65df6a2f6c0f6caf6bdf678f621f6cdf573f53ef53ef557f595f5eef53df68df6d8f609f72ff73ef71af7e1f69bf63df6f7f5ddf5d8f5f6f530f663f69df6daf605f72ef74cf748f736f719f7e6f6c2f6b5f6adf6c2f6ecf611f745f77ff7a5f7c2f7d1f7bcf79bf771f735f709f7f2f6e0f6ecf611f73af779f7c8f70bf84ff88af89ff89ef88af855f81bf8e7f7b0f799f7aaf7ccf70df85cf890f8b4f8c7f8b7f8a4f89cf888f876f86bf857f858f881f8bbf808f959f98af9a1f9a9f99cf98df980f963f944f928f909f904f91bf937f95af982f99ef9c0f9eef917fa3cfa57fa59fa52fa49fa39fa34fa38fa32fa36fa49fa63fa91facbfaf8fa1efb3bfb43fb44fb3ffb26fb08fbe6fabffaabfaadfab7fad7fa09fb3cfb7cfbc8fb0efc50fc87fca3fcaafca2fc8cfc75fc5bfc38fc20fc10fc00fc00fc14fc2afc4afc72fc96fcc1fcf1fc1cfd4efd82fda5fdbcfdc6fdb9fda5fd97fd8cfd8cfd98fda1fdacfdbdfdd2fdf2fd18fe3afe56fe6afe77fe84fe8ffe92fe91fe8afe7cfe78fe8cfeb9fef6fe33ff65ff8dffa8ffbdffd2ffdfffddffcbffacff89ff72ff70ff86ffafffdcff0800320054006b007b0081007d007e0087009900b600d900ff0022013e01580172018101870185017a016a0160015e0164016b016e0174017f019501bc01ef01250258027e029502a802b902c602ce02cc02c102b402a702a302b302c802d702e602f102f502020315032803400354035e036e0385039f03c503f003130435044804430434041604eb03ca03b503aa03b703d503fa0331046f04a804e00409051b0524051f050905f604e204c604b204a1049604a604c604ec0428056b059f05ce05ee05f305e905d205ac058c056f0552054805500562058e05c905ff053706660682069b06ab06a906a40696067e06730670066e06740676066e0671067e069406be06e70602071e0732073a074d0761076907710772076b077107750774077f07870788079907ab07b207c307d107d607ec070a08230840084e084b084f084f084f0862086c086508660860085708690881089708c008e508fe08220939093a09400937091a0911090b09020915092c093a0954096509650972097a0979099009a809b209cd09e109e509f609040a070a170a200a1f0a320a440a480a5a0a670a600a610a5a0a420a380a2c0a1a0a210a350a500a830ab60ae10a1b0b490b620b7d0b7c0b5a0b390b110beb0ae80aee0af40a0d0b1d0b220b3a0b500b5d0b720b730b600b600b620b6c0b950bb40bc10bdc0be80be70bfe0b0e0c090c0f0c060cf00bf60b010c070c230c2c0c1a0c170c080ce70bdd0bd60bc60bce0bdb0bea0b180c470c6c0ca60cd40cec0c0a0d100df50cdd0cb20c740c4a0c1f0cec0bd80bc80bbb0bd50bfc0b230c640c950ca70cbb0cbd0cb00cbb0cc50cc50cd10cc90ca80c950c790c560c4e0c3d0c1b0c0d0cfa0be60bf70b0b0c150c2d0c330c260c280c230c180c250c260c190c240c2b0c2b0c440c520c4b0c4d0c370c080ce60bb60b790b570b330b0c0b070b060b010b1a0b350b480b700b8e0b9b0bb30bb90baa0ba30b890b560b2a0bf40ab70a940a780a5a0a4f0a410a2a0a260a230a1c0a250a240a160a160a120a080a130a1d0a1f0a2b0a2f0a220a140af209bc0986094209f908c4089808700860085f086808820896089d089f088d086d0854083e08290822081b0811080d080808fe07f307d4079f0765071e07d306970665063b0621060d06010605060f0620063f065b066c067406680649062006e605a1055e051705d1049c0475045d04580457045704580450043f042d041004e903c1039403670346032b0319030f030403fb02fa02f602eb02da02ba0287024a020502bd0175012c01eb00be00a500a100af00c800e400f90003010001ef00cd009c005a001100ceff93ff61ff3eff24ff0efffcfeeafed4febefe9ffe77fe4dfe20fef3fdcffdaefd93fd84fd7afd73fd70fd64fd4dfd34fd15fdf4fcdafcb7fc8bfc5bfc1cfcd8fb9ffb6efb44fb26fb0bfbf8faf6faf6fafefa11fb13fb00fbdafa95fa43faf9f9b3f97df961f94cf946f952f95af962f96df963f944f913f9c2f869f81cf8d4f7a1f78bf77af77bf78df796f7a5f7b9f7b1f798f76ff724f7d4f691f648f614f600f6f2f5f9f514f620f628f632f618f6f3f5cdf58cf543f501f5b1f472f455f43ff445f467f478f486f497f48ef486f483f45df428f4f4f3a6f362f343f328f322f330f327f31ef323f312f305f304f3e4f2b9f293f255f227f215f2faf1f0f1fff1f9f1f9f10df208f207f212f2fef1e7f1d9f1b1f18ef17af14ff12ef126f10af1f7f0f9f0e1f0d1f0d3f0bbf0a9f0a8f090f083f089f07cf07ff09df0a4f0b1f0cbf0bff0aef0a7f07ff05bf046f015f0e8efcfefa6ef97efaeefbbefd5effbeffeef01f013f00ef014f028f01ef017f01af003f0fcef0cf0ffeff2efecefc8efaeefaaef95ef8fef9aef91ef9aefb8efbeefd0efeeefebefebeff8eff1effcef19f01cf029f043f041f043f04cf036f028f023f000f0ebefe7efd0efceefe7eff1ef11f043f05bf076f09af0a2f0b8f0daf0def0e5f0f0f0dff0ddf0eff0ebf0f4f00af1fff0f6f0f7f0e1f0d9f0e5f0ddf0e4f002f10ef128f153f169f18ff1c9f1e9f10bf233f239f23cf246f239f236f243f235f22af22af215f20ef21ef21ef229f246f250f266f28ff2acf2d7f214f33bf366f397f3acf3bff3d7f3d4f3d7f3e5f3dbf3d0f3cdf3b7f3adf3b4f3acf3b1f3c3f3c6f3d9f304f42af461f4a5f4cef4f3f419f526f538f550f555f55ef56cf569f575f58ff59af5aef5c8f5c8f5c6f5c6f5b4f5abf5aff5adf5c1f5ebf512f645f681f6aef6e4f61df73ef75cf776f776f775f77af776f77af784f782f787f791f792f7a2f7c0f7d2f7e7f701f811f82bf855f87ef8b0f8e5f809f927f941f94bf95af96ef979f984f993f998f9a2f9b7f9c7f9d9f9edf9f7f9faf9faf9f5f9fef916fa30fa53fa83fab1fae1fa15fb40fb66fb87fb9cfbaafbaefba3fb96fb8cfb81fb80fb8dfb9ffbb7fbd2fbe6fbfdfb1bfc3afc5cfc7bfc8dfc98fca1fca8fcbafcd6fcf1fc10fd30fd49fd65fd83fd99fda8fdadfd9ffd91fd87fd82fd89fd99fdaafdcafdf6fd21fe52fe84fea6febffeccfecafec8fec8fec4fec5fecffedcfefdfe31ff68ffa1ffd6fff9ff0f001d0019000b00faffe4ffd5ffd4ffe2ff090045008600c500030137015e01790183017c016d015b014d014c015e018101af01df010902310255026b0277027d0273026502620268027b029f02c602ef021a033d035b0381039e03b203c603cd03cf03e203f903120436044e045304590455044a044c044d044f04620475048904b804ee041f055d059405be05ec050a0616062d063e06480663067b0687069e06ab06ae06c106d506e40606072307340757077d07a107d70708082b085b088808ae08e808210952098e09c009e009090a280a350a460a4a0a3f0a420a440a440a5f0a830aa70ae60a250b5d0ba80bed0b220c620c970cbb0ceb0c0d0d210d470d630d700d8c0d9a0d950d9e0d9c0d8b0d8f0d8e0d880d9e0db60dce0d070e3e0e6d0eb80efc0e2c0f690f900f9a0fb20fbb0fb10fba0fb20f930f8a0f780f580f5b0f5a0f4a0f550f590f520f730f980fb50ff30f261042107910a710c310fb10261135115a116c1160116c11681146113a112311f910f710f210e210ff1021113c118811d71117127b12d2120913531386139813bf13d313c713dd13ec13ea1311142f143314551467145d1478148d149214c114ec1409155815aa15f4156e16de163117a117fc172f1875189f189f18b118a1186f1868185d184018591874188318ca1812194c19b519101a481a9e1ad71aed1a2d1b5c1b6c1baa1bdb1bef1b301c611c6e1c9d1cb01c971c9d1c861c4c1c431c311c081c201c401c561cae1c041d401da71df51d151e4f1e631e461e4a1e321ef41dea1ddb1db51dc81dd51dc61ddf1de41dc81dd71dcf1da71dae1da81d871d9a1da61d981db41dc01dad1dbf1dba1d931d891d5f1d0e1dd91c871c161cca1b6e1bfc1ab71a6f1a201a041ae319be19c619c019a619ad19981965194319f91889182818aa17121795160a167f151c15b1144114f2138e131913b9123d12af113411a3100a10910f140fa30e610e230eee0dd20d9e0d580d140da40c170c860bcc0af9092c0950087f07d2063006a4053a05d00473042a04d60383033503d2026702fc017e010801a4003b00e5ffa0ff57ff1cffebfeaefe72fe33fedbfd79fd0afd81fcf7fb6bfbdefa6cfa0dfabff997f981f976f989f99df9a8f9b4f99cf95ff917f9acf82ef8c2f74cf7ddf696f652f61cf60ef6fbf5e6f5e3f5bff584f54ef5f2f488f430f4c0f359f31df3d9f2a6f2a1f28df27df285f261f221f2def15bf1bcf024f067efb2ee23ee82edffecb8ec65ec2dec2aec0bece4ebc9eb72eb01eb97eaf3e944e9ace8f0e742e7c3e62fe6b6e571e50ce5a7e459e4cee331e3a2e2e1e126e193e0e4df54df07dfaede7cde8dde87de8edeadde8bde57de25dea6dd1bdda1dcecdb45dbccda2edab3d978d924d9f5d8fdd8ddd8d3d8efd8d0d8c2d8dad8b9d8afd8d8d8d2d8e8d82ed942d96cd9c0d9d3d9e6d909dad9d9a4d97fd913d9bfd897d83bd80ad81ad806d81ed873d89ad8dbd842d96dd9a6d9f7d906da28da67da68da83dac4dad2da04db5cdb75db9edbdddbd4dbd3dbdfdba1db6ddb4ddbeedaaada91da5ada57da88da9cdadeda4adb90dbf6db72dcb3dcfcdc43dd45dd4edd60dd49dd53dd74dd7eddb9dd12de5ededede72dff1df9ae04ae1e0e19fe262e30de4dee4abe55fe633e7f3e792e84de9f5e988ea45ebfdebb5eca4ed9ceea4efecf03ef2abf354f5f8f6a5f875fa29fce2fdb5ff5a01f902a50415067707e408160a430b7d0c850d960ebf0fc710ec1136136b14c7154417a818321ad11b4e1df01ea3202d22ce237225e4266928e929372b8e2ccb2dc62ebe2f893004317931bc31b231a73179311f31e630ac306c30673071308630da302b316d31c831f031dd31bc31423179309d2f762e232de52b892a30291028e526ce25f8240d241d234a223c210720d81e6a1de01b6f1ae1185e170916a71463134d121911e80fc00e4c0db30b090a0e0802060f040b023900c1fe73fd7ffcf5fb8cfb5dfb65fb4ffb22fbd8fa31fa49f935f8d9f664f5f5f385f23af125f03bef96ee2ceee5edc8edbfedb4edb3edaded9eed9beda1edc2ed0aee62eed9ee7aef1cf0c7f083f11bf28af2d7f2e0f2b8f277f20cf2a5f15af115f108f141f194f126f2f1f2aef376f441f5bff512f641f60cf6a2f51df546f463f39ef2b6f1eff06ef0e2ef81ef6def47ef2cef36ef05efc2ee8dee0fee74ede9ec17ec37eb79ea82e98ae8c8e7dae6ede52ce52fe428e342e217e1dedfcede8cdd4ddc48db1fda10d950d880d7d1d66bd6e8d578d53ad5c4d441d4ced30dd337d272d173d07bcfaacebacdf5cc76ccfbcbc8cbe4cbf7cb3acca2ccdbcc2bcd86cd9bcdbbcddecdbbcdb6cdd1cdc2cdedcd56ceb1ce59cf47d02ad155d2b9d306d58ed640d8ced983db47ddd2de6fe0fde137e37be4a2e55fe618e7b5e7e9e71ee846e819e8ffe7eee7a0e780e782e772e7ace72be8a9e873e988ea89ebc3ec2fee5def98f0e1f1ccf296f34ef498f4b1f4a5f425f471f39ff26cf12ef008efb9ed8feca9ebcdea3cea02eacde9c7e9e0e9b4e968e9f9e821e821e712e6c2e478e35ee24fe18ae031e011e036e09ee015e192e1fee149e276e272e24ae220e2e0e1a6e194e17ee177e195e196e17ee154e1d4e01fe053df50de6bddecdcc4dc63dd04df83e132e50eeaa2ef00f6d4fc6403b0095e0fc71333178d19781aa01a451a38195018e117a7174918d019ac1b3f1e4f2124241e27122a722cca2e233127338b356e388d3b7a3f0c44d1481f4e76533858b85c7160e762ab647d653965c36416643463fe624b63ed63776569674e69726b1b6dd06df16d026de86a4f680d6562611b5e1b5bb7588c57245794571a59d85ab05cc45e16609f60bf60b95fc05d7a5b6a58eb54a851204e924a734712449440493d5f39f5347a30512bcb259220501b6e169012600f330d690c670c480d230f0911eb12dd14ff15661676169015fa1361125f10370e960c0d0ba609d7080d08140743060e0546035e0109ff4cfccdf977f76cf552f409f48af444f6dcf810fc160062049408e70cd41011140d177a19371be61c5d1e7c1ff0208f22132403262028ff29032ce12d2a2f48301631473159314e31063108315e31f531383306353037f439f83cff3f3c433f46c848264b004d3c4e4f4f02504c50925090502f50c64ffe4eb54d3c4c2b4a764782440f41483dbd394a362c33e730432f642e962e6b2fd730e332e334bb366b384a396639f53881375435d732c22f7e2c82297226a2236d21501f681de41b301a531878162c149a110f0f530caa09520716054c0317022001a400a0009400a300ce00a70063002800b6ff4cff18fff9fe01ff66ffe5ff74002a019a01b2016a0180000aff25fdd3fa57f8f1f5cdf33af25bf143f115f2adf3e4f5aaf89ffb7dfe2c015303c804a005b50523053304d7024701deff79fe31fd4efc87fbd4fa56faabf9c2f8bef74df68bf4baf29bf06dee90ecbeea36e94de893e72ae74ee760e75ce787e757e7dce665e67ce54fe446e3fae1ace0b6df8ade52dd52dce1da25d95ed7ead402d2fcce50cb63c7b6c3e6bf78bce7b9a2b713b690b553b592b579b621b7acb73fb816b885b7dbb677b5e2b38fb2f1b093afd7ae1aaecead26ae59aecaae96afebaf32b096b060b026b034b0eaafedaf83b0ffb0eab168b3bbb44eb623b876b9b0bac1bbffbb1bbc19bc55bbdcba98baf6b9efb951ba84ba2dbb2dbcb1bc47bde2bdc8bda1bd7ebdc5bc3abc09bca6bbcfbb95bc41bd65bed7bfafc06fc1ecc147c128c09abef3bb12b93eb6fdb24ab06aaeb8acf1ab24ac70ac49ad93ae5faf19b0adb052b095af95aed6ac15ab84a9c5a78aa6dca53da52fa57ca586a5b2a5bca526a56aa454a3a3a103a0559e789c249b209a3399d798a0983698f39767977c96b895e6945f94e894639651996b9e55a549ae6fb9bcc5e9d287e018ed53f8e9018808750c150ebb0c65093905060001fb52f791f481f3aff424f717fb8e0041063f0c93122e187c1df422f5271c2d053335391b40f04702506d58d8605668216fd6745a78037a237abc7830779975e4733b737e73537425769d78f27a287dca7e2e7f697e557cf478d3742a70886bb167c5644563a06353656e68e26c83710776397adc7cdc7d6c7dc47a4e76c170c1690062445a3052624a56435e3cce35d82f9e2967236f1d0c17b710cd0aeb04c3ffa4fb29f8faf51ff5d8f48ff509f745f88ef9bbfae3fa5efa4ef91af741f428f175ed8de9c1e5cbe1dadd0bda0bd6e1d193cdf2c824c45bbfaeba69b6eab26ab01faf47af0ab164b43cb95bbf67c611cee7d56ddd61e46bea40ef05f3a6f506f7b0f7d7f76cf70bf7f0f6dbf646f750f879f90bfb19fd08ff130169038505a207150a7a0c080f1d1277153a19a11d6d22ac27642d3d333d395a3f0245724a7a4f94531657bd59525b1c5c0d5c0c5b6c5939576d545e51214ec24a8a478344b541633f8e3d443ca13b843bfe3b1a3d8c3e5b40784268443346cb479848b5484448ca468144b541033ec7397535b530e72b7627f822a91ed81a10177c1353101f0d100a4a076904b3015bff0efd33fbf4f9edf877f8aaf8fff8b8f9e3faeafbf3fc0ffebffe27ff66ff23ff87febbfd7efcf8fa48f940f7fff49bf2f6ef2fed69eab0e732e50ee355e12fe0a8dfd5dfcce069e296e442e729ea21ed14f0c1f209f5ebf644f810f96ff96df926f9bef84df8f4f7b2f783f788f7acf7cef704f82cf81bf8faf7b8f72af799f60df65bf5ccf476f430f444f4c6f478f592f61ff8cff9c4fbfbfd15002402180491059e062f07ec06010676040a0205ff9cfbb4f7acf3c4efe8eb79e8ade550e39de1abe018e0fadf4ee09ae0eee054e161e12fe1ebe041e05adf85de8bdd9bdc00dc7adb18db07dbfddafada17db03dbb8da41da5ad91ad897d6a3d47dd249d0decd94cb91c9a1c725c64ac5ccc4f7c4ebc54ac747c9e9cbc5cefed181d5d8d82bdc68df25e29ae4bee63ce869e94eea9feabeeab4ea32ea94e9d8e8a4e75ee606e545e38fe1f9df36dedadc0cdc6fdb78db40dc4addecde24e158e3bee545e84eea11ec8fed45ee98eeb1ee28ee70edbbeca7eba1eac0e981e83fe703e639e445e245e0c1dd3adbefd872d64ed4ccd277d1b9d0c4d004d1a8d1b9d296d367d441d59dd5a7d593d50dd541d471d373d25ad14cd03ccf20cee3cc8dcb20ca68c895c6dac4f4c219c1a3bf43be11bd58bcbdbb36bbf2ba98ba32baedb99db9a9b97aba13bc17bff4c390ca64d375de15eb3bf94a08ef16d22425318b3a0a4177442144ea408c3b0b34e32b3224191dd81712154414f115ff193d1fbd25362d22340c3afb3ef242c646aa4a884e1a535258d75d0f64696a4770eb757a7a4d7dfa7ef67eec7cf5791f7675713b6db069da6688659065a066e3689e6b516ef070aa7248731473ac716f6f0c6d686a2968f2666e660267ce68e26a3c6da76ff57021712770256d7b689e623d5b1053bc4a1f42f7399a32a92b95254e20291b7516fa11180d4e08a203befe6afacff6a7f3b6f1fbf0e0f0d5f186f302f56df664f7fdf670f5bff270eefee8d5e2f7db00d569ce42c8e9c27cbecebae4b784b55db364b16eaf61ad6aaba8a954a8cea753a827aa88ad68b2a2b806c030c89dd0c0d82ae060e6f0ead4ed0fef84eeafec1aeadce68be3c8e087de23ddf5dc92dd02df64e116e40ce77deadced37f1fbf4daf8f7fcc80101079d0cd5124419b11f0326c62bd830163528383a3a6a3b9a3b453bce3a273ac239ee396e3a563baf3c143e513f38407540ea3f893e573c8b39623630335730252ef22ce32cdb2dd72f94328c357b38f53a5d3c9a3c8b3be538fd342630762a8024b61e3019631477102a0d9f0ab008df063205860378013cffe3fc4ffaf1f7faf554f467f343f39cf394f4fbf555f7a1f8a4f9eef997f995f8c2f667f4b0f1afeebcebf3e857e618e423e262e0e2de6dddeadb6fdadfd853d70bd60ed590d4d8d4d1d58ed71bda25dd85e00fe450e70bea13ec20ed3ced76ecd6eabae861e6efe3d0e131e011dfafdeefde84df83e0aee1a5e28ce345e496e4d8e423e560e501e62be7aae8bdea59ed11f0e9f2b9f50ff8eff940fbc3fbbdfb49fb56fa59f982f8abf732f721f714f734f771f747f7cbf602f68ef4a7f283f0feed86eb6ce98fe74ee6e4e500e6bee620e8a7e943ebdbecf7ed99eecdee4fee50ed0bec63eaa8e818e796e55ee492e3eae274e233e2d9e16de1ede027e04bdf6ede6fdd9cdc13dca6db9adb00dc7ddc38dd32de00dfcedfade045e1dfe1ade264e350e498e5dbe652e804ea66eb9bec97edbded44ed4eec68ea00e86fe56ee289df1cdddada41d989d825d86dd872d97adab8db2bdd1adecbde63df51dff7de8fdea3dd9cdcc0db8eda60d966d808d7a2d55dd4acd2f2d05fcf7dcdc8cb76ca1ac92ec8dac793c7afc738c88ac8e2c84ac92ac9c0c82fc80ec7aac540c493c2f6c093bf3ebe2fbd58bc88bbedba52ba85b9c8b8dcb798b64eb5d1b30fb26cb0c7ae1cadccabc3aa25aa55aa46ab4aadbab065b598bb82c39ccc01d781e21feeb3f9d404560e2f16251c501f3020261fdc1b6f17c012c40dab0936071306ff06240aa40eb314f41b3e23b12afd314338fc3d2e437647a44bdf4fe7537c587b5d6662a867bb6ce9708d742377257824781177ed743172956ed96a8d6886678e673469df6b1e6f0d73d676157aec7caa7e517f547f5a7ecd7c467b7879d477bb768a7574749b731972f76f486d50695464ab5ef357c550a6496942bd3bf135a430552cfe28f1257a236321ea1e771c021af716f41323110c0e5b0b37090e075d051f049002f60039ff98fc5df9a3f5eef0abeb2de63ee05bdaded4a8cf18cb54c71cc4a6c1ebbf87be93bd0cbd9fbc71bcabbc18bdd7bd23bfd2c0e8c298c5b0c8fbcb89cf0ed32fd606d962dbe4dccadd25deb7ddefdc1ddc10db43da21da72da8cdbbbdda1e063e41de94dee02f43bfa6900a906fb0cd4127118e91db62221275b2be92e1032fc343437f0384d3ade3ae93a823a5839d63738365434c332db31883151327734c737763c5442e148f04fe856235d6a622b6607682e6879660a638c5e2b595153b94d7c48e14357408b3d5d3be2398038ff3673356f330731912edf2b4f295927d52521257a255d26dd27f129c22b2f2d252ede2d692c072a5a26c821e41c9e177912000e150a0307ef04710391023102c2014401a9009bff57fefefc78fb2dfa3bf981f84ff897f8fff8a5f956fa9efa93fa1afaf1f84af746f5eaf282f035ee1cec6dea1be915e858e7a5e6e4e504e5c7e349e2b1e0e8de47dd28dc7cdb89db93dc59dedbe00be467e7bfeae2ed53f005f2f1f2d5f2f6f18ef094ee7aec7eea82e8e3e6b9e5a8e4dee351e388e2afe1d2e091df44de24ddf8db2cdbfcda13dbbedb1bdda8de80e09ee269e4f3e53ce7c9e7cde76ce75ae6fbe48be3c0e103e089deecdc76db3ddabfd83bd7cad5f9d31ed273d0b0ce49cd83cc11cc61cc9acd39cf71d135d4d5d65dd9afdb2cddfadd27de54ddecdb33dafad7d2d502d44bd225d1abd061d093d031d1a3d12ad2c7d2f9d224d36bd36cd39fd330d4afd484d5c3d6dfd725d991da84db4edcf0dcd9dc7ddc01dcebdac5d9c5d874d756d68cd57dd49bd3fdd2fdd110d151d022cf17ce67cd70ccc8cbaccb71cb8ecb22cc67ccc0cc3ccd11cda1cc10ccb0ca04c953c717c5e9c217c127bfa5bdc4bce4bb72bb7dbb4abb2abb2abba4baeeb933b90cb8ddb6d9b5c4b4efb35cb3dab2a5b27fb230b203b2adb1feb067b0b3afd1ae40aecfad72ad8badccad22aeceae79af46b089b109b340b5afb827bd33c33acbaed4b9df35ecf8f8b505d511e81bc0231729f72afb29bb2610215c1ad3139f0d1d093907a507030b481150190723c02d0d38e541d34ada51ad57795ca15f11628c641c67756a6a6e6072a8768d7a117d657ee67d0f7be576aa717c6bbb65f060495dae5b135c225e0162f2664f6cef71e876c97ab67d1a7f1a7f527e887c347a0a78b1757a73c671cd6f926d326bc9676763595e16581951074aba42e83b26363031882d3e2b8e29a02823280e2792258d233e20351cc817a812b60d6b098005a402f500c1ff3fff33ffa3fe93fdd7fbbcf892f49eefbbe992e3b5dd39d8b5d377d049ce4acd53cdd0cd97ce60cfa5cf5bcf99ce4bcdc0cb65ca6cc92ac9f3c9c1cb84ce3bd27bd6d0da0fdfc2e278e555e74de835e89de7e5e607e699e5f6e5d8e67de8f4eaaaed9cf0b6f36df6edf863fb7ffda9ff44022005a008050deb115d17341dcb220828b42c4930ef32b9348135d7351536443603378b38a43a8b3d1241a1441a481a4b094de74d934dec4b5449204699424d3f923cb03af339323a593b503d853fab419343a944d9444244aa425a40b63db63abd371c359c326e30982e982c722a22282b25ae21db1d86191e150a11490d550a78087c078f079508ff09bc0b800da60e2f0f070fcf0dd60b5d09590649037f00e7fdcffb46faf9f8f4f712f7e5f573f4b2f26bf0d9ed36eb95e84ce699e496e373e31ee471e55fe78ee9adeba3ed23ef06f067f02ef078ef93ee86ed86ecd4eb57eb24eb4aeb78ebaaebe6ebd6eb96eb48ebb3ea1ceacee990e9ace961ea4eeb94ec49eedeef5cf1d0f2b3f325f456f4e5f328f378f288f1b8f063f01af018f094f0f3f044f1b5f1b8f161f1f3f01cf01eef3fee50edbbec83ec8aec02edbbed73ee19efa0ef8eef03ef1aee79ec6fea4be8dae581e38fe1bcdf43de45dd5bdc92dbebdafbd9e6d8c3d753d6e6d4b1d392d2ebd1e3d141d242d3d7d48bd66ad848daa2db8fdcf7dc8ddcabdb72dac2d821d7bad560d486d334d306d33dd3bad306d465d4bad49fd488d487d45ad4a1d47ad588d649d8b5da2adde6dface2b3e435e60be79be66de5a5e3ece011de68dba3d889d65bd58cd49ad47fd568d69ed705d9c8d943da89da08da5cd9dcd81cd8c1d705d853d814d94ada29dbe6db6adcf3dbcdda1bd96dd65ad34bd00fcd4aca58c800c7a7c64bc760c8f6c9cbcb43cd6cce18cff8ce64ce70cd18ccdecae0c914c9c1c8b9c8ccc804c9f4c866c866c795c512c34cc023bd06ba9fb7d0b5f9b47fb5efb652b9a4bc10c094c325c702ca89cc2dcf8fd16fd48dd89ddd35e4a8ec1af67300440b1a15831dea231b274727ae241b1fd21707103e0809028afee9fde6008107ce10751c6d293a365342d74cdb54a15a285e7f5fa75f185f3b5efb5d4b5e175faa60466264632564d6633762d35fa55c2a59ff55f7521451a3512e5479588c5e4f65426c0f737678507cb67ee17e557dc87adf7667722a6eb0697565d361ed5dea59da55dd50554b97452d3fea387933a22e452bcf29a3291a2bf92d0c312a34c636a537cf361d34fe2e2b282220fa16db0d5f0588fd32f779f2d0ee7fec2febfae9f1e8f4e74ee65de45fe207e0f7dd6fdc42dbcbdaf5da52dbdedb3ddce4dbd5daedd801d66cd283ce87ca02c75cc4cfc294c2b3c3f4c51ac9cfcca6d03cd45dd7e3d9b0dbfcdc0bdeffde2be0d8e1f8e39ee6c8e90eed40f030f369f5dcf695f76bf7b4f6dbf5eff479f4fcf473f622f933fd3a0207085c0e8914461a541f3723fa25ba27582849280528a927bd27a728632a2b2dfd306c35403a173f5a43be46e04872498f483a469442303e8139fb343f31a62e6e2dd42db22fd432f236663bb33f7043f8450c4799466644b540f33b4b3643305f2ad0240020241c15190217d3151115bc14ab1474143214e6135b13cd124b12a9111c119d10ef0f320f450ee90c3d0b3709b906f4030001d3fdbafabff7d2f430f2c9ef7bed76eba0e9dee779e66de5bbe4c1e47ce5e0e623e910ec52efd8f22ef6d4f8a9fa45fb60fa22f882f4a7ef1dea30e445de07d9c2d4aed11dd0f3cf04d145d355d6ded9c6ddaee166e5f8e830ec02ef91f1b0f34cf56ff6dbf677f653f546f362f0deecc1e857e4ffdfe7db77d8ffd57dd41ed4edd49dd622d952dcbbdf4ae3dfe61bea13edd8ef2ef238f4fff53af7fbf730f87bf7edf583f301f0b4ebd6e673e11fdc49d710d300d062ce11ce43cfdfd157d58cd924de61e21de628e90cebeaebe9ebe3ea39e93be7e6e49ce293e09edeeedc87db1ddad0d89bd73bd6e9d4bad388d2b4d16ed18bd159d2efd3f1d577d876db70de67e142e495e67ae8f4e9bbea16eb1deb9aeadde900e9c5e77ae632e5aae335e2eee0a3dfb9de48de1bde9adecddf4ee16ae309e68be810eb77ed1aef1df086f0e3ef91eed4ec73eaece79de558e389e167e09fdf68dfb7df0ae087e018e138e122e1dfe013e025df42de2add54dceddba3dbc8db67dcfedcb0dd75ded6deeedec7de18de17dde5db6ddaf8d8a0d75fd66dd5b3d41dd4d3d38fd334d3efd27ed2d8d14cd1b4d016d0cacfaecfd0cf5cd018d108d233d34bd485d503d788d882da3edd8ee0f5e4a4ea30f1d6f85b01ce0903126e19ef1e7a22d1235e22c91ea21922139e0c1307f3027601030348079f0e661862234c2f163b6945454e20555c59bf5b875cbb5b7d5a2859bb57fc56b8568556c756f25685560f564d551c545b531a5376532555d157635b6c6044663c6c47727f77697b2c7e3a7f9c7ee17cd379df75b6711d6d74682f64c55f615b4957e1526c4e5a4a4446a34200400f3e423ddc3d3d3f6e4127446146f0476348c2463943d13d31363c2d8e234019770fd70646ff84f9b8f53ef345f27ff200f3caf3a0f4dbf4bbf448f433f3e4f173f097eea3ec85ead1e7b2e405e170dc49d7c3d1d9cb1bc601c1adbc90b906b8fdb774b95bbc4dc0e4c4d3c9abce10d3e6d60fda73dc45dea6df95e050e1efe13ce257e23ce2a2e1b1e090df1bdebcdcdfdb85db37dc61ded4e1c4e640edacf4d9fc8a05eb0db415ba1c6622ba26e129a52b532c442c6e2b262ab028f7264925d02365225921de20d72095215223f2259c294a2ea4337639663ff544c8497b4dc74f9150bf4f7c4d174abf45f040203c75374f33ef2f292d132ba229682860277c265c251b24d2224e21d71f9c1e741da11c2c1ccd1baa1b981b2e1b8f1a9419d4179815df12600f870b81071703b8fe97fa85f6dcf2d0ef3bed61eb55eae8e942ea51ebc8ecaaeebaf098f22df423f528f548f459f24def7ceb12e74be2b3dd99d93bd6f9d3eed217d374d4c9d6d0d939dd9ee0c3e367e64ce884e912eae0e934e934e8d2e65fe502e49ae25de161e07cdfe1dea5dea7de20df1ae069e130e357e59be719ea9fecdaeeeef0b1f2d7f3a6f423f516f5def499f414f4a6f35ef3f0f294f24df2c5f12ff197f0bbefe2ee2cee6aedf2ececec1cedbdedd1eef2ef3af192f281f321f46df4fef306f3a8f1a9ef5fed14eb97e836e62ee43ce293e05ddf55dea9dd7edd88ddecddcbdecfdf0de18fe2eee326e52de69ce67ee6e0e57ee496e266e0d4dd32dbd1d89fd6e0d4bad3ffd2d4d23dd3edd303d578d6fbd7b1d99ddb75dd63df63e122e3c6e446e651e70de877e84fe8d0e708e7cee58be45be316e228e1aae057e07ee01de1dbe1f3e24ee483e5dbe64ee878e9aceaf3ebf5ec0fee4aef2ff00bf1ddf11af2f7f175f11cf03aeef2ebf9e8c7e5aee28edfeedc18dbd6d996d963dabbdbc8dd67e0e9e25ce5a3e727e910ea6beadee9b7e82ce70ae5a9e240e0a4dd27dbf8d8eed646d514d42cd3afd295d2b3d214d382d3c9d3eed3afd3f6d2fad1a5d012cfa1cd60cc86cb6acb07cc79cdbbcf70d297d502d930dc39df23e2a0e42ee720ea53ed53f158f6ebfb2b02c508ba0ed913a9174219e018ab168d12960daa084704c701d4015804dc09ff119d1b67265b31033b204330498d4ce64d9e4de34bdd490c488346fc455f463447ac483a4a4f4b384cb24cb14cff4cb04dec4e73511d55af59555f5b65256b8370a0740f77ea77da7629747670d66bf6667f624c5ec65a2f58e255ea533c521350994dfc4ad047a344fd41bd3f743e5f3ef93e584010421c4356432642a93e3339cf315628f31d6113df08b3ff72f8f2f2c4efb7eeefee4ff037f2b7f3c6f409f50df444f2bcef5decc3e801e5f4e0f9dcdcd841d46fcf4ecab8c434bf07ba59b5c6b1a6af0caf2eb000b321b722bc7ec1a5c60acb50ce52d0fbd072d01bcf46cd62cbe7c901c9dac87cc995ca0bccb1cd0ecf3bd062d152d281d36ad5f1d78edb97e080e636ed97f4bafb450201082e0cc70e0410b90f800e050d720b8d0ae70a5b0c510fe5137c191a208927f42e37361c3dfd42ed47e74b874e0d509d500050984eaa4c304a8d47f644794278400f3f513e923eb13f82411c4422473b4a554d0050f0510f530a53db51aa4f654c65480044243f333a8135e630b82c2b29ec2530231121331fca1dee1c3b1ce31be71bd81bdf1beb1b831bce1aab19ad1720150b12260ef309a5051201c4fcf4f876f5b7f2cef061efa1ee7bee89eee4ee68efbceff6eff5ef77efa3ee6cedb7ebbfe974e7cfe419e255df96dc32da33d8a6d6c5d580d5ced5bbd613d8aed96fdb13dd87debbdf8be01be178e18be18ce187e152e11fe1e8e070e0dfdf2ddf27de1cdd20dc1fdb80da60daa3daa6db6add9edf6de2ace5e8e838ec73ef36f2a8f4aef6f5f7b8f8f4f873f88af746f67cf48ef291f062ee79ecf9eabde929e941e9b3e9b8ea38ecc5ed84ef56f1bbf2d8f3b6f4e0f494f4ebf397f2eaf005efc1ec6eea49e846e6aae4a0e30fe321e3d0e3cee418e67de78ae83ee985e90be905e89de6abe486e283e08adee3dcc5dbefda7ada78da95dad6da47dba5db05dc71dcc2dc2bddbcdd47de00dfdfdf9de06ce147e2dde268e3e7e3ffe3e9e3ade3fee225e245e121e000df0ede22dd87dc5ddc75dc04ddfadd12df78e0f8e139e370e46ae5c6e5dde5a9e5dde4ebe3f1e2a4e175e08ddfa8de1bde02de11de73de1ddfc0df92e072e11de2e7e2ade322e4c0e47fe5fce59ae64be78ee79fe779e7b4e69be54ee49ee2eae061dffadd0edda1dc86dcdddc64ddcfdd26de1cde92ddbedc72dbc8d930d89ad629d544d4cad3bbd345d417d553d6e7d76cd938db25ddc7de90e089e245e45de611e903ecd3efbff446fab500d007a00eff144b1a781da51e9c1d071afc14300f2909b104a9023c038707550f6e19a425b732b63e33494351ba55335702563a525e4d4b484e43a03f763d6a3cff3cbe3edd40b943e046c549214dca506054a4585b5de6619f66046b4d6ea770af710e71536f826cdf685165f261185f815dd95c015d315ea05fdb60ec6112622a619b5f1f5d105a23573e54d3515750534fda4ed34e464e044dd64ad64640416a3a0c3206292a2081170410590a2906da036803e9033f0509074308ed08df0875071305ed01aafdd8f8bbf306ee2ee860e252dc77d612d107ccdfc7e6c415c3c9c21cc4cec6b7ca8ecfa1d478d99ddd79e0c3e15fe139df8fdbe0d69cd155cccdc77fc4a4c295c251c469c7b1cbced0fed5f8da8fdf50e35be6efe8f6eadbecebeee2f0fbf248f541f703f9a9fac9fbbafcebfd47ff5f01b50408098c0e33151c1cf7226729792e02320f34583473332532bc301130c230bd323b36133b7540f745094bd44e1c51b7518e50304e104b8f47704413429c405f403d41ed424245b847fc49e44bfd4c4b4df34ca74b99490747a943cb3fb23b22377a32082e9529a2258a221320a11e461e741e3f1f65202d2191213f21951fca1ccd186a13580df506620084fabaf5fbf1caef1cef85ef00f1fff2c1f415f67ef694f573f31ff093eb71e60ae191dbc9d6e4d2ffcf72ce0ece9fce21d036d295d410d731d9d1dad9dbf2db2fdbafd945d729d4aad0cfcc08c9c9c531c3a0c15cc147c279c4cfc7dccb6cd00dd51ed970dcb3de8cdf3edfefdda9db08d974d61bd48fd20bd275d20ad495d6aed965dd5de10ee58ce892ebb9ed4fef48f06df035f0a4ef89ee62ed41ec09eb47ea08ea1aeae0ea4becffed2ff099f2b5f49df604f867f805f8edf6f1f49ff249f0dfede9ebb3ea11ea4dea76eb18ed20ef52f11df36ff41cf5baf479f37af195ee3eebe0e772e469e125df74dd8bdc93dc28dd39deb8df2be179e28fe317e436e4fee32ae3fde1ace0f7de2add8ddbded94dd804d7cad5ded46ad439d48dd485d5d2d69fd8e4da37dda9df08e2bbe3cce426e569e4e5e2d2e016de34db8ed828d691d413d47cd406d688d862db81de86e1c5e34de5f9e55ee5eae3dfe12edf8bdc61da90d88ed774d7d5d7ded876da1bdcf3dde2df7ae107e38fe4b6e5dde608e8c7e862e9d0e9a2e92ae976e836e7d2e573e4e2e289e18ce0b8df5fdf77df9fdfffdf80e0d4e020e150e12ee1e6e06be0b1dff0defcddc0dc7adb0ada6dd800d7d7d504d5c4d423d53cd609d844dae7dca1dfdce1a8e309e5c6e57de6c6e7c7e936ed79f242f98601a70a5e13d71af01f7a216e1fe71952116f07c4fda6f532f17af18df6c700240f8f1fa1305e40a04cb9541858805633514d49e33feb36782f0d2a8f27a6279829662d3b326037323d45434549d94faf56545d1e64666a546fd172337426733470846bd0654b60415b6b57c055e355c257875b0c608c64d368e46b746dd26db36c716aac675264f860255e8b5b785901586156ba540a539250954d384ad545d740a63be93541301d2b2d26e8217f1e8c1b81194a184b17cc1679168d154e149512cc0f600c3e08ec02fdfca8f6caef29e913e35fdd99d8ead425d2b1d084d036d1cbd2cfd4a9d64dd85fd96fd98ed88fd641d3fbce06cab4c4a5bf4cbbf3b7f8b593b5c3b676b981bd70c299c785ccd0d0f0d3d0d5a2d64cd618d593d3f4d1b9d062d0e5d063d2d2d4a1d7cbda49de92e1dce46ae8d6eb85effbf3e2f879fef404860be611e317a41c07202922aa22fc21b520f71ea61d871d921e4021b125272b6a312838753e04449748a14b464db64df24c804bb34991478345ac430442d7402d40fa3f6b405941ae427c446b463d48cd49904a4d4afe486946de42c73e3e3ade352632142f162d4f2c412cde2cc52d282efd2d032da92a57274123411e0619f313f90ebd0a7807e00441036e02de01bc01c0016201d500d3ffdafd34fbcbf766f38fee68e9eee3bede06daded5dbd214d176d038d103d36dd554d81edb4fddc1dee7de82ddcbdab7d696d117cc9ac6a8c1d8bd58bb6fba35bb48bd83c088c49ec888ccfbcf70d2f8d395d412d4cbd2f1d081ceffcbaac988c724c6b1c525c6ebc7edcad1cea5d3e6d8e3dd85e243e685e88ce93ee983e719e55de288df69dd42dc08dc27dd74df88e287e60deb8bef13f43af879fbfefd89ffc0ff02ff4dfd83fa49f7f0f399f002ee77ecdfeb8cec63eedff0f0f335f708fa50fcccfd1cfe80fd1ffce8f94df793f4abf1ffeed5ec15eb0eeae9e967ea9aeb7ceda4eff1f12af4c3f58cf669f615f5c4f2d2ef5cecd5e8b8e526e36ce1cae017e13be20ae413e61fe804ea78eb82ec2ded4bedfcec62ec61eb29eae6e881e71fe6e4e4c1e3e9e286e28ee223e33ce49ee547e703e97ceab5eb7eec81ece8ebbaead8e8a7e670e434e265e045dfc5de2bdf79e05ce2d0e48de70eea4bec0beef0ee32efdbeec4ed64ecf9ea76e94be891e7fbe6b2e69fe664e62ee6ffe59ae540e502e5bae4bee427e5bde59fe6a8e76fe8f0e80fe9a5e8e5e7cee662e5f3e37fe20ee100e044dfabde5dde3dde21de30de7dde16dfffdf0de14ae298e38de446e5d2e5d9e5b2e5ede5ace692e83eec98f198f8cd002609d010b0168619fb18d714300d880370f950f068ea24e9c8ecc2f552038713dc243d354842f44a734e704c3946173d4e320d28951f71199f16f816ac199e1ee924902ba932b5393940c246f34c3252c456185a775b265bf358e254e54f7a4a6845fc4180403e41af44fe4961508457215e566304677f68b46743654c61785cb3572053454f9f4cd84a1f4a934a8a4bf24c994e924fc14f094fbf4c2a498e44ad3e29389531042b5225f720c31d1d1cd71b2e1c291d531eda1ed61ef01d891b09187d13ac0d5707cd0002faaff316ee21e963e5e7e262e10fe19ae16fe290e392e4ebe4b7e4c1e3b4e1d3de2fdbbbd6e2d1f5cc22c8dcc37cc033be45bddbbde0bf23c350c7dbcb23d0a5d3ecd59ed6c7d58ed32ad048cc8bc84cc544c3e4c203c4c9c634cbafd01ed761decfe543ed87f4e6fa3e006104a30620070006140324ff17fb5cf71af538f5c3f72efd6905760fc61a7626fd30a839ec3f104360435c414f3d3938f8320e2e722aad28cb28202b782f3835273cae43004bbf514a57f85aab5c395caf599c556d50af4a19450b40fd3b583909382838a339e03b9f3eac416944a9464c48ce480e48ef452742043dcf36b52f8828d521db1b6c17d814e313ba14eb167919f91bb51dd31d5e1c3f196014790efb072e01f4faa3f544f142ee69ec50eb12eb4aeb87ebf2eb33ece1eb2bebd1e991e7b9e437e10addaad834d4f5cf7dccd2c910c881c7e3c7ffc8c8cac6cca8ce4dd049d182d108d1b7cfcecd9ccb2ec9e4c618c5d9c37bc322c49dc5f8c7f2ca0cce2cd1fdd310d67fd734d811d88dd7dcd614d6c8d50fd6c3d630d82ada53dce1dea0e13ce4f4e6a3e901ec52ee67f0f0f11ff3bdf37ff3c7f2a5f120f0eaee4eee5dee9def0ff252f56ef9f0fd1202a1052c081f09aa08f6060b04920011fdb7f913f76ef5a4f4e3f411f6b3f7b1f9cffb88fde3fedcff1b00c6fffafe67fd35fba0f880f519f2c8ee81eb90e858e6cde42ae4a1e4dde5bfe70fea2decdbedf1eef4eeefed17ec46e9dbe55fe2ecdef5dbe7d99ed833d8b2d8b2d921dbeadc97de16e04fe1d7e1c6e13ae1f6df47de67dc2cdafbd724d693d4b5d3c0d363d4b7d59ed790d98adb66ddabde75dfbbdf32df41de2addd1dbb2dafad966d944d9a8d94ada75db28ddfade0ee141e321e5d9e64ce80fe94fe901e9eae77fe607e583e373e2f4e1d5e156e260e39de428e6c5e7fee8eae971ea65ea17ea9be9dbe813e843e762e6b9e544e5fde419e55ce599e506e67ee6e0e661e7f1e775e809e9ade978ea6feb4fec09ed75ed23ed36ec05ebabe9c1e805e9c4ea70ee41f4cffb9404840d1c15421adc1b19197312c10829fddbf1d0e874e363e327e909f41f03751467250e34913e8f433143ee3da6347329031ea413240c3908af079b0a341045176b1fd827c32f4737ee3d2a434e47024acf4a224ae347e943043fae39703480306d2e892e58315c36e53c9b445c4c24539e580a5c015ded5bec5874546f4f3e4a634581419c3eeb3cb03c913d7b3f4b4243450e485b4a604be94adf48d644233f39385a307a2865216f1b58175515fd145b16ea18a41b321eed1fec1f401eec1acb159b0fdb08b80105fb20f50ff05becf8e977e8fae725e85fe8cee83ee92fe9c8e8f1e746e600e439e1d9dd2bda4fd648d275ce1dcb6dc8d3c682c656c73fc902cc29cf4dd212d5fbd69fd7dfd6b7d45fd17bcdacc973c680c42fc468c554c8d4cc3cd231d84fdec9e363e825ece0eef3f0aaf2e2f3e4f4c1f516f632f645f605f6f2f58bf6d2f792fa73ff4e064b0f101a4f2520307239db3fd34218427b3df135b72c0b23ea1ad11577149417ec1e5a29e7351f43444f3559e75fae62cc61aa5d0857354f0c47483fcd38f633f73015301b31df332a385a3d23433849bc4e30532256ab567d54b24f58482f3f2535012b03220d1b8b1639150717111bd3203027972c6530ef3185307a2c1526941d14146a0a330192f9e2f30cf05fee65ee77ef9df136f46ef630f8e6f8f3f798f5d1f1a5ecaee61be034d9bdd202cd6cc8b5c5c8c472c5b9c7faca93ce3cd245d51fd78ad727d60dd3acce60c9e9c308bf10bb86b8bcb78db8fdbac2be2dc3d9c738ccb2cf35d29cd3d0d331d3d6d1dccfdecd0ecc8bcaeec944ca75cbdfcd58d19fd5d8da84e012e668ebdaefe6f2c3f43cf548f499f26bf008ee50ec89ebd4eba0ed9cf04ff4b2f834fd550133057708ce0a7b0c5f0d620df70c240cd30a6509d8071906ab04cf0391035204120680088b0be70e1412e514fb16d6176e17c215ca12030fe50aa306b70280ff03fd83fb32fbd9fb5cfd90ffe7010904c1059a0671064b05ff02bbffe6fbaef790f31bf060ed8bebc5eab6ea2beb0fecf5ecabed24ee13ee8aedb8ec7deb0aea9ae8eee618e54ee368e198df2cde07dd4bdc1cdc37dca2dc52ddd8dd1bdef8dd12ddaadb0eda37d8a2d6a3d5fbd4dcd465d535d64ad794d893d93fda9ada7cda48da31da01dafad915daf1d9ddd9d8d9aed9dcd976da22db15dc55dd82debbdfcce022e1d4e0ebdf4ede96dc29db0bdaaed926da2ddbecdc39df9fe10ce426e687e75fe89be82de880e786e60ae560e393e1a6df14de2bdd19dd1ade17e006e3bde697ea39ee5cf150f30bf412f4b0f3a6f3dff4b2f750fc70022809a70fbc140d172f16ee11750a5a015bf805f16eedc2eefbf4f2ff640e211e632d003af541b9440f42793a083076244619a210800bfa098d0c9d12ee1ae3243b2fc3385b416c48934d60517b53825314521c4f904a7e456240ac3b74381c37f937ab3bb2416a496a52385b9f624368446b576b1d69c464e95eac5897526f4d084a50485d48274ade4c2f50d853ee563359815a145ae7572f54b44e0248b640f6389131242bcc254322bd20bd205a220f25b627072a7e2b362b43299725e81fea182511dc081e0171fadbf4f2f0b4eea9edf6ed30ef87f0d4f185f2f2f156f0b0edd9e959e56ae012dbe6d538d125cd17ca14c8e4c696c609c712c8bdc9cccbe4cdc1cf08d16ed1e1d05dcff3ccc7c91ac64fc2d5be4bbc4bbb04bc90beddc25bc89ece49d596db0fe169e514e813e9c4e847e744e572e3eae126e1a1e12ce30be67beafcef7bf6d6fd41058b0c9213a1199f1e6e226924be24cd238c21b91e141ccd199918fb18dd1a951e0f24872aa031af38af3e5e43784698471e47544566421c3f0a3c94394f3848384e394f3bc83d5340d042c84402468a462e460e459243cb41f63f4d3e923cd23a2a396f37e035963443331d32383149308e2f0d2f472e2f2d842bca2844252621741cca1764133d0feb0b8809d8071207d1066206b1055b04010205ff74fb52f73bf354efa1eba8e861e698e46ee37be25be124e096de9cdc94da6dd82dd62ad440d273d00ccfd0cdc6cc0acc49cb8eca09ca96c95ac97ac9aec9e9c928ca22cae0c967c987c877c75ac619c515c494c388c32ac476c524c743c9a9cb06ce6fd0a7d25bd4bed5ced672d70bd8a7d830d9f4d9dedac2dbeedc50debadf69e13ae3fbe4f1e608e91ceb5fed8eef5cf1f4f22bf4ddf45ff59ff585f563f535f5fcf425f5a4f551f667f7b4f8f4f94cfb95fca0fd9bfe59ffafffd2ffb6ff57ff01ffa2fe1bfea8fd2ffd94fc23fcd5fb8afb72fb78fb70fb81fb9efb99fb88fb50fbc6fa0bfa18f9e9f7c3f6aff590f493f3b2f2c6f1fff069f0e1ef89ef56ef09efadee43ee98edb1ec87ebfce92fe83fe63de48ce259e192e070e0f9e0d1e1f3e24be44fe5c2e5c5e5d9e42ce341e1eadeaedcf3daa1d9f5d813d9b9d9e5da68dcc3dde9dec1df04e0eddf91dfbfdebfdda1dc44db18da47d9afd89fd805d98cd974daa3dbbddce7dde7de5ddf83df49df95dedfdd35dd80dc1adcdddba4dbcfdb36dca9dc74dd4fdef8decbdfa8e079e18ee2a2e380e447e593e55be5f4e40de4b1e258e1dadf6bdeabdda3dd7cde75e01fe345e6abe996ecd6ee54f077f06aefaced69eb80e9f1e822ea9fed7ff30afbaa033b0c1f136b174018ed141b0ee504b0fac9f10dec9cea86eeacf7d9049f14b424b832153d37427a41cc3b46328e261d1baf11970b0e0a040dd913ce1d3929a8342a3f6e470e4d6c5062515a502b4ecd4a98466342763e1e3b15397938af39283d73427649be51ef594361fb66f0690c6a9667a2623a5c6b55c74e6949ff45834459453948224cbb505255e758725bb25c245c345afe564052964c6346c93f8b39dd33b32ecb2a3c28c126e1266128632ac32cdb2eb22f3d2f312d2a29b8231f1d9d155b0eea077e02e1fef5fc14fc4afcfbfc44fd34fd66fc3efa1bf725f364eea3e932e514e1cbdd42db34d9f6d744d7aed65ed603d63bd563d491d3b8d234d2f9d1bfd18bd128d16ed079cf17ce37cc2fca34c892c6dbc56ac654c879cb88cf0dd46ed832dc29dfffe080e1e1e074dfc8dd8bdc31dc1fdd4ddf1fe23ee54ee8b0ea70ecd7edcceedbefd7f119f53bfa8d015c0ab413901c6023202783274224271e5916f90df8060503ef0273075010021c2d2941367741e149d14ed24f664d36481c41b5392433fd2df22a022abc2a122db03034357d3a01404945264afa4d5c5041513150e84ca147924082389e30ca290e250b239823a626ce2bf9316a38373e044239439641fa3c3636342e95256c1d6716c110340de30b4b0c340ece100713a6145315b5144f133a11380ea00a7a06bb01f3fc42f899f35aef6debd2e73fe5eee3cae3ece4bae665e8a6e902ea33e95ee758e41fe034dbf4d508d150cd1acb7eca75cb60cdb4cf21d228d480d5fcd565d5f5d310d209d07ccec1cdb0cd2dceeace7dcfebcf37d05cd0a9d02bd1d8d1f8d299d4b5d672d961dcf0de0fe18ce24ee3bde3f1e3f5e328e48ce42fe584e67be8d9ea9aed42f070f261f419f6a0f760f946fb20fd0effd50036023f039503e1025b0130ffd0fc24fba7fa88fbf8fd8f01a905f609ef0df010b412f1127811b10e310b8e0778044802fb009400eb00cb01430329050c07bf08240afe0a770bd90bf70ba20bb20ac608d2051702c4fd55f962f525f2fcef56ef2cf07bf21df63efa1afe1e017f020302ebff33fc35f78cf170eb7ee58ee0eddcf1dacedaf1dbfeddbee087e314e642e86fe97ee9a2e8c7e669e40fe296df31ddf9da7ed802d6f3d327d2f0d09ad0d5d0cad1a3d3f1d599d835dbdfdc6dddd0dcc8dafbd7fad4d0d11ccf3ecd0dccf0cbffccacced6d00ed394d479d5c6d54ed588d49bd352d20ad1e0cfcdce4ace55cea1ce5ccf50d03cd183d217d4b3d57ad717d914da92da9dda55da1bdaebd9d0d9f1d9fbd901da56dab6da29db24dca8dd0ce003e4b9e928f1d4f98702290a8c0f70119d0f3e0a900100f768ec64e317de26dee7e338efe7feb910b1228132d73da1434443bf3cbe3145245316a70a25037a003603d50ae6153b230c31783d9047494e08518650354d8f47fb40363a9c33492ed42a8329e62ad02ecd34973c21458d4d8355de5bbd5f1f61915f1e5bcf54644dc5452b3f153aff365f36e4375f3b7740f645154b514fb9512e5204510e4ea4494b44023e5137cb30902a39251c21fd1d371cd71b621cf51d44205522d4234d2407233720171cb416ca10c60ad504c3ffd1fbe4f860f7fef608f76cf7c0f770f79ff638f509f36ff084ed5cea7be7f7e4bde201e181dfe3dd41dc81da8fd8bad61ed5c5d3ead29dd2e0d2b5d3e0d424d644d7f3d702d862d71dd655d428d2dacfc5cd22cc54cbabcb0dcd6fcfbdd280d67cda8bde3fe27ae527e8e7e9d8ea2eebd0ea2beaa3e919e905e9e9e9b8ebd7ee86f340f9c9ffae06010d7a12cd165f195a1aed1903186c15f212e5102010181187139017fc1c13239229ee2f42354e39c13b4b3c6b3b8539da362f34ef314230b32f6130303233350539273d5d411a45f547eb49aa4a174a7b48e1459442243fcc3bf138e3368135f2343535dd35ec364a386039123a423a7539c4374635d831df2d9529ff24bc20181d021ae617a516b6153415d5140514e9124a11ac0e5c0b6607c9023afe01fa26f62bf3f8f04aef6cee0feeb7ed65ed94ecc9ea48e808e519e11ddd2ed95cd51bd262cf35cde9cb44cb0fcb4ccb9acbdccb41cc96cce2cc43cd64cd30cdb5ccbccb6fca07c970c7e6c596c470c3c7c2c2c23bc353c4ddc574c728c9d1ca3bccaecd13cf32d059d175d264d388d4ced5ffd656d8a2d9bbda06dc73ddf7def5e02ae360e5e8e780eaf4ec91ef0bf21ff417f6bdf7f0f80afad7fa2cfb55fb33fbdbfaddfa4cfb45fc29febd00c3035107f10a310e0311fe12da13d61306138a11d00ffa0d190c760a20092708d0071a08ed08590a310c280e2d100a125a13f613bc1371123210480de1095c0622035a003bfefefc90fcebfc05fe79fffe0068025303a7038b03df02b001320030fea7fbdcf8bff57bf27cefc7ec8aea1ce962e864e835e95dea8feba1ec09edacecbceb11eae1e781e5d1e20de08cdd2fdb35d9e6d702d7a0d6e5d66ed737d84bd93cda08dbb2dbe4dbc7db76dba7da98d96bd8d1d618d57ad3bdd13dd03bcf86ce68cefecef9cf73d142d3ead475d6abd723d81cd890d747d6bed430d394d183d03ed09bd0d6d1c6d3f6d55bd89bda5fdccadd9edeb7de87de06de36dda6dc5adc32dc7bdc23dd13de88df60e186e3f6e525e8d0e901eb5aeb00eb8bea26ea4deab8eb99ee25f357f97200bd07360e8b122814cc12490e9207efff72f8cef27bf014f212f80f02a40e601c56298333ed39d23bfe38af323a2af8201119f9133c126d141c1a15225f2b9034603c5d42e445ca46e2457943fa3f8f3c8c3901378f352d35b0356f37313ac93d50422547d64b4c50a75363559955c553e64fcc4ad744d43eea398a362f352f36f738223d3342f346bc4a324d8d4de94bd8487c448e3fca3a3c364c32262f712c592ad72869274f269525cd2448242024d0236123a122fa20801e2a1bd7161f12490d69083f04070199fe62fd35fd67fdd3fdf7fd23fd5cfb8ff8b9f479f028ec14e8ece4d0e2a2e17de1e0e122e20ce231e149dfacdca2d97fd6e3d331d298d132d2c6d3edd52ed8f8d9f1daebdad4d9e1d76cd5d4d286d0e3ce3eceb7ce2cd084d285d5bcd810dc73df8ce25ee5fce719eac3eb22edfbed69ee8aee33eeaded43edf5ec45ed6dee25f0acf205f6b1f9e6fdc202e207740d89139d19911ffd2400294c2b752b1129c024371f221907141311d8102414ff1a97242b30563c6a4759500756bb57c4557d509e48aa3fd1362d2f072ae627e728f92c4d33043b5343084b5951dd55da572a571854ad4e7e476f3f16376d2f53292a259223a724ce27b22c7932bb37cd3b053e9c3dcf3af3353d2f9d27c51f1e1894117b0cc108c5063606750694071009340a130b410b380a4a086805780106fd16f89cf21aed88e706e23edd3ad90fd642d494d3c0d3e1d45ed6a7d791d888d854d735d51fd26bceaacaeac684c3edc009bffbbde5bd5cbe3ebf64c054c10dc28fc29ec286c278c25dc295c233c3efc3dfc4c1c520c621c6bac5e7c44bc430c4b6c463c622c9a0cceed089d5dad9d9dd04e1f7e204e41ce458e375e2a2e10fe159e179e25be44ce7e8eacceef5f2dcf62ffa2bfda0ff88014603a50480051e0652060f06be056405190553052706a907150a260d8010ec13de16ed181c1a421a5819bf17a91549131b11690f4b0eeb0d3e0e040f1a10551173125e13011438141014a013dc12e011c210550f980dad0b7e0935073005730320026c01240125016a0190015801b90066ff64fd07fb59f8a4f552f347f18def4bee30ed33ec79ebaeeabee9c9e87ee7efe568e4c4e224e1bddf3edeb1dc47dbc6d959d839d714d6f8d407d4f5d2f8d14dd1abd039d011d0dbcfc8cf0bd053d0b5d021d10fd183d085cfe5cd11cc55caa6c887c73ec7a7c717c97acb2fce04d184d305d595d533d5c2d3bdd16acfefccfacaddc9bbc9fbca60cd73d024d4e9d73edb35de74e09ae1d3e117e181dfaeddf3dbb4da67dae8da3adc81de3fe136e46fe75aeac9ec0def33f1a6f3eff6fbfab9ffc6042209430ca90d930c32091304aefd7cf71bf399f128f425fbb605db12db20752d3737c63c143d9a383f304a25351a1c115c0b5c0a340ee0157b20502c7337e2406c47464a034a0f471b42c93ce937e3338631bd3037313a3360364c3a203f2944e4486b4d0951515387542b541052da4eb04a21464042573fbf3de53d3a3f764185447247cb49754bb04b7e4a734891456c42b33f343d133b6939a937e4352934fe31a72f642df32ada287d277526db258225a3242e231821171ea71a0e173113a70fa80c000a1808e906e105ff04ff0360025400e3fdf1faf4f708f523f2c5effeed9beccbeb42eb71ea44e983e704e51de20bdf09dc8fd9d1d7f4d62fd761d841da8adcb3de3fe0ebe083e000df8cdc6bd9fed5a7d2f3cf6cce4aceabcf82d24bd68adae5ded7e21de6a0e820eabbeaadeaf8e90de94fe8a2e748e788e73de8bbe95fecf9ef95f40dfaacff31054e0a540e3a11f612261330129710920eef0c500cc60cb00e12126d16ae1b6a21cf26992b5e2f8e316a3236321731be2f9b2ecb2db52d612ea62fa6311c34ac3649398b3b1d3d173e503ec03db93c423b8839f0379236ac357235a2351e36b736e936a636fd35b134fe321831da2e8e2c6c2a542889260b2583231622b220131f891d121c5d1aa418d1169d1459120210540d900a96073304de00b8fdc9fa8bf8eff6acf5edf464f4b0f3e1f299f186efdcec8fe9c4e51be2beded3dbb4d933d82bd7bad693d686d697d670d6f4d53fd531d4f3d2bcd177d04acf51ce65cdadcc3ccce3cbb8cbb3cb99cb89cb88cb84cbbccb2fccbbcc8fcd87ce7bcfaad0f6d131d393d4e7d5fdd61ad827d914da32db5fdc84ddecde73e009e2f7e3fae5dde7c9e974ebc1ec05ee1fef0af016f118f201f321f453f585f6f1f762f9b7fa26fc8ffdeafe76001902c103990576073609ed0a630c650d0d0e480e100eaf0d4d0df70cf00c4f0df80df10e201040113112dc120c13ce123d12521139102a0f1e0e330d960c1a0cb90b850b340baf0a120a2609f007b6065e05fa03cd02a30170005bff1ffeaefc36fb6ff95df743f5eff28af07bee9aec00ebfae934e99de85ae8f8e74fe76de6e5e4bfe24ee07adda7da58d86dd625d5bbd4bdd41cd5cfd532d622d6a6d550d456d217d077cde7cad5c820c72cc637c6ebc666c88ecab3ccbece78d03fd132d169d0a0ce57ccf0c96fc773c553c4eac391c443c67dc851cb77ce4ed1dbd3dad5dad625d7c7d6b1d58bd497d3d3d2ced28cd3bfd499d6e2d833dba7dd01e002e2e3e36de579e653e7c0e78fe71be750e62ce531e483e34ae3ece35de5a2e7d7ea8bee78f27cf6e7f964fc02fe86fe2efe94fdfffcfcfc00feedffc30232065309ab0bc70c130ce409e506b00384016301a903bf084e1030197822c52a8a302f334d32e02d1e27441f8417ab11c40e210f2a13421a2023d72ce935ef3c82412043c1416c3ec1396c34b42f0e2ca129fd28e929092c792fab333038173db5419445c948b14aed4ad14931474043dd3e623a6d36da33b2321e335435a0388f3ce340a4445147d948b84809475244a7409b3cd1384e3572327f30032f012e6c2da62cbe2bd42a932942282527f225d124c9236d22cd20d31e251c0d19ae15ea11510e300b660857061c055804180431042b04fb0367032102610033fe92fbf5f889f639f441f28ef0cfee01ed02ebade83de6e6e3d9e182e023e0bfe055e2a7e438e787e917eb7deb88ea41e8e7e4e4e0cddc35d996d66fd5fad50fd87cdbd0df4ee47de8f3eb3eee69ef9befe6eed5ede3ec2dec1dece1ec27eee9ef12f249f4a7f63af9d6fbc6fe16027e053609240db210dc137616fd179c188b18d117fc1670164b161017d7185f1bc81eb8228326082aee2cce2eeb2f683056303430263022306030b630e330f830bc301a30542f722eab2d6c2da82d642eb52f2e319332cd337c3490341a34ed324431592f1f2df42a0729212777250f249e225b215420441f631ea71dc61cfc1b3a1b2e1a07199917861515134510f90cb40985064b037200f5fdaafbf3f9bdf8c0f730f7caf638f6a0f5c0f44df374f1fceecdeb58e8b7e41ce110de9bdbb7d998d802d8c7d7f6d741d87cd8b4d8b1d874d831d8ced75bd7f0d657d693d5b3d49fd38ad29dd1d3d065d06ad0d3d0ced154d332d560d796d97ddb13dd29dea7ded6deb3de42dee0dd93dd66ddb8dd7fdea9df64e17de3cce57ae84ceb14eee5f067f361f5fcf612f8a4f811f953f96ef9b8f92afac9fadffb58fd14ff2f017403b4050c084f0a580c3f0edb0f0311e5117e12b912c812aa1238129311d010e50f0c0f6b0ef30dc30de50d2b0e9e0e3d0fba0f08101e10aa0fb30e610d890b4b09f2066204c80184ff85fde7fbe2fa27fa9bf94df9dcf83ef8a0f7abf662f504f43cf219f0ebed6aeba4e8efe515e349e0fddd10dcb3da2dda1bda72da46db0bdca4dc13ddbedc92dbbad9e3d65fd3b6cfe5cb65c8b9c5bac3abc2bac26cc3b9c47cc60bc85dc967cab6ca85ca01cadcc86fc7efc52ec49cc27ac19fc072c006c103c2a3c3c0c5ddc711ca1ecc8acd8bce11cfecce9bce3aceb3cd85cdb7cd1fce20cf95d02dd218d404d69ed732d99edad0db3addbfde42e011e2ebe3a6e57ae70ce932ea2debc0ebf4eb47eca0ec10edeaedf5ee2ff0d8f1b9f3eaf598f856fb17fee300330302057e065c07d8075c08f208120a1c0ce00e70127d16301a3b1d301f6c1f391eee1bc518d015f613a913b9153f1a91203128f02f5f36d43a823cf53af0361d315a2a622440207d1ed11fdc23a92997306737fd3c1c41324319439441da3e523b0b383535e532a231223132313132d23300360b39673cb63f03439045f6465d474b46bf4356402b3cd5375134cf31b1305b313833f1354739423c763ec43f963f113eb63b85380f35f1310f2fa52cd42a1f298a27162655248722e720371fd61d021d581cf21bbb1b201b151a7418de159c12d90e950a7306d202b0ff89fd74fc14fc69fc21fda1fdc0fd2dfd9cfb4ef96bf618f3e8ef19edb1eae9e8a1e786e686e566e4f1e246e178dfa6dd25dc28dbccda2bdb28dc8cdd0fdf51e004e1f4e007e053de12dca1d970d7d3d528d5a9d52ed791d996dcb2df8fe209e5dce622e816e9c0e96dea54eb48ec61eda1ee9fef63f00bf168f1d2f1baf231f4a6f655fae9fe4904160a6f0ff0133217951843188d16a5137210cd0d230c2c0c2f0ec811c8169b1c58229727db2b9c2e01302730222f992df42b632a5b29ee28f1287d29642a792bdb2c5a2ed72f7031e53214341735b135ca357a3599343f33af31f02f532e212d382cbb2baf2bad2bab2b942bfe2af929912895265f242922e21fec1d5b1ce91ac319c91891173d16ad148a121d10760d720a8907df0459025700d1fe83fd9afcd8fbd9fabbf940f820f6aaf3dbf0a5ed75ea61e765e4d7e1b4dfe9ddabdccfdb2cdbe0daadda6bda39daead965d9ccd8fed7f3d6c6d55fd4d6d257d1e4cfbfce23ce10ceb2ce12d0ecd122d46ed664d8e4d9c1dad6da65da92d97bd899d717d7fbd69bd7e6d8a5daeedc82df0de2a3e408e7ffe8baea17ecf9ecbeed67eeedeeb6efb7f0caf133f3d2f474f64ff839faf0fb9afd06fffbffbb0042017b01c5013302ac028203b004f8057207f108100adb0a3c0bfe0a650a99098a088d07ca0614069e0571053c051305fe04af044104d60331037102b401b5008bff4cfeb3fcdefa01f9e4f6c3f4f3f24ff102f04eefddee9bee87ee28ee61ed40ec77ea34e8d6e551e308e16fdf5adedbddffdd3dde62de67dee7ddfadcd9db60dad7d887d73dd629d568d498d3c8d20dd223d150d0d1cf7ecf8ccf05d084d016d1a3d1c6d1a3d13cd156d051cf67ce8fcd3fcd91cd3cce5ccfb9d0dbd1dcd294d3c0d3bdd39bd355d379d31bd415d5aad691d854da0cdc7bdd66de28dfbbdf10e091e02ae1c1e1ade2bbe3bce4f6e538e761e8cfe95febefecb8ee72f0e2f134f333f4def494f542f607f73ff8baf964fb64fd53fff0004302050336031e03cc029202c60255036b041406e907d309be0b480d770e780f51106111ec12eb147417341a861c201e881e481db11a22171613ae0fc70def0dc9102516471d73254b2d69331d37a237c234532f1b28302047195614fb11dd1293164b1c6b23a92aea30bd356438b13843374c344e30522c8e283b25f32297212021eb21aa233726b0296d2d123193342a377038883809370a344430002cde27b724ad22092206231025e0273f2b432e8330ea31f231b430a72ed82bc128e62543232621bb1fa61ef41d901df51c321c531b0f1ab7188c1765167e15e7144414a013d9129711fd0f020e7b0bca0815065103f7002effcafdfefcadfc74fc53fc11fc67fb78fa34f98df7dff53cf499f23cf110f0d9eea6ed55ecc2ea20e983e706e6fce484e4a7e47ee5dbe672e805ea3debcdeb99eb91eac6e86ee6d7e35ce161df46de49de70dfa3e1abe419e894ebceee69f143f353f48ff439f494f3b8f2f5f17cf12cf130f1aef186f2ecf308f6b4f804fce3ffeb03ff07d20bd70efa101b12f111d110160fee0cfe0ad2099509b10a360dc7103d15211ac41ee62228262128fe28d528b42722266c24b2225e218e203c209a209221fd22e124f226f228e12a712c7c2d212e372eb92de22cb02b422ad4285727ec25b0247b237422c2213421ed2004212f216b21aa21952127215a20f41e2d1d221bbb1852160e14ce11dd0f4f0edf0cb40bbd0aae09aa08a807730643051604c00280014e00f3fe97fd1bfc3bfa1ff8ccf537f3b9f078ee7bec09eb21eaa4e9a8e9fde95ceabceae7eaaaea15ea1fe9c7e738e687e4d5e25ce131e06bdf21df3adfacdf69e047e138e222e3e2e37ce4ede42ee562e587e590e59ce5a3e5a1e5cae51ce683e621e7dbe791e869e95aea54eb7eecbeedf5ee40f078f17bf271f339f4b5f427f590f5eff590f676f781f8d4f94afba7fc04fe41ff2900e4006601850172013401b3002900abff25ffd4fecafee0fe48ff0600cf00ac01890203031503c502dc018300e9fef7fcf2fa17f94bf7d1f5d9f41ff4b5f3a9f39af389f385f338f3adf203f2f1f095ef20ee53ec59ea70e86ee692e422e3ece115e1b3e068e041e058e055e050e065e03ee0ebdf8bdfd8def5ddf4dc8adbe3d926d834d683d473d3f0d247d383d433d63dd85cdafadb09dd5adda6dc50dba0d9abd711d61cd5b4d424d555d6e9d7ead90edce2dd7adfa1e019e142e12fe1d4e0a9e0b5e0d4e056e125e211e366e403e6abe78de965ebdbec15eed5eeeeeebeee43ee92ed3ced5eedfced70ef83f1d4f350f684f80efafcfa1efb82fa9ef997f8adf76cf7d5f7d3f87bfa78fc6efe4200ab018602ef02db0277021d02cf01a601c101e101dc01b6015e01fb00cf00fe00c7013f0338059207ff09f30b1e0d440d440c7a0a66089306b4051e06c907990af00dfa102513cc139512e00f340c5d0895059a04c1053c09680e3c14d619021ecd1f0a1fb21b4b162a10620af8050904c404ce07c70ca31242180d1d452098216d21f71fa91d681b7319e4171c17da16d4163a17e317c918461a381c851e52212a24b226ea285a2ab92a422ae528d726c424f422c621b1218a222a247c26e9280d2bcb2caf2d9a2dcf2c4a2b5d298a27df259924f023a323ad230e2463249924ac244f249f23cb22b12189207a1f4b1e1e1d0f1ce71acb19c5188d173f16e2144613b0114410d60e980d990c9d0bc80a1a0a4d096a085607c805f203f001b0ff87fd98fbbff926f8def6bdf5def43af496f3f6f253f28cf1d0f045f0d7ef9cef94ef80ef48efdcee0deed5ec4aeb79e9a6e741e692e5e4e56ce7f6e918ed6ef06cf396f5cbf6f8f62ef6d3f444f3daf126f16bf19af2b8f46bf71cfa92fc97fef1ffdf0094012102eb021e04ab05bd07310a900cb90e6f105e11be11c21185117811d8119d120314f41519185f1a801c1b1e401fef1f282038203a202f2051209620ea206921f3215d22b422e022de22dc22d822e122172353239023da23fb23e5239b23f022f521ce20751f261e081dfc1b2a1b991a131ab0196c1904198e180318311748164615f5137912bd108b0e2c0cbf09470728057e0322024401c5005e002900fcff8cfff5fe15febffc33fb72f96af758f530f3d8f09cee90eccaeaa4e921e924e9b0e983ea5aeb25ec9cec89ece2eb84ea85e842e603e427e203e196e0d1e08ee17ee279e35be4efe43be549e520e50de541e5c1e5a9e6cce7d5e8abe920ea0eeaaae903e92ae87be712e705e7a5e7e1e885ea9bece1ee05f110f3def445f676f75bf8e0f842f977f971f974f970f943f92ff932f941f9b1f996fad3fb8bfd8bff6d0116033a0482041104f7023f0166ffc5fd7cfceefb34fc05fd4ffec7ffe200760163016900c6fec8fc8bfa7ff8fff6faf595f5caf529f693f6eaf6c3f622f627f5acf3ebf134f078eeefeccbebd4ea1feac1e970e938e92fe9fae89ce829e857e73de60be594e307e29ce031dffedd34dd95dc3adc26dcfddbd1dbbbdb83db5edb72db81dba7dbe5dbe6dbc1db79dbd6da16da61d9a1d831d839d889d84fd973da89db97dc7cddf3dd41de81dea3def5de72dfd4df47e0b3e0e4e028e182e1cbe153e222e31fe49be587e78ee9a9eb77ed91ee27ef43eff5eeb2ee8bee68ee90eefaee8aef79f09af19bf288f349f4e3f4c9f525f7e5f802fb06fd74fe3fff4aff99fe8efd4ffcf8faedf96cf9a4f9c6fa9efcc5fedd0072025803bb03b1035703d8022c025c01a1002e003800d100ce0110036e04b905fa062208eb082c09c0089e072206b904bb0384030d04190596063b08a909c30a2f0b940a2609320732050204160477052f08c00b890f3d133b16d717e9172c16b912860e720a3d07cf0545064308a60be40f5b14c9187d1cd01ecb1f681f041ea61cc41b701bea1bd21cc41df21e42208421d022c7233924a4244025522645289a2a942ced2d3c2e882d762c422b0d2a26296f281b28b528312a582cd92ebb3066310331ba2f162ec02ca32ba52ad329fe286c287528c6281729172933289926e52450232d228c21d420d01f9d1e391d051c2f1b451a181993178d158a130312c810c20fb30e210d400b87091e084207ca061506fd049603eb017a007dff88fe65fdeefbf6f9dcf710f697f47af3a6f2eaf189f1e8f11bf316f571f757f93bfaf2f968f8e1f5c3f232ef79eb35e807e693e55ae729eb40f0b4f584fa00fe02008400a1ffb3fd03fbf7f763f5e7f3c0f30af55ef705faa7fc1fff6501b8031e065808540ae70bf30cbe0d5c0e910e5f0eb80d970c7f0b010b710b100db60ff7128d16201a531d0120c92141226e217f1fe31c621a8d18ab17d917e718a31af31c951f4522b0245226f226a226892509247622c820001f1f1d2e1b8c1988182c188a185e193b1a1a1bdf1b421c451cb21b371a0b187a15d2129e10ec0e750d290cbb0a00095807d5054f04eb028301f3ff9bfea3fd02fdbdfc5efc6ffbfdf9fef79df55df33af112ef11ed2ceb78e952e8aee74ce701e75fe64ce516e4e4e2f5e182e146e113e1ece09ee02de0a9dfc7de71ddb4db99d992d712d635d522d5bfd5acd6e8d766d9ecda7ddcdcdd93de98dee8dd96dc2edb00da1cd9d0d809d98ed999da17dcc8ddcbdfe7e1c2e37ce5fae60be8ece87be985e94de9d2e80fe87de736e731e7cee709e9b3eafceca5ef36f29ef484f693f70df80bf891f70bf786f6e1f563f510f5d3f4fff48ff540f62af729f8f3f8c2f9aafa8ffba6fcd8fdcffe80ffbfff43ff33fea3fc8afa4df846f69ef4c8f3f7f3edf47ff64df8c6f9c6fa46fb2afba6facef976f8c7f6f6f421f3b2f1e8f098f0aef0fbf02cf148f15ff13ff1dcf012f0aaeed6ece9ea1ee9d2e71be7bde6bde620e7d3e7fee88eea0dec26ed8eed0eede8eb64eaa2e8e0e62ae57ee340e2bbe100e22ee3fde4e0e6a1e81cea3ceb38ec0eed89edaeed70edd3ec38ecc4eb5deb0eebb3ea31eae4e911ead1ea44ec23eef9efaaf119f33ff45df568f626f798f7a6f752f7fff6dcf6e6f638f7aaf70bf876f8ecf852f9aaf9c1f977f905f9a6f8a2f851f99dfa32fcdafd4eff6000250197019101ff00cdff24fe68fcf0fa01fab2f9c3f903fa6bfa04fbf6fb5bfd0fffe0009002f3031605f3055c062c0623051a036d00a3fd4cfb0cfa22fa71fbdbfdf70043046e07e5091f0b190be809ea070806e204be04e2050808ac0a990d58106f12cc131f144313c011f20f430e730da30d9c0e7310d21262155118681b561e25216c23d024842568256e24072337210f1f321dda1b451b011cfa1deb20d3241e29412d0e31de333135153561335530d52c60297e26d8245524cc2437260728db299b2bce2c542d792d1e2d6f2cbc2bc12a73290e287a26ff2405245f230123dd228222002299212021a62025201a1f7f1d941b62195d17d7158b147c13a912cd111f11c3105110a40f920ec50c8a0a5108330678041b03b801630046ff59fee5fde9fde1fd92fddafc8cfbfbf979f803f7b1f583f455f362f2e4f1d3f136f2d6f23af32cf3a5f297f13af0d4ee82ed7dec07ec3fec37edddeecff099f2ddf34af4d5f3c2f255f1d1ef91eed0edb2ed70ee23f0a3f2b4f5f1f8d8fb20feaaff7300c000c900a10078006b006d00a4002801d701aa02990382048105c4065808510a930cc70eab100812b412d712b41281128b120313e7132a15a016ff17081986195d19a41894177a16aa155815991561168c17fb18801ae71bfc1c731dfc1c8f1b441963167813e410c80e300de90bc50ae70972099109760ae40b660db10e550f080fe70dec0b14099f05aa0170fd7af912f66df3d4f123f127f1d4f1d4f2c6f37df495f4e4f3a2f2fbf045efe7edd0ecd8ebedeac5e959e8f2e6a4e590e4d4e335e393e2e5e106e11be061dfdedec4de37df0fe049e1d5e262e4dae517e7c9e7e5e75be70ce642e443e242e0b5ded5dd92dd0fde30dfb3e0a6e2e6e423e75fe960ebdeecfbeda6eebfee82eee3edc7ec8feb76eaace9bee9d7eacbec98efd1f2eaf5b2f8ccfae9fb35fcb2fb6dfaeaf869f702f61bf5bef4c4f457f567f6bdf768f937fbd4fc3bfe48ffcfff09000200a1ff1aff73fe91fdb7fc10fc99fb87fbe3fb6cfc17fdc1fd2ffe79feb8fee4fe28ff84ffa7ff6fffb5fe3cfd31fbecf8a4f6b8f46cf3b0f283f2dbf283f37df4c1f509f738f829f984f942f981f83ff7b5f529f49df220f1bbef3aee95ecd5ea02e96de77de662e659e75fe902ecdfee8bf17ff383f487f464f335f12fee89eac3e665e3c8e04bdf04dfb3df3de175e30fe6fae80eece4ee3bf1cff25df303f3e7f132f03bee2eec14ea41e8f4e650e6b2e632e894ea9deddcf0c5f30ef672f7cdf749f700f61cf411f22bf0a9eef9ed48ee8fefd9f1f0f470f807fc3aff8b01ba0291021d01c2fedefbe0f84ff66ff46bf37ef3a9f4d6f6e8f981fd2a017204df06320869089407fe05fd03bd0178ff65fd9cfb5dfaf5f992fa67fc5fff0f030007880a040d4a0e620e800d2f0cd00a84097b08b0070d07c606e9066f076c089a099a0a630bd40bec0b230cb00ca20d3c0f4e1171137f15041791173917fa1516144f120a1184100e114f12cd137e1514176818cb19291b591c861d7d1e241fcc1f5620ab20fc200621a4202b20931fea1e961e7e1e911e141fdb1fd1202322772388246225a8254225862464230422dc20e81f481f521fdc1fd6205c220d24b72552276628c6287b2838271b2586227b1f491c6919de16ee14fe130014041503176c19de1b071e591fc11f571fe61d961ba91817154411b80da10a550805076c067a06250722087209090b790c940d3c0e310e900d8a0c000bf0084f06ed0208ff22fbabf741f54cf4aff438f692f82afba9fddeff7c016e02c1025902370171fffdfc00fadff60cf41ef2a1f1aef208f529f846fbbbfd49ffdcff97ffd6fed0fda9fcb0fb1ffb1bfbcffb24fdc7fe7000cc019e02f102d7026a02f601b701dd01a6021004d00596070109cd091e0a3e0a740a000bd80bb90c7d0d0b0e660eba0e130f4e0f470fdb0e050efe0c130c870b820bfe0be30c0e0e560f9710a81155127712fd11f310860fee0d5f0c110b170a790947096309ac09130a690a880a730a0a0a370905086406650451025700affe91fddcfc61fc02fc80fbd8fa48fad9f997f988f952f9b1f89df702f616f43ef293f033ef32ee57ed98ec11ecadeb81ebabebfdeb67ecdbec0aedd7ec34ecfcea6de9e9e7a8e6f7e5dde5ede5d9e574e5ade4f4e3c4e33ee461e5c9e6d5e755e850e8f4e7bde7d8e707e82ee81ae8ade756e774e723e880e936ebb5ecc3ed2eeee9ed56edb1ec20ec07ec82ec7eed15effff0ccf263f49cf568f622f7dff771f8cbf89bf8aaf758f60ef539f462f489f54bf769f97efb30fd91fe8ffffaffe9ff61ff79feacfd47fd4bfdbffd4cfe72fe26fe76fd77fc96fb10fbd4faf8fa77fb1dfcf0fcd6fd7dfed2febffe1dfe2bfd21fcf9fae6f905f92af871f7eff66ff6f1f572f5b6f4ddf316f358f2d1f194f15bf11ff1e9f099f066f08bf0ebf086f137f27df221f210f125efb9ec49ea1ae89fe61ee66de67fe72ce9fdeab6ec1eeec9eea6eecfed50ec93ea01e9bae7fee6d0e6eae640e7b3e7fde73ce896e80ee9eae942ebc8ec3bee37ef58efc1eec0eda9ecf5ebb0eb86eb48ebcaea0cea8fe9bde9c0eab2ec3cefd2f122f4c8f571f626f6edf4f2f2c6f0e5eeb4ed91ed5ceebcef76f131f3b8f426f665f763f838f9d4f94afadbfa7ffb16fc83fc67fc90fb27fa58f879f6fcf40cf4daf398f441f6d3f826fca3ffb702e504bb054b05110487024601b900e300b201eb0222042105ba05bb054d05ad04fe039803a4031204ff046d063f08860a050d3b0fda108b112a112b10ff0ef60d6a0d3e0d1f0d110d100d2d0dc70dd90e2a10b41130136f14aa15ca169f174a189f1886185c1833180a18151831184e18c21883196f1a7d1b101cb41ba71a2d19e317b817d218de1a771dc41f3f2114224e222b221222c8211e214020121fbb1db11cec1b661b481b501b741bf01b961c641d871eb31fcd20ee21b222dd2270221e21fd1e901c1c1a1e181117cf162f170118ab18f418e518471842172c16f814d41301135212c2116011e91068100610a90f730f800f810f5b0f030f270ed60c500b9c090408d706fd0578053205c90429046a038802d701b4010d02d102d2039404de04b20403040703f701ca009dff99febbfd36fd33fd7dfdddfd28fe16feb4fd60fd5afddefd03ff7500d801f1028703a303760308036a02bd01040163001c003700ab006b013a02fa02be038904620551062307a507d407b50773075a0789070708ce08b0098c0a520be00b1e0cfe0b680b6e0a470930087a076307ef070309670ac80be70c970dbd0d6e0dcf0c130c870b490b4e0b750b630bbe0a7509a1079b05f903220340034a04ce0543075408b6086308a307a20689058d049b03a102b401b40097ff7dfe44fde4fb92fa57f95df8f4f712f894f850f9cdf9b7f904f99ef7bff5d3f300f279f075efd5ee93eebdee1bef93ef18f056f02cf0a2ef98ee3deddbeb85ea67e99be8f7e777e720e7dce6d5e62be7bde78ae870e915ea68ea5beacde9ece8dde7a3e680e598e4e5e393e3a5e3f6e3a7e4b7e50ae7bee8a9ea74ecfeedfaee27efbbeedfedbcecbeeb0eeba9eac5ea61eb65eceaedb2ef4ff196f238f312f38ff205f2b8f1fff1b9f28bf366f424f5c0f597f6b2f7d8f8f2f9b0facdfa90fa48fa33faacfaa8fbcdfcf1fdc6fe13ff01ff9cfedbfdf6fc02fc02fb4afa11fa63fa6ffb24fd2cff58014e039004f7047004f602f100d9fefbfcaafbfbfaacfa9dfab2facafa12fbadfb77fc60fd3dfebafed8feb6fe51fecdfd31fd3ffcf0fa63f9b4f750f6a4f5bdf594f6e5f721f9eef917fa72f93bf8b9f60af575f330f23bf1c7f002f1d3f12ef3d1f42ff6edf6ccf6abf5e4f3f0f124f0e8ee61ee5deebbee41ef9aefb5ef86ef09ef8fee59ee7dee1def0cf0e1f065f177f114f191f02ff0faeffeef05f0d0ef68efd5ee27ee9aed40ed25ed88ed84ee2af085f23ff5d9f7f9f943fb9efb45fb6bfa3bf9e4f768f6eaf4b1f3e6f2c1f25af379f4f1f5abf781f97bfba0fdbaff9f011e03fe0353044304d5033b038c02c4012001d600fa00ba01000382043406f4079709440bdf0c200efa0e460fe80e340e600d8a0c080ce40b100cd30c290ef20f36128c146f16c1173e18db171b1740167b1542158d152e1641178018a219b81a851bec1b3c1c701c971c111dbc1d6e1e4d1f12208b20e8200121ca2091204120ea1fec1f3020ae2097219622642307242c24bf2313233222612117214721ef211a234224102575251725fc238a22d820371f161e601d0e1d211d301d1f1d0d1ddd1cc41c091d721ded1d641e5f1ec11da51ce81abc187d1635143012c010d00f6d0f8c0fc00fe70f0310da0f900f4b0fd10e160e1c0db30b160aa1087607de06eb06340775076e07b9066505b903d8011700c7fee9fd8ffdbbfd35fee9febcff6800da000c01cf002a003afff7fd89fc35fb1efa6cf93ef973f9e2f96efaf2fa71fb04fca4fc43fdc3fdf0fdb4fd29fd74fcc9fb58fb2bfb2ffb58fb97fbe6fb4efccdfc51fdc8fd1ffe45fe45fe38fe2bfe3afe7dfeeefe7cff15008f00c300ac005700e3ff83ff57ff62ff9bffe8ff34008700e00037018701ae0183010e016c00b7ff2affe7feddfe00ff40ff74ff95ff9dff6cff06ff7efedbfd51fd15fd18fd47fd7ffd72fd0dfd6afc91fbb1faf3f93df995f80df889f71df7e7f6bcf692f678f64df621f612f6f2f5a4f517f512f4b4f252f113f03feffceef8eef5eec8ee24ee2bed27ec26eb5aeadde96fe90fe9d8e8b8e8dbe85fe900ea9cea0aebf3ea67ea8de957e803e7c2e583e491e32be340e3ece30be516e6e1e645e70ae772e6aee5a8e498e3a2e2c5e16ae1c8e1b2e21ce49ee59fe619e71de7aee642e6fce5a1e54fe50be5c9e4f4e4ace5a6e6cae7b1e8e5e8a2e826e89ae77fe7ebe79fe8ace9e0eae9ebd9ec7aed79ed11ed67ec9feb4beb95eb3eec35ed1bee8aeeaeee9dee5dee42ee51ee6beed9eeb5eff6f0ccf2f4f4ecf679f83df9f3f8e3f747f652f48df244f18af09bf05df17ef2e0f341f56bf685f795f892f9a0faa5fb6afcf4fc28fddbfc26fc0efba3f946f846f7d5f633f740f898f9f1faf5fb67fc6cfc39fc01fc0dfc73fc18fde7fda7fe0fff0eff95fea1fd68fc17fbc5f9a5f8d9f771f79cf76ef8ccf992fb7afd20ff4f00ee00f2006f0077ff08fe41fc4afa5af8c9f6d1f575f5b0f565f663f7a1f81ffabefb50fd94fe39ff15ff23fe7efc6cfa3df835f6adf4edf314f415f5adf66af8e0f9ccfa2ffb44fb44fb51fb60fb42fbd9fa38fa9df95bf99ff952fa2efbcbfbddfb6efbbafa13fae0f943fa22fb66fcdcfd4cffb100f501e902800395030b031402d40081ff8afe24fe62fe7dff55019403140678085d0ad20bdd0c870d240eab0ee70ef20eab0e120ea80da20dfc0ddb0ee40fa61038119c11f711d6123e14f5150218fd19971b151d6b1e791f752017210e219020961f411e291d7a1c551c271dc71ef320a3233426152845298129e62822286827d826cb26fb263827b8273d28ad282f2965293129ec288d284e28a5284c29072ad22a372b1b2bd12a302a4e2972285b271b26142521245c230623c1227b2262222d22ed21d92197211b218420801f2d1ee11c761b241a42199c1849186f189e18aa188c18d8179c1625156a13b31157102c0f4f0ee80daa0d980dc00db90d6d0de70cdc0b5f0ab208c306d1043803000266019b015a027403bb04b60548068d066906f9055e056d042b03d00171005affd3febefef5fe45ff56ff19ffbdfe57fe16fe20fe57fea4fe06ff6dffe2ff74001401b1013b029002ab0293024202cf016001100104015b010402ce027903cc03ae0332039702280210025a02fb02c9039c04640509066c066906d505a70408034501d4ff27ff66ff89005402540423068a0759088e0847088c0779062c05a303fd016600ebfebbfd0dfdd7fc15fdc4fda7fe94ff750009012001990042ff37fdd1fa67f87ff685f564f5f3f5f2f6e1f785f8e0f8d2f86ef8d2f7edf6def5cff4b2f3a1f2a4f186f05bef57ee80ed1aed4cedcfed73ee04ef20efc8ee14eeeeec84eb04ea6be81be771e66ce61ee74ce847e9b8e97ee987e85be77ce60ae634e6d4e66ce7f0e759e879e88ae89ce85de8dce728e729e642e5bfe491e4dce47ce5fbe556e67ee649e614e616e62ee68fe62de7a5e708e852e84ce83ce843e83ee86ae8cce824e995e914ea5feaa5eaeeea0beb2deb4ceb1debbeea34ea66e9bfe87de899e852e98eeaf2eb82ed10ef43f01ff174f1f2f0d0ef49ee9fec75eb20eb90ebc2ec50eebbeff7f0ecf18bf225f3c6f341f4aff4eff4c8f465f4d3f316f37cf218f2dcf1e9f11df24ff2a8f22cf3d5f3d5f411f649f77bf883f944faeefa7cfbc1fbb9fb35fb18faaff846f72af6c8f530f637f7c7f89bfa63fc0efe68ff30005e00dfffaefe13fd45fb75f9fbf702f79ef602f72cf8e5f9fefb22fee7ff2701d501ed019901ed00e1ff8efe08fd70fb16fa31f9c1f8c0f8fff834f951f96ff9a6f927fa06fb15fc1afdd6fd0cfeb4fdedfcd5fba0fa75f962f87ef7e3f69cf6bbf647f724f82df937fa14fba8fbedfbecfbb4fb53fbcefa1efa3df929f8eaf696f55cf460f3cff2dbf299f302f50ff785f90efc69fe4c007c01f601b801c9005dff9afdb1fb0ffa00f9b2f85cf9d6fabcfccefeb00018022603f00382041d05bd0538069b06ce06b30686065b0634065806d2069707e408b10acb0c340f99118e13111508167716c71619175e17b717ec17c51779171217a2168016aa160d17e3171f19b31ac91c191f452130237624e524c0240924de22ab218120881f311f7e1f6220e2218523e6240426ad26fb264c277c2771272c275326e42445238721e11f9f1e801d6d1c991bf61abd1a491b631cdb1d871fd3208521a821f620741f571d7c1a2217d213c5106c0e3a0d080dc20d510f2611eb126c142115dd14bf13ba11210f6e0caf091107c0048e029a0032ff5ffe56fe3cffb8007f024e049f0545065106b40598044003a901e9ff2cfe76fcfbfa00fa93f9c3f987fa8dfb98fc8efd3bfe96feb2fe75fecefdd0fc84fb20faf9f848f835f8cdf8e9f959fbf5fc80fec3ff9700d5007f00d0ff1effc4fe01ffcbffde00e0018402ac0274020b02a2015b0144016601cf0187027f038b047005f7050606b3052e059a041404a503490312032903a5038904ac05c706a0071b083e0830080d08bc0725073906fb04ad03ac022b023502a5021b034d031f038402a401b300c1fff0fe62fe18fe24fe88fe09ff74ff9cff45ff6ffe3efdb9fb0efa72f8f4f6d5f55af582f54ef692f7caf8a1f9e6f967f94ef8e2f634f57bf3e4f162f01fef3bee8ded22edf8ecd4ecdcec3deddaedcbee03f019f1eef170f261f2e1f10bf1b2ef08ee3fec5dead7e80ce8eee79de8fde988eb12ed6cee2fef6def38ef72ee6eed73ec7aebd2ea93ea7aeaa1ea08eb6bebeeeb91ecffec48ed6eed4bed39ed74ede3eda5ee8bef0cf01ef0bcefd4eedaed1ded88ec41ec32ec04ecd6ebbbeba6ebe4eb84ec4ced4cee5aef18f097f0ccf089f013f08befe4ee5beefdeda9ed97edd2ed44ee12ef0cf0caf02bf1f6f008f0c9ee97edb1ec84ec13ed20ee94ef25f181f2a2f358f469f4eff3e6f25af1baef52ee5fed41ed09ee8cefadf107f428f6d9f7d9f80df9b4f8f4f7f0f6f5f50ff536f491f325f3ecf208f371f30ef4e4f4e4f504f75ef8e1f962fbbffca9fde1fd6cfd69fc13fbd2f9ecf87ef899f827f9fbf9fcfa07fcf9fcc7fd67fed0fe14ff3eff4bff3dff0dffb0fe30fea3fd20fdc1fc94fc96fcc1fc0cfd6afdd2fd3afe94fed8fe13ff59ffbeff54000e01b9011b0206025d013b00e6feaafdcdfc81fcbcfc54fd16feb9fe11ff1affdffe89fe57fe62feb5fe54ff1000bb00440182015d01e7001d0011ff0bfe3dfdd7fc19fdf3fd37ffc0003f02760376043405b105150643060e067e057e041603b10195000c008100ef011c04e006bf09420c600eed0fd7105c116311c710af0f190e2b0c850a820965098d0abe0c940fe81241163b19dd1bd81deb1e3d1fb21e551daf1bfd198418d517f317cf18841aa41cc41edd209022bf23c52496252d26c9261a27ee268526cc25ee246f2439243c24a224132576251f26ef26df271a292c2ac72a012b9a2ab629da28fa2726279726ea2503252c244723802244225b22b2225f23ec2330244b24eb2314230c22a9200c1f931d161cb21aaf19d1181f18cc1786173417eb1653167915b014f3137d139013d11309141314741322125d10210eb50b77095e079f058b041b047504ae0552070109620ae60a710a3c09670751055a038401f3ffd0fe12fee6fd6afe66ffa900f801ef027b03b803ae0385035103e6022f022a01ceff50fef4fce2fb4efb53fbe2fbeffc57fed6ff3b015c0214036c037b034803e102430266015d0055ff84fe20fe3cfebbfe6fff2500c3005301e90192023e03bd03e3039f03fd0230026f01cb004000b1fff6fe13fe1ffd43fcb8fba1fbfcfbc3fcd2fde6fed0ff5d006200eaff0fffe7fda6fc66fb28fa0df932f89ff777f7b0f70df86af89df87ff830f8c8f73df79df6dbf5d5f4b1f39df2a9f109f1c4f0a5f0a7f0b9f0aff0a0f08cf04af0f2ef96ef22efc8ee98ee67ee3fee1feee0edaeed9bed79ed50ed12ed8becf4eb85eb33eb27eb4feb49eb12ebb9ea33ead7e9cfe9dbe9f4e9f7e9a0e92fe9e6e8c1e8fae888e90aea82eaf1ea25eb5debb0ebe3eb12ec3fec29ecfaebbfeb3beb99eaf2e926e984e835e80ae826e882e8d7e851e9ffe9a4ea5aeb09ec52ec57ec33ecd1eb85eb6deb45eb1eebe8ea63ead6e970e920e92de99ee927eadaeaa3eb38ecc2ec44ed84eda7eda3ed35ed8cecc0ebccea18eadbe9f8e98dea6beb22ecaaecefecccec90ec6aec49ec6decdaec5ded1bee0cefebefc2f06bf194f15af1d2f0ffef42efc8ee71ee50ee44ee0ceed1edb7edc5ed46ee4bef9af02ff2dbf346f568f620f730f7b4f6c9f575f411f3d7f1c6f012f0ceefedefa5f009f2e6f31ff662f835fa73fb0dfcf1fb52fb49fac4f8f0f603f531f3f3f199f11cf265f327f5ebf68cf801fa3cfb61fc6efd2cfe83fe5cfe9ffd7efc2efbcdf997f8b1f714f7dcf60bf781f73ef82ef926fa1ffb03fca9fc0bfd1cfdd1fc4dfcb2fb16fba7fa72fa70faa9fa12fb98fb38fcd9fc65fdd7fd20fe3bfe35fe09fec1fd7cfd49fd3bfd5bfd7dfd76fd29fd8afcd3fb65fb7cfb41fc97fd17ff780091015102e7027303d9030a04e7035e03b3023002f6013202ca0279033d041205eb05f60626083e093f0a110b990b0d0c6a0c8d0c910c680c0a0cca0bc40bea0b600cfb0c890d430e370f65100d12fb13d5159117ea18b2192a1a491a031aa5192a199d186b1899181a191e1a561b751c971d801e111f951fe81ffe1f222032201a201a20fa1f9e1f591f161fee1e481ffb1fe5202b227923b62423267e2795286b298229a82831272d25fd224421fb1f281ff81e111f601f1a20f320ce21c5227623cd230024cf2338236b2222216e1fb21de91b591a5d19c2188d18e8189819a31a1e1c8a1d921e021f651ed61ccd1a79183f166f14cc1254112610240f8b0e930ef70e920f33106a103310b30fd50ec90db80c870b650a8c09f108b108ca08e108db08a7081e086707a806cf0502056304ee03d40321049204f60408057a046003ef015000d3fe9cfd9ffcf6fbabfbb7fb2afce5fca3fd40fe9bfea9fe9bfe8cfe76fe59fe0bfe6ffd9ffcb4fbdafa48fa05fa0cfa61fae7fa84fb2bfca6fcd0fca2fc0ffc3bfb5afa82f9c6f82df89af70cf795f635f602f60df63bf689f6f8f675f70ef8c4f86ef9f6f942fa26fab5f913f94ef898f708f781f607f691f5fff46bf4e9f372f32df32bf356f3bef358f4eff478f5d4f5ccf56df5c5f4d4f3dbf206f25af103f10af14af1ccf176f204f369f386f32cf380f2aaf1bcf004f0a6ef8eefd4ef6bf024f107f2f3f29af3edf3ccf313f302f2caf07aef50ee58ed7decf4ebe0eb3dec2fed8aeee4ef17f1f4f15cf291f2b4f2b1f29df264f2e7f166f10af1d5f0e8f020f12cf113f1d7f078f03ff043f062f0b2f025f19af13bf201f3bbf36df4f6f429f52ef513f5ccf482f437f4daf3a7f3c1f32cf40bf53bf665f769f817f94bf935f9eef87af808f8a2f742f721f757f7dff7cdf8faf91cfb18fcc3fcfefceafc9cfc18fc8cfb06fb81fa29fa15fa50fa02fb26fc8dfd0bff52000d0125019f0096ff5afe2cfd28fc74fb1dfb1efb91fb7bfcc0fd3effb100c60153024902af01b60091ff60fe4ffd7ffcfafbcefbf7fb52fcc6fc42fdb6fd2afea6fe13ff57ff56fff4fe44fe78fdc0fc48fc21fc33fc62fca2fce6fc35fd91fdd8fddcfd7efdaefc97fb94faf6f9f4f996fa9dfbb2fc96fd1cfe44fe2ffeeffd8cfd0afd5efc8ffbbafaf9f964f916f911f953f9def9a0fa7ffb5ffc1ffdaafd05fe38fe47fe2afecbfd14fd15fc01fb24fac5f906facffae0fbf5fcddfd8cfe14ff81ffceffeaffb9ff2bff57fe5dfd62fc93fb04fbbbfacdfa39fbf4fbfbfc2ffe69ff9900a4016602d902e3026e02a001a600b9ff31ff30ffa0ff6f005e012d02e2027703dd032e0452042804d2036203ef02c202e2022b03a3031d047404d7044e05d705a20699079408a609b00a890b4f0ce70c2f0d560d4a0df80c950c150c720b010bd60a000bc20bf00c440ebd0f1911351252135c143515ee153b16e9153b154d145b13ec1208139513a014ce15dc16eb17d7189b197b1a501bfd1ba71c131d2c1d331d141dda1ccf1cca1cad1c981c501cd21b771b421b561bf71bdf1cce1db61e351f331fee1e5b1e981deb1c301c6b1bd81a611a251a651aed1a9e1b6e1cfc1c2c1d241dce1c4c1cd61b3a1b641a5e19ee172e167114c8127611b91062106010a510e3100f113a1136110d11cb104110780f870e5a0d130cda0aa3098c08b607080798066d065b065e0667064106e5054a0553041b03c4015d001eff21fe53fdb7fc37fcadfb2bfbbcfa5cfa22fafef9caf981f916f986f8faf77cf70bf7b0f64ef6d4f555f5d6f46bf433f41ef413f409f4dcf38cf337f3e1f298f263f218f2a2f103f130f04fef96ee0feed2ede6ed19ee59ee93ee9bee7aee48ee05eedeedf3ed2fee96ee1cef8cefecef3ff065f06af049f0d4ef23ef50ee60ed94ec11ecbeebb2ebe6eb36ecbeec80ed4aee16efbbeff4efd3ef6befbfee18ee95ed22ede8ece9ec06ed60edeeed79ee09ef86efc3efe8ef03f0fceffeef08f0f7eff5ef09f010f028f036f0fdef96ef05ef47eeaeed5ced3eed7ced04eea3ee73ef5bf01df1bef11df20ef2ccf17af121f104f11af12bf148f15ef156f165f18cf1a0f1b4f1aef16df12bf100f1eaf024f1a7f14af224f317f4f0f4bef567f6bdf6e0f6bff631f656f525f4a0f22bf112f090efffef53f13ff395f5fbf71bfaf8fb72fd55fea3fe32feddfce3fa81f807f605f4cdf27ef239f3cbf4d7f628f96afb50fdd5fedaff3d00150057ff08fe76fce3fa8bf9c7f8a5f8fef8bef9aafa93fb8afc8ffd94fea1ff8d001c014401f200240010ffd7fd92fc7dfbb4fa44fa52fad6fab1fbd1fc09fe28ff1f00d30023011701ad00ebff02ff13fe26fd4ffc80fba8fae4f95af933f99ff999faebfb5dfdaffeb3ff6d00dc00f0009f00ceff73feb9fce3fa3cf90ef879f770f7e0f7a6f89af9abfabefbb1fc76fdfdfd3afe35fee8fd4cfd6cfc5afb3bfa48f9aaf86af87cf8b9f8faf839f97ff9e1f973fa2afbe9fb92fc0cfd4cfd5cfd3efdeefc68fca8fbbdfacef904f985f86cf8b1f845f912faf7fadffbb5fc5ffdd2fd10fe1ffe12fefbfdd6fda1fd54fde9fc71fc09fcbffbaafbc9fb08fc69fceefc99fd7cfe8dffa4009b0142026f022b028b01ab00bcffdbfe14fe8afd51fd76fd1afe34ff990027029b03b9047905d905dd05b0055805ce0429046a039e02f80191017201bb0163025703a1041c069307e508d509380a320ae20975092d090209cf088d081f088b071707de06ea064e07df0782085609580a8c0bfd0c670e7f0f2e104f10f00f5b0fa70ee00d2c0d760cc70b600b4c0b9b0b640c6d0d860ea90fa7106d111112691267122d12b5112511bd1073103f102a100810e20ff10f3510bd108f115f12fb125f1365132313cc125012ba1126117b10d30f5d0f0b0fee0e1d0f710feb0f97104111d31144125d122712ca114011ac102010740fa90ed80dfd0c4b0cf00bd00bea0b310c720cb80c160d6c0dbd0dfa0dee0d9f0d250d7f0cd40b310b6f0a91099e089207ab061706d305eb054d06c3064e07e7077008ef0852096c094609e8084d089907cf06d405b6047b032f0214015200eaffebff3900aa0048010c02e102cb039e0420054305f7043c0443032002db0097ff5efe40fd72fc08fcfefb5bfcfbfcb3fd80fe49fff7ff8c00e100cf00590077ff40fefafccffbe5fa6afa51fa81faebfa5ffbbbfbfdfb15fc05fcebfbc2fb8efb62fb30fbf7facafa9efa72fa55fa31fa02fad6f9a6f97bf970f97cf99ff9dff921fa56fa80fa84fa5cfa12fa9bf907f974f8e9f77cf748f749f782f7fcf79ef855f90efa98fad9facffa73fae4f952f9d2f87cf860f868f88ef8d1f81ff977f9dbf934fa75fa9afa8bfa4bfae9f96ef9f8f8adf899f8c8f839f9c9f95efae5fa48fb89fbb9fbdafbf6fb16fc29fc2bfc1dfcf7fbc2fb94fb75fb76fba6fbf5fb56fcbbfc0cfd48fd7efdb1fdeafd2ffe67fe80fe70fe2dfec9fd63fd0ffddefcdafcf0fc17fd54fdabfd2ffef9fef9ff11011102bb02e9029d02e801f400f6ff09ff42febcfd7efd99fd19feeffefdff20012502e8025d037b034a03df0245028b01ca00040047ffa8fe34fe06fe41feebfefaff4a019702a5035504980483043804be03170343023b011a0017ff5dfe13fe46fed9feabff9f0094017a024203ca03fb03cd03400374029101ab00d5ff16ff68fedffd97fd9ffd02feb1fe80ff4f00070196010402520270025a020e028c01ea00380073ffa3fec9fdeffc41fce5fbeffb61fc15fdd3fd7bfef5fe3fff68ff6fff42ffdefe3bfe62fd7ffcb4fb19fbcafabffae9fa45fbb7fb2afc98fcebfc22fd51fd75fd8dfd96fd6cfdf6fc3bfc3ffb26fa2af966f8f9f7faf75ff81ef92efa5cfb7cfc66fde2fddcfd65fd8bfc7dfb71fa7bf9baf84af826f859f8eef8c4f9ccfaeefbfbfce3fda1fe1eff5dff62ff14ff7efeb6fdc4fcd7fb17fb8dfa52fa75fae3faa1fba5fcbdfdd0fec1ff6900d800230146014f013201ca00250064ffaafe3bfe3afe91fe30fffdffd500d2010003450482057306c206600668050f04b902ab01f2009a009300bb002101c9019e029c039f04720509065e066c0659063106f005a6054d05dc046d041104d003ca0305046d04fc049205010641064a061d06e605bd05ab05be05e305f405e705a9052d058b04ca03f4022b0286011b0117018a016f02ba0337059e06b80750084908be07d806ca05d5040f047303f70282020b02b0018901a8011202a0021e0374039a03a303bd03f80344048504890435049d03e2022f02ac016201470153017e01c20123029502040363039f03b303a6037d033f03fc02c402a902b902eb02210337030b039602f0014401b60059002300fbffd3ffb1ffabffddff4e00e9008501f70122020b02cc01860153013c0139013a012f010d01d30085002b00cfff7bff38ff0eff06ff21ff5effb6ff1600620081005700daff14ff1ffe24fd51fcc8fb98fbc6fb42fcf4fcc7fda2fe6cff11007a0096006300edff4dffabfe27fed3fdb6fdbffdd3fde0fdd6fdaefd71fd25fdd3fc8dfc5dfc4ffc71fcbdfc23fd91fde4fd06fef5fdb9fd69fd26fdfefcf1fcfbfc0dfd21fd43fd7dfdd4fd49fec1fe1eff50ff4aff14ffc3fe5ffeecfd72fdf3fc7dfc2ffc18fc3cfc95fc00fd5ffda4fdbffdb4fd8efd51fd0cfdd7fcc7fceefc53fddcfd5efeaffeaafe49fea7fde4fc26fc92fb35fb20fb5ffbf3fbcffcd8fdd6fe8effd9ffa2fffcfe19fe26fd49fc94fb01fb86fa23fadff9cdf9f9f95efae7fa76fbeafb2efc40fc26fcebfba2fb5efb36fb43fb94fb24fcdbfc88fdf5fdfafd88fdaffc9afb7efa8ef9edf8a9f8b6f8fff86cf9e4f960fadcfa4efba8fbd4fbb8fb50fbb2fa02fa71f926f926f966f9cff945fabcfa32fb9bfbf0fb2bfc3cfc25fcf2fba7fb50fbfbfaaefa7ffa86fabefa1afb75fb9afb77fb21fbc0fa94fac1fa2ffbaffb07fc08fcc0fb64fb1efb19fb5afbb6fb12fc63fc9ffcdffc30fd7afdadfdb4fd7bfd1ffdd0fca6fcbffc16fd7ffde8fd46fe8efedafe32ff78ff97ff70ffe3fe09fe0ffd1afc67fb18fb2bfbacfb8dfca2fdc7fec6ff57006f001f008cff0dffdcfe01ff7cff2900d0006301cb01e2019d01e600b0ff36fec7fcacfb38fb7ffb51fc86fddffe28005b016a022b038c0365039b025401c7ff30fee5fc0cfca4fbb0fb12fca3fc5dfd2bfefafed6ffbc009c0177022e039703a4034a039302b401d000f5ff2cff5efe6ffd77fc9bfb10fb19fbc4fbf0fc69fee0ff180101029902e402f502c50248029001af00c2fff9fe6afe17fe04fe1dfe50fe9efe00ff75ff0a00c10090016d022f03a803ba035b03a502d30117018d003200e7ff90ff33fff1fefafe71ff46003f0115029002a3027602430239026902bd0212034703550346032d0317030803f702dd02b4027f0245021102ed01e80113027102ff02a4033a049904a6045704bc03fa022f027b01f4009e008100a7000e01b701950283035804f0042805020599040c0486032803f102df02e802fb021b0351039003d003fa03e8038e03f3022b025f01b800440009000a0034008f002501ec01db02d803ac043205550503055404720377029001e40078005a008e00f9008f0148020a03d1039b044505b805de059005d104bf0372021f01f3fff2fe29fea5fd66fd8efd4bfea0ff8701d2031a060b086809fc09ce09f908830787052e03a10041fe86fcbbfb12fc77fd80ffbf01dd039305de06d6077108ac087d08c6079b063305b70368027301d20084008500b30003017201e1015502e2028803560453054b061a07a407c70799074707dc066706e5052a0530041f03210284018601160204030b04ce0433055c0564057a05ad05bf057a05c704a40360026b01ff003701f801ea02d1039c043f05d2056b06e70628071f07b5060206340552046d039302b901f5006e002b00370092001601b8017b0246030904a904e5049f04e903e302dc012101c100ad00c500d400d200e0000c016b01f6017502c202d102a00250020702bf0170010f018900f2ff77ff2dff27ff61ffaaffe4ff0200fbffe4ffdbffdaffe0ffe7ffd4ffa1ff5cff0dffd0fec3fee6fe38ffaaff1200540060002b00c9ff5fff07ffddfef3fe3bffa4ff19007700a800a4005e00dbff33ff7afed6fd6ffd59fd9dfd2cfed4fe5cff98ff6cffe7fe44fec0fd9afdf1fdb3feacffa3006101d3010b0225023a0250024c02080270018b0084ff9ffe16fe00fe52fee0fe77fffcff6c00d4004601ba01180240022002c1014a01e900bb00cb0001013e016c018a01a201ce011a028302fe027a03e6033a046e0477044a04e6035703c102530230026102cd02400384037e033603d9029d02a7020303a50370044a051a06c0061607f70649061a05ab03570275013a019d0168025e03510433051206f306c10758088d084b08a507c506d705fb043d049403040397025d0260029802ec0247039703e2033b04b0043905c30525063c0600067d05c9040f046903e0027a023202fe01e301ed01210289022503d9038204ef04f20471046b03f5014900a4fe40fd5efc29fcaefce4fd9dff800132036104d50488048f0301020100aafd24fbc8f809f74ef6dbf69af811fba8fdd3ff4101f6012202e801580168000bff63fdb6fb47fa3ff98ef8f5f742f776f6c2f576f5cdf5c0f61ef89bf9f5fa20fc20fddcfd36fe03fe1bfda3fb02fa9ef8c4f77ef782f76df707f756f6a1f537f53df5aef55ef61ff701f834f9cbfaacfc70fe6eff2aff91fdf6fa0ef89ff519f48ef3c1f33ff4b5f403f524f534f563f5d0f5a6f604f8dcf9f4fbe6fd31ff87ffecfe9ffd18fcc7fac8f904f950f875f776f68df5f1f4cbf426f5dcf5c9f6d7f7eff812fa35fb2dfcd6fc1efdfdfc98fc32fceafbd1fbddfbcefb6ffbaefa90f94ef83ef79bf68ef620f725f872f9e6fa4ffc8afd76fedcfea7feebfdd9fcd3fb38fb25fb7cfbf0fb12fca9fbd3fad8f92bf931f9fdf95ffb01fd6cfe4dff82ff03fffffdbdfc75fb65fac4f99af9e8f99afa77fb50fc0afd86fdd0fd0efe56fec4fe67ff2600df006d018f011401e9ff18fef1fbfdf9c2f8a9f8c1f99dfb9efd26ffc8ff90ffdffe12fe74fd1bfdd5fc81fc31fc13fc67fc55fdb5fe28004001a9016201b200f2ff7eff7cffccff4000aa00dc00cd007400b2ff75fec1fcaefa98f8f5f619f637f648f7fef8fcfaf9fcb8fe22002d01d00118021602da0187012f01c300360079ff76fe3bfdeafb95fa54f942f874f70ff73bf709f862f9f3fa42fcedfcc6fcf2fbf4fa60fa91fa97fb1dfd85fe51ff44ff6ffe35fd04fc21fb9efa5efa30fa03fadef9d5f9fbf93bfa62fa42fabbf9dbf8e8f72cf7e6f646f745f8acf940fbb4fcbffd46fe57fe21fee8fdcbfdc1fd97fd09fdfafb9efa50f973f847f8aef850f9d7f90afaf2f9cdf9cef905fa64fac2fa0efb62fbe9fbc2fcedfd2aff1f007d00180011ffc4fd9cfc06fc47fc47fdb9fe35003e0189011b012300f0fed1fde1fc14fc52fb87facaf956f96af938fab9fb9dfd7dfff200b501cc0190016d01cd01dd026f0426068b0741084008bd07e506e005b4042f033701ecfe8ffc81fa1af980f8b3f8a0f92cfb4efde3ff9d0229052e076d08f9081a0915092009430958094109e60837083807e4052c043a02660014ffb3fe6ffffa00cc0252041d052505bb0443040d042d048804fe047505e1054e06ac06d006a1061c065d05a604350428047f040905940512067806be06fb0635074f07400701077b06ad05a804830368028a0112011901930169027d039f049d054f067d060006e704770323027f01e101410341052a074908470832076a058303ea01c4001100baffa7ffe6ff840076019502aa038f0436059c05c1059a050005e1036302cb006fff9bfe54fe70fec8fe43fff2ffff006302d603f1044805ad046703fe01f6009400bb001001420132010a010e015001a801ca017901ca002500faff7f008b01a00249036f034d035703d9039d041505bd045b0339010eff84fde8fc18fda2fd28fe94fe0dffcaffe000260259034804ec046f05fc0590061207630767072507ac06e205a004d6029a005afed2fc91fcbafdf7ff78025504fb045c04d8021201afff20ff84ffae005002f4031205650501052a045b031303710342043705fe058006e8066a071708cb082809d808b807d2056903e20086fe92fc39fb92faa0fa50fb6cfcc2fd3bffcc008a028804a0068b08ef097b0a320a6e099f082a08380881089608230800076205bf0362026401bd003400a3ff24ffddfee6fe4cfffaffd200c901eb024704c70526072f08ba08a70816083b071006980408039e01ce002101b2022505d607f709070b220bc30a7b0a9b0aea0add0af90909085a0595024900c7fe0ffed3fdd4fd0efe90fe82ff040100035005c707230a330cd00dbb0ee80e880ed10d140d950c390cbf0beb0a810987075605410386015400a0ff4dff5cffd1ffc0003c022f046a06aa08900adc0b6b0c220c1e0ba009da071906ac04a7031e032703a9039004de055a07b508ae09ff099709b608bc070c07e0060f073e0711074b060605a10367027f01e6006000c3ff2affd5fe1eff3900000219040a064b07a407380749065305e7044e05950681086b0a8f0b6a0bd6092c073404b2011c0073ff3ffff9fe58fe5afd4bfc98fb74fbdefbc8fc1cfed9ff09028d0420076309fe0ae00b340c210cb60bc60ae208c5059c01f8fcc6f8fdf51af50ef657f825fbc1fdd4ff56018302be03440516070309a30a710b010b31093c06af023cff95fc16fbaafafafa97fb1efc76fcc5fc2ffdc3fd7afe29ffa9ff0400700020011c023003f103e403c302bd0071fea0fcf3fbb8fcb0fe37019c035705220614066d055704e1020b01cefe2cfc5df9baf698f439f3b7f2edf288f343f406f506f6c1f7bbfa20ff8b04090a540e5510a80fbe0c9e0885046d0192ff8afea4fd2dfcc3f995f632f33cf045eea7ed5dee29f0aff28df56ff81ffb94fddffffa01c3030c058805f8047b038401a3ff6afe21fe90fe2bff53ff91fed1fc5bfabcf78cf53af4f9f3cdf458f603f850f9dff997f9e2f859f866f82df954fa2bfb39fb73fa47f997f834f95cfbb1fe4402d4046a05a803dafffcfa4af6d7f240f167f195f2f6f3d7f4f4f4b4f4b1f458f5daf6faf820fbe6fc1dfec6fe1dff41ff1effa0fe9afdd4fb5cf952f6d3f24fef59ec6eea06ea43ebb5edb7f09af3d3f560f79ff801faeafb56fed600ed020f04c3030d022aff67fb53f772f31bf0b3ed71ec41ec04ed51ee70efeaef79ef28eeb5ec14ecedecb0ef30f484f9adfeba02cf048d04ff0184fd11f8eaf242ef04ee44ef1ff248f560f795f733f62af482f221f216f397f4daf529f615f5f8f274f0feed22ec35eb2eeb22ec14eec5f00df4a8f713fbeefde1ff8a00defff5fdfffa9af75ef4a5f1cbefcdee35eeb7ed12ed26ec5ceb33ebf5ebeaede5f042f477f7edf918fb05fbe6f9e9f7a2f58cf3c9f1a2f02ff033f0a5f079f165f238f3a9f339f3aaf119ef12ecade9e0e82cea94ed2ff2a0f608fae6fb24fc6bfb51fa06f9d6f7def6fcf542f59cf4a2f312f2beef9aec26e903e6b3e3c9e298e324e66dea11f03bf600fc450021028301f4fe6afb3df855f6e6f5bff611f8cef860f89cf6c8f3ccf08cee76ed92ed2cee39ee37ed3beb12e940e8f5e959eea9f432fbfafff001470145ffbffd01fe28001803d604b6035fffb3f88ef12eecd9e974ea0ded22f059f25af386f389f31df48af58ef7bdf99bfbdbfc9afd27feeefe6900c002ac0589084b0a020a6507ca0228fdcaf783f37cf06beeccec6aebb6ea48eb6fed0bf161f57bf9d9fc96ff470288056e09700db61070125812ca10540e6b0b2908440479ffeaf92df43cef05ecefeacdebffeda7f035f3a0f521f803fb6cfe2202b505bc08fe0a820c680dbf0d760d7b0cdb0af008400747063506a506c106ab05b802ddfdf6f754f24ceee9ec72ee42f238f72bfc47006303dd054108ed0ac40d391095114611360fd10bc107c303740010fe9ffc1cfc72fca1fdabff3d02da0400070a08a80736065404ba0219029a02d4033b055606f4063e077b07d7072708ef07e6061505b20243005efe2dfda4fcc8fc93fd2affbb011a05e908b50ced0f53120c141115411584149412600f560b0607f60291ffeafc02fbfdf902fa4cfbe4fd4c01dd04fc07140a0a0b340bdd0a5e0a260a620a2c0b840c030e380fd10f850f8b0e790d8c0ccb0b160bed090b08d705eb03e8024103bf04b50663082e090d096808a007220730078507d60721086008d408f209d90b630e1d112613e4135413b111b00f1e0e110d280cf90a0909740606047f024f027e036d05780767093d0b440dac0ff51167136f139f11520e9c0a7607b405cc0558079509ca0b200d420d870c6d0bb50a230bd20c690f521294147615c0146d12ec0e070b5e07a8048403f403bc058608810b140e3b10f7117f133315ef164518c318df1780151912270e560a440703059103fc021503d7035a0549075d098f0bb50dfa0fd5123d16d519191d131f0e1f041d3b195d14440f5e0afd057d02160049ff9d00e903a608f60d76122815ec15f114ea12d710390f480e2c0ebe0ef00fd4112d14a916d618ed19721950176f133f0e9b081f0382fea0fbd5fa3bfcb8ff8b04d209e40e231376163d19951b5f1d351e491d241a0715b30e8908f3039801a501d1032e07f90aa70e5b117512cf11540f7a0b4e07be039a018901a703c007430dfb1283179b198018c41425108b0c760b270d211048120312bb0e78094504d1000000b901dd043808fe0a910cb90c8f0b32093a06ba03b602e1032607580bf40ebf1032100e0ece0b830a8d0a770b0b0c660b9a0971072e06c6060d09fa0b250e530e4d0ce2084505b102d8017d02f3037e057706ae0651069f0511051405c1051b07eb088e0a6d0b470b140a32082d064b048e02de003fff26fe4afe3300f403b908ec0c2d0fce0ef10ba3074f03ebffdefd2cfd98fdf3fe2301e703af06a9081409c207240530022700e4ff6701ff037f06af07e9065004b80072fdbcfb28fc8efe2602c6057308c909fb098409dc082b082c076205b5028dff90fc88fa00faa6fa84fbc4fb03fb78f913f8ecf76ef92bfc31ff84019b02be02dc02ae0346053007a208cf08950776050d03c300abfe7ffc0ffa91f796f5dff401f607f971fd5702b106b9090b0ba50aed08690684037d0046fdaaf9c1f5ebf1b3eedaecdbec7dee10f1b1f39bf592f6ddf6fef68bf7cef8b7fa30fdfdffbb022405d00632072d062504b501aeffb2fea7feccfe0cfe83fb0ef761f1d1ebfbe7e2e6a9e8c7ecf4f1a6f6e3f92dfb76fa70f807f6edf3c4f2cdf2b7f330f5f5f6b6f881fa90fce6fe5a0176037904ca0314017cfce5f686f189edd0eb48ecebed7befbcef0dee1deb48e8bde643e789e943ec5dee59ef67efaeef61f1caf48df9bdfe21030f06700768076606c6049302e9ffd2fc3cf946f5f2f054ec11e8d6e411e325e3c2e4d7e68ae83ce9b0e8a7e722e7c2e71aea38ee66f3e8f8cafdc100fb003dfee0f85df2b8ec9ce901ea80ed6cf2e0f642f9dbf87bf698f37af11af161f234f48af583f59cf34df052ec2de887e4a7e17cdf6ddedadebae022e4b5e862ed69f167f431f64af744f81ef9b9f9b0f98bf87bf606f4b6f129f057efaaeee7ede4ec97eba3ea6deaafea14ebe6ea49e94de67ce287deb7db00db67dc9fdfcce3a1e780ea6eecdaedddef4ef31cf8a6fd8d023805ec049101a8fb97f4b3edcde7aae367e16de037e00de042df21de60ddc4dd3fe0eae4c0ea93f014f54cf786f7a2f672f5d3f4f6f454f57ef5e0f4e8f2acef72ebb1e688e202e0b2dfdee1bee5b6e985ec5ced23ec01ea5ae80ce878e902ec75ee19f0a2f04bf01df0f1f0f2f2e8f5d4f868fa15faddf75df4f8f0b0eea3ed70ed08ed5aeb6ee809e556e2bde1d9e323e88fedb4f260f637f854f83af7e7f506f5cff454f513f641f697f51ff442f2daf043f009f069ef73edc0e922e5fde0b2de25df06e23ae6dcea59efb4f36ff87dfd0e0233051c06b2040b02a9ffa3fe35ff5d006f0018fed6f860f186e948e348e05ae109e608edc1f475fbe2ffc601620167ffdefc66fa1ef807f6ecf39bf148ef64ed53ec58ec65ed38ef7ef1d5f313f64cf888fadbfc5fffef01510449066607550725060f048001fcfeadfc68fae3f7f2f4f1f1d3ef9deffcf1c8f6d5fc7c024d067c073a067f036a00dbfd39fc6cfb27fb21fb32fb79fb3afca9fdd2ff6202ad040206d305f803e8005dfdfaf941f77af5c1f454f577f71ffbd0ff94045308580aa40af0094e096609300a280b8c0bdb0a35091f072705b403be0207026a01e2009400ca009a01e5025e047b05ce054d0531040f03c002b903e0059508c10a730b840a81088206b7059506b808340bed0c390d3d0c800a9808d9061105e002230017fd98fad2f97afbbbff1f06630d12141a19c41bf91b4d1a73172f143911cf0eeb0c690bd409e407c505b9033a02da019902f0033405b1053a057b0478041b06ac094e0e7a12ad14f913c810a90c4e092908cb09550d4e116e14ba1520158813e111ec101111d61165121a127910990d4a0a530749057b049304f3043405380571059a061c09210d5d12bf174b1c5c1f3d20b51e2c1b1f167e10be0bee089208870aa90d9a108c124d137c130f142815351655168c14d410660cad08d606630796094d0cdf0e1411491314166b19d41c951fbf20fe1fa91d131ae315f311ad0e740ca00bce0b630ce40cb60ce40b470b920b460d86107b1406187c1a831b541ba91af51974192819aa18ce17a5161615661320127311ad1117131e15ed16de173417db14b411b30eaf0c2e0cdf0c330ecb0f4d11d312a31477160118fc18db189a17bf157913fd10b70eb60c350be20a2f0c570f2f14aa19871ebe217722ad20071d1c189d12390d3308110496010e019702f305240a450ef9110515b917901a3a1d111f811ff01d941a8a16ec128f10ae0f650f870e480c6808c8031b00d8fe0a01c906b30eba16cc1c1a1f111d8e1738104d09cb0479032f05f108170d8410e1121a14c0149d15bc16e117cd18e218b3175f153b12e90e390c910afa090d0aed090c096007340552035c0224022802f7015601f5001f02b205d00b8813ec1a66204f23b82374224020de1ca8174e102907d9fdcef6cff345f51bfa0c00ec04c007e008ab09890bf30e5d137417a519fb1856153f0f0508330120fc0bfa7ffbd4ffaf054e0bd80e8e0f170ebd0bed0990093b0aa00a9509b406b50228ff8efd8ffe98013c051d08700937093c085207b7065406e80532056c043304fb04e5068909ea0b050d4b0ccc0959063a037a018a01fb02a3046205a1047702aeff40fda7fbc5fa2dfa80f9dcf8f3f894fa22fe49030609ff0d0d11ba115910980d370ace067d03080043fc41f855f43bf1c9ef75f043f3bff7f2fcd101a7053b08cc09f20a4c0c1d0e1d10941191114a0f8d0add034cfc2ff5b4ef75ec7eeb6deca6ee94f1cbf4f8f7d4fa32fd12ffa3002e02ed03e805be07c0086908ac0601045c01cbffe4ff7901b80371058905600315ff6ef98ff3c0ee2dec57ecf3ee32f3e7f7ecfbbdfe7b00800122025602a501caff08fd2efa64f887f890faa6fd89002b0248025a01190017ff70fecffdc6fc0ffbb8f824f6b1f3b2f190f07ff06ff133f34af5eff6b3f78bf7c2f618f649f699f7f6f9f0fccdfffd010e03a102b900a6fddbf909f6d4f26ff0bbee70ed52ec97ebcaeb77ede7f0a4f5a0fae0fea301a6026e02a101830035ff93fd45fb56f80af59bf169eeb6eb82e9fbe755e79fe7f4e828eba3ede0ef7bf13af28ef249f31af565f8c8fc0b01c403bd037d00e4fa94f440ef50ec1beccaed2bf002f26cf290f129f0f6eeb4ee88efc2f08ff123f114ef06ec3ee9fde74ae935ed92f2def7b0fb2ffdb6fc50fbf2f94cf942f901f9e2f793f539f2b8eef4eb48ead7e945eae9ea80ebf5eb38ec8decfeec46ed68ed6ced4bed62edeeedbfeebfefb6f041f178f1a7f1f2f195f283f357f4eff443f56bf5f5f52df7cff872fa5bfbb4fa68f8daf495f07fec31e9b4e621e584e4e0e487e683e958ed60f1a9f460f69cf6d8f5a9f4c8f341f371f201f1e1ee47ec16eafbe8d8e848e9b7e9aae985e915ead9ebe1ee82f2a9f5ccf702f9f9f9adfb3afea900c001390098fb09f56aee61e918e765e7e6e84eeac9ea34ea6ce969e98feac2ec2eefc8f041f1eaf07ff01ef146f384f608fab6fc9cfdc7fccdfa4cf8e1f5acf346f16bee18ebbde749e56fe467e508e875eba0ee0cf189f24ff341f404f6b9f85ffc54006203ae04a703020050faa7f323edfce72ee535e51de84aed91f383f990fdb8fe28fde0f973f698f4f4f4def617f910fac3f88bf590f11aee39ec16ec03ed4fee82ef7ef0abf155f360f588f753f95bfac1fab8fa4dfaa7f9b9f859f7c3f578f4f3f38ef433f66cf8b1fa80fca6fd5efed1fe07ff02ff89fe79fd20fccefabbf916f98bf86af75af55cf2dbeecdeb10eaeee934eb3ded55ef3ff131f391f5a3f818fc3aff61013302ef01620135018e01240247025c0162ffbffcfaf98af779f588f39ef1e3efcfeefaee9bf074f3e4f60cfa57fce3fd0dff4a0004020d049a05e80582046f016afd97f9e9f6c4f5c9f517f6c7f56af46ef2e7f0fef079f347f866fe7a045a094e0c3f0d820c4d0aba06ef0130fc31f61af101ee78ed6cef07f302f73dfa14fc7ffc03fc65fb58fb3ffc0ffe7000df02e2044c063b07ff07ec082e0aaf0b310d4a0e8a0eaf0d7d0bcf07f2027cfd1ef8b8f3f9f0f3ef5df0ccf1c2f3eef547f8b4fae8fc8efe75ffb8ffbeff1a001e0195020d0440053c06a607610aac0ed8138b18ff1aed196a15940e09077e00f6fb76f985f878f897f873f8f4f748f7dff645f7eff8f3fbc2ff83037a063508f1088909bc0ad90cb50f9212a114791504158a138911300f770c5109890508012afc77f7aef3baf126f2f4f4acf93aff7004a708b10be50de60feb1191132214d4126d0fa20ac40551025201ac026a053408af096509ef073a064505c30560074a09dd0aa80bcc0b050cd60c4a0e0c105e11b1111811f40fd60e1e0e5f0dd20bea08860468ff19fbf9f8c9f963fd7b026907d70aef0be90ae3080d077f06e807f70ad40e8e1220151516b7157f1420134d121f126512df12e012d3118c0ffa0b8b0745032300dffeb5fff2018904a306cd0776089c09cd0b040f9d1255155d16e3159a149b13bb13a9146f150e15c712de0e830ad206a4043504c1046e05d905d205b2052c067b077509c70bdf0d780fcc102912f3134a168318b1190019e215d210350b84061d049a043807b20ae00dd30f8b10cd101f11ad113f121212ae106a0e140ccd0a770bee0d591183141f16b715a5137410f20cd90943073405cf03ee028a02c3027c03bd04d106ce09b70d4d12b916051a6a1b701a8217a913e60f310d050cdd0b000ce60b230b050a73090f0a170c3e0f5912311428143c124d0fc60cac0b5e0c670e8b109911cf10e20d6109530499ff2dfcf4fa43fc28005a06cc0d2915441b201f7320a61f441de919fd158111a40cef07f4037701070154029504e3064f08a3087e08a908e509840ce20fdc126f1407140112970f140e4c0e14101f12e51255113c0dbf07af0269ff8efee5ff71026905ae08640cc710a615dd19fb1b171b2e178a115f0c8c09d909970cc60f4011c90f730bc305d8002cfe32fe4700fb0218053e069e06c6063507dd077508d5081009ab09340ba80d881008133d14cf1317129d0ff80c990a7d089106f904d6034a036303e3038a044e054706a7077209350b530c4f0cfb0acf08b2065105f0046c053706cd06ff06cc065a06ca0514055004be039003f303d3049b05a2058a044a0260ffa4fcb7faeff957fab6fbe5fdea00a404b708a10cb50f611184116e10970e420c70090606fa0198fdc7f995f7a6f709fa14fe6a02ba054907f40646054d030002e301f802cd04a306b80792071d067f0301001afc49f805f5cff209f2a8f22cf4e3f52ff7ddf76bf8d2f9e2fcc001c507ae0d1d124b144f14ba122d100c0d4e09b9046cff08fa7ef5bef242f2ccf397f6c6f9a9fce6fe8f00e801f5027d03510336020c003ffd97fac4f83ef807f96bfa55fbf4fa09f925f67ef358f261f35cf654fa2efe0b01a70279031604c1046f05b805f304b70206ff37fa07f56ef05bed83ec0eee95f156f64dfba7ff2f03fc052508cd09ba0a490a1408180494fe44f813f2a0ec5be890e553e4a7e47fe6a2e9b2ed24f274f658fa80fdb9ff11015e01620054fe88fb50f864f56bf382f2a4f293f3c5f4d7f594f6d1f6a7f650f613f671f6c7f717fa2afd4b007a021d0309027eff43fcfbf8c5f57ff2d7ee8bea06e618e298df3cdf0ce165e495e8c2ec2ff0c5f287f455f56ff51ff58bf441f4e9f4caf611fa77fe0603a00639081107400396fd62f729f2efeef5edf1eedcf074f208f327f2b9ef66eccfe836e512e2b4df21ded1dd5adfefe28ae887ef8bf645fcb8ff8a006fff89fdc3fbd0faa8fa9cfa1efac2f855f637f3d9ef94ecffe961e89ce79ce7fde729e821e830e8cbe8c7ea71ee2af30ef8ecfb99fdfefccbfaeaf770f5e3f3f9f23df237f1b5ef48ee94eddbed0fef65f09cf00bef9eebe8e65ae251df77def3df0ee38be6b0e921ecebedd8ef90f213f628fa17fed700f60174019dff2ffda2fadbf7b5f4d0f0e3eb7fe6a6e149de64dd48df55e39fe805ee85f2ddf50ef825f96df9d7f818f764f416f19aedc6ea1ce979e8aee854e9e2e94deaabeaf2ea37eb56eb10eb9aea3aea41ea4beb81ed86f01df4caf7ecfa64fd21ffcdff44ff5dfdf3f969f580f023ec68e9c6e8f2e94deccdee75f01bf105f19ef081f0c2f0f7f0dbf029f0d2ee5fed3cec75eb30eb60ebd9ebd7ec99eefbf0b0f31af687f7cef733f752f608f6aaf6e1f728f9b9f9fbf829f7e8f4ecf2eaf113f2f9f2f7f353f4b3f379f258f124f1a7f2d0f5bff973fdcafffaff34fe25fb7bf7f9f311f1beee02ede7eb6deb84ebe4eb46ecb6ec73ed17ef67f283f7b7fdcf034e082f0a7f0910070804700165ff41fd59fa51f677f1f0ec06ea75e93feb9fee71f2cdf53bf8d6f909fb08fcd9fc6dfd8afd25fda4fc6ffcc7fcddfd90ff6301c40228032c02a9ffcafb32f7c5f245ef52ed3fedd4ee9af121f5eef89afce9ffac02cc046606ab07b0084709f3083007b603c6fe6af90df5daf263f36af6f5fac0ffa403d60518069004b70171fecbfb8bfafdfac1fcdffe320007008cfeb4fca2fb36fcabfe4702de058a08c0096a0905082306250462022801b2002e019702aa04de066f08d208ef070c06cd030e025401c1012d032c056e07e309700cef0e141125126111830ebe09e60351fe1bfae1f7b3f7faf8f8fa42fdbaff8a02f305c809800d5d108711a9103c0e260b9808b907fd08140c2110e1134e16f416d915a3132611b60e680c200a8307b2048402bd01dc02d905a509bd0c0a0e310de70aa40894072308e0097e0bcd0b6f0acb07f5042303f0025f04e8069c09f40bdc0d520fc410ba122215a517cd19ac1a96199a163912920d210ac0088b09ec0b8f0e38105b10f00e980c3e0a5208ee0606065c0500055a05a406f7080e0c140f6311c4123513331357139c13c31384137112b810150fef0d760d8a0d7a0dd40ce50b3d0ba30b860d2b1038127a123710f60b6d0768042304cf066c0b9b102a154c18001a9c1a241ac018b81622147611580fdd0de90c560cab0be10a810aee0a750c2a0f5a121a15bc16b5160b155212110fce0bf6089306c204b8038f03990410078e0a970e9e12cd15b2176c182d186917b21635160b163f167f169b168116e415b0140213c0100b0e2b0b1d081b05a002f5007e00a80159042508740c61103c13c514fb1457149213221356132c140b15531580142a129a0e9a0adb062204f5020c030004930571079409310c100fc211ce13ad14581459135912fc117d125813db137313b111c50e510bca07970411024b0076ffd1ff5001bc039f062109b00a310bd20a440a5e0a790b930d4d10ca125f14dc1447141a13091270116d11e61156122c12f3102e0eaa09a703bffc16f615f1e7ee40f007f53bfc8e04b20c76134d18241bfe1b3b1b7e19471711152c135d11400f8f0c300987054502e0ff88fe23fe42fe9cfe2dffe7ffb4007201f4015d022903e604f5070b0c21102f13a6149a14eb139a13e11331148313d910180c360696007efc88fa55fa0ffbfefbccfcb2fd29ff6c0158046c07e8093e0b3f0b1e0a86084507ec06bf076a09fc0a6d0b060ab00643023ffe21fcd7fc4f005c054a0a850d2c0e740c60092906c10363029a01cc00abff57fe74fdb7fd59ff0002eb044907a108f408a008110865075d06a8041302b0fefafaa9f769f5b7f4b0f51bf887fb53ffd902ae0596078308a30839088407cd0658063d065d0656069f05cc03db0066fd75faf2f830f9b5fa50fcc4fc8dfb20f9bef6c8f5e3f6acf9eefc46fffdff69ff92fea0fe3500ff02fc0514088e0861071a0558028cffe2fc3bfa77f7b6f443f286f0d4ef53f001f2a9f4e9f75ffba3fe4601180315044d0406048603d002e501c70045ff52fd19fbcbf8b7f652f5eef4a7f559f796f9cdfb67fdf5fd68fde4fbbaf982f7d1f5faf42ef53cf672f72df810f81ff7faf586f541f61df876fa52fc20fdf8fc72fc6cfc59fde3fe4400a50080ff1afd2ffa72f770f54ff4c8f39cf3aaf3c7f3e1f3d7f37bf3ecf27df291f2aff3fdf507f931fcb7fed3ff5fffaefd2efb8df85ff6c1f4a4f3def220f252f17ef0b4ef23efe7ee0befcfef5bf197f36df65ff990fb86fc21fc81fa5df86bf6daf4abf3bbf2c8f1f7f0b3f037f18df26cf448f6cff7cef832f934f9dff819f81df72ff661f5d6f43ef4d6f236f06eec04e83ae441e28be2f5e4c2e8e6ecd9f07ef4dff738fb70feed002702b5015fffa4fb5af758f385f04def61ef2df0d1f086f04bef9aed22ecb8eb98ec49ee47f0f5f1d8f231f360f379f3a9f3dcf3b2f327f368f295f123f169f166f212f424f6fef732f977f9b8f86cf70af6c5f4baf38af29af0e1edb7eac2e709e619e6b9e761ea29ed40efaff0dcf12ef32af5b0f7f2f954fb64fbedf987f710f521f332f252f20bf3d8f32ef4a7f359f294f0dbeeefed28ee6aef7ef1b5f347f503f6d7f5c6f442f385f178ef52ed43eb60e91ae8cde788e863ea39eda0f040f48cf7dbf9effaacfa43f976f7eef5ebf48af462f4baf355f252f011ee4aec78eb9beb7eecadedd9ee28f0b9f1a1f3eef518f876f9e7f969f934f805f73cf697f5e8f4eaf355f271f0baee6eeda7ec3eece9ebb1ebdbebd5ec10ef6ff26bf665fa97fd86ff50001300e8fe1afdbefaedf72ef5eef258f183f00df058ef2deea0ec1deb71ea21eb40ed9ff0a7f4a7f84bfc4eff7401c5022d038802fd00cffe50fcfef93cf84ef757f722f84ff973faf5fa69fad7f877f6dcf3e8f12ff1e0f1d8f358f661f850f9e6f876f7f2f547f501f636f847fb4bfea300020275025302ce01d8005bff59fd1efb3ef93cf84ef83ef977fa7dfb26fc8ffc26fd50fef9ffe001c4035405810676070608b307f105340271fc7cf5c5eee0e911e8b6e929ee0bf4cdf948feff003202c0029d035c052808a40bf90e551131126911560f850c5909f5052f02d8fd3bf91ef591f293f253f5dbf994fee001af023a01d8fe21fd3cfd66ffdb024e06a1086509e508d6070407f2068e077e085b09ab0938094d083c075d061d067d0601073907c8068c05f303b90269022d03a6041b06e206a8069f0557044303a5028f02d3025b03620406063f08e50a760d6b0f8510ad100210d20e3e0d600b76099f07f905aa048c0375028901fa0023017a02f404ff07e80af30cc80dbd0d640d490db00d480e870e1e0ef60c670b0f0a3a09ec08f708e9089308370815087908a209410be10c3e0e130f590f4d0ff50e460e5a0d3d0c390bdb0a4d0b600ca50d420ea20de60b84093607b3050405c704ab047a04810467056e075b0a820dc90f7a10c30f5c0e650dea0d15106e1321170e1a901bab1b861a99188f169d14d6124c11a70f8a0def0ac2073c0405019ffe62fd83fdc1feb7001b0396050308560a3e0c860d2c0e320e060e610e950fb71192144f173419091ac019c118cb172417be165c16581539131210210c0c08b8049402be011502fe02f303d1048b056606e907260af00c0110c512c914fa155e163716c915ed1480136011400e540a5006c80282003d00f2013d059d09100eb011271449153f15a214db1326139b12fa110711ab0fcc0d970b61094f07a005a3044e04a804b305130795084e0a260c2e0e991023135d15f31688171417f2156a14c4122e11700f6f0d4f0b1409f2062d05a3033c0221015300f5ff55006d01090314057307360a830d3d110d155918391a201a03182d14800f180bac07c20584057406fa07a309d50a500b520b0a0baf0a860a6e0a200a79095a08e00670055004aa0380039703c203f4032404820437051206e1067b0792072907a0064a068a06a0074e091f0b9e0c420de30cc20b250a5d08ab0609057c0341029001a801a10214045905dd054805cc030d02aa0017006f005b016d025f030104510464044004ff03b5035b030003a4021d027a01f700b500da007b0158022b03e40389043305f3059206a506e9057404c6028f014301d3019702a7027f0134ff66fc0dfaedf831f99cfab2fce5fee4008f02b6033004f1030d03ce01ac00080009008e004c01f7015b02650219027201680025fff3fd32fd3cfd19fe57ff3400f8ff58feb6fb12f9a2f73ef8e5fac3fe8802ed045105fa03bc018bff01fe15fd53fc41fbb6f90cf8ecf6d9f6eaf7c6f9c0fb39fdfcfd38fe5cfecefeafffd600dd014e02ec01b800e3fee0fc28fbfcf975f973f992f983f926f978f8a5f7e7f64af6cef57df570f5ebf532f749f9edfb95fe99009a019b01e000e3ffeffe00fe01fddefb9dfa8ef908f908f949f950f99bf81cf743f5c9f37af3b7f433f73bfaeafc76feabfec5fd31fc93fa70f9f6f83ef939fa87fbb4fc4cfddffc53fbe7f824f6d6f3b0f20af3fef427f8a7fb98fe2100b1ff7efd60fa6cf7cdf51df6f7f772fa70fc05fd1ffc6bfad9f859f855f97afb16fe45003001840058fe19fb90f779f43ef220f1fdf069f13df286f350f5c2f7bcfa9afda1ff32000effc4fc56fab4f892f8ebf9ecfb96fd0dfeddfc67fa8df72df507f44ef48af519f75bf8e5f8daf898f86ff8a7f82af98bf993f934f987f809f827f8edf837fa92fb58fc4efc88fb4ffa3ef9cbf8e9f858f9a2f93df915f86df6acf469f3f7f238f3ecf3b4f428f549f53ef539f59bf592f6fcf7c0f99afb20fd2cfebbfed1feacfe6ffeedfd01fd71fb0ef934f694f3daf1a5f111f37cf50bf8def95ffabaf992f894f75bf7faf7f9f8d7f920fa9af99bf8a2f70cf731f70ff83ff95bfaf1fa9bfa60f983f766f5acf3c2f2a8f241f33df435f529f658f7f1f81afb9efde2ff6101c201ff0087ffd4fd21fc9bfa3df9fcf720f7f2f674f78af8c0f977fa7afae0f9e0f8ccf7a7f615f5e9f256f0f1edc5ecadedc2f06df574fa74fea300e100a2ffd1fd40fc5cfb58fbfffbcefc55fd30fd21fc6bfa99f830f7a4f6f6f6a9f73bf855f8f9f7a9f7e3f7bbf8eef9e4fafefa3bfa1cf94af85bf854f996fa63fb2ffbf5f951f802f782f6f5f6f7f7e4f86ef989f950f91bf916f91df908f9b8f818f856f7acf638f61df65ff6f0f6dbf71df996fa29fcacfdf7fe26006401c302380458056905e2039400dbfbb0f62df20def98ed85ed3aee5defe1f0f2f2c8f535f995fc28ff5300e5ff6afec4fcaefb90fb4cfc45fdd2fd8dfd70fce3fa6ff98bf86cf8e3f897f942fab5faf5fa42fbbbfb3dfca7fcccfc84fcfafb75fb14fbcbfa6dfabef9bef8b6f718f749f75ef813fafffbc2fd33ff6d0089017502fd02c7027d0119ffd3fb02f81af48ef0c7ed36ec35eceaed3df1c0f5c7faa8ffc803b1061a08d707ee05db0270ffa5fc5dfbe6fba5fd66fff1ff95fe94fb18f8a2f53ff50ef745fa99fddaff8400e0ffa2fe8bfd1cfd4cfdadfdc9fd53fd33fca2fa05f9b7f7e3f67ff65ff666f6a9f688f78bf9fffc99016a06110a4c0ba109af05fc0055fdfafb03fd5aff5a019a0193ffecfb27f8daf5edf559f834fc1800da02fc03b103a5029701e9007d00f3ffe9fe46fd6ffb23fa0cfa6cfb01fe1101a5030c052805580445038d026a0295028e02e8019b0022ff40fe91fe2a0076026e041905f903570123fe72fb04fa12fa4ffb29fd28ff27012f0344053d07ce08a909a409ec08e807ed062206750592043503600149ff62fd4cfc77fc02fec20028045c0792093f0a4109f006f8031801ebfec5fdb5fd95fe1b00fc01ed039a05d706a4070b0826081d08f0079a073607e606de064207df074108f907b906a4046b02d80079006d0135030a055306d906ce06ac06ca062c078f0792070707140603053f042104a604b1052907da08960a410c9e0d760ec40e890ee50d110d0a0cb10af708d4067004350280008dff79ff1e004201bc025704e605480757080b098c09000a960a690b510c190da50dcc0d900d150d5e0c810bc20a4d0a520afd0a0e0c020d6a0dea0c760b7b097307be058a04b4030f03910245025a0206033904d705d007f209270c660e6310b91128128411fb0f1c0e6a0c430bb50a4b0a7909f1079905d4026100ccfe60fe2effd300d202e304cd068008240ad10b960d7b0f5411db12bf139f13601238107b0da90a35081f064f04d502be016a016902be04de07eb0ad00ce50c750b6409c6075a07fe07ed0844096e08a606c5048b03610323041105830565050205fa04f5050c08dc0ac90d15104c115c116810d80e2a0d9c0b510a4a0924089706b504b9023501f0003102b604e007b90a7e0c0e0db60c0a0c900b540b0f0b5d0ae408c60685049802780161010e022f039704fd055107bf083b0aa80bf50cd80d070e6b0d090c270a4808de063a066706f6066b077207db06e10500056d042d041d04ea0375030703f3028503d2047a0605082509b509f1093f0abe0a650b0b0c5b0c300cad0be90a010a1209fb07a8062e05a3033a023801ad009400d5002f017401a301ca012c0215037e0427069b073c08c5077e06fd0409043e0489055407de086d09d0086c07dd05bc046404b0044f05f60564069706b706d306f0060307d8064a064d05e30351020a017300e9008202cd0411078e089608ff0644042b018cfe11fdd7fc8cfdb4fedcffe9001202a303d1056f08e00a6b0c830cf40a2608f104290276001f00e10036029003630464049b033c02a70053ff8cfe6ffee2fe9fff74004d01340246038c04ce05c406380710077506b40506057904f4034a035a022a01daffa3feb8fd47fd7ffd6afecfff4b014b023802d90082fee1fbcdf9fef8acf995fb36feff00750340052406ec058a044802c9ffd4fd1cfdebfddbff1102ae03150435038b01bfff46fe4afda7fc15fc74fbeffad5fa62fba5fc69fe320083011f0208027101b9002900c0ff49ff6ffed5fc63fa5ff756f4fdf1f0f06bf13ff3e3f5abf81afbfdfc63fe92ffcd00160255035e04fc041805b304cd036702830032feabfb46f965f75bf63ef6e4f60ef85cf982fa76fb29fc75fc52fca3fb41fa56f84af67df459f328f3cbf3fff484f61af89ff910fb62fc80fd41fe9dfec3fee8fe3dffe7ffa300e20035005efe77fb2df85df5a3f353f335f48ff5b1f623f7c4f6eef52cf5dff445f540f66df789f86bf9fbf965fad4fa3dfb94fbc0fb93fb16fb6efabff942f917f938f999f90ffa64fa7dfa28fa3ef9e9f756f6b7f482f3f4f2e6f233f397f3b2f387f34ef32ef35ef3edf3a7f46af52af6eff6eaf733f9b0fa45fcb2fdaefe3eff67ff21ff8ffeb8fd8afc22fb8ef9c6f7ecf510f42bf271f009eff5ed5bed41ed8ded5eeec6efaef116f4c6f640f930fb5bfc97fc1afc37fb2dfa4ef9c8f89af8c9f83af9acf9f9f9e3f936f918f8baf65af572f437f47bf40ef588f565f594f451f300f252f1d0f192f371f6daf9f1fc12ffc7ffe6fed0fc1bfa53f718f5b2f3fdf2caf2cef2bdf2a6f2b6f20cf3d9f30ff562f6aaf7b6f85ff9d1f926fa5cfa93fac8fadafae3faebfaccfa8dfa14fa29f9d7f744f692f41cf326f2b8f1d9f164f21af3f0f3dff4e3f524f79bf816fa7bfb93fc21fd39fdfbfc76fce4fb5efbc7fa1bfa41f91bf8c4f662f50ef40cf37af248f27af2fbf2a3f38bf4c3f542f714f918fbf7fc77fe5eff7bffe5fec1fd39fc9ffa25f9d4f7c1f6d6f5e8f40ef477f367f341f424f6bff88ffbd1fdd5fe72fee8fcbbfaa2f816f733f6f6f532f6b2f680f79ff8eff959fb9efc6bfda6fd4bfd74fc7bfbb2fa44fa52fabbfa22fb38fbc1faaff94af8f0f6eaf574f57ef5caf53df6d4f6a0f7daf88afa79fc54feaeff3a000b006cffbefe69fe82feccfef0fe7cfe27fd1afbbcf893f638f5fcf4b9f509f75df83bf980f964f950f9b0f9a8fa0ffc9bfdfdfe17000a01f001c8026c037e03ac02f80098feeefb74f978f71cf672f574f50af61cf76af89df97cfafafa38fb88fb32fc50fdcafe5300990161028b0210020c01b8ff73fea9fdb0fda3fe3100a6014c02bf011b0013fe94fc2efcd0fccbfd1efe23fd02fba0f826f76bf76af93cfc99fe97ff23fff9fd33fdabfd7afffd014104810579057104e8025201ffff07ff75fe63feddfec6ffe700ea0182029e025402c9012d019f001d00aeff59ff1cffdbfe71fecafdf9fc41fc07fca1fc16fe250065025504b1058206d906d0068806fb0528054b04af038c03f603af042f05f504b0038001fffef0fc03fc8efc4efe9900a002a6035e0311025b0005ffcafef1ff42022905dc07c309b10acc0a890a5b0a460a040a4009ac0768051c037701f100a201fe022f04a1041d04e2029f01f50037015e020404b0050507c507ed07a407f506fe05ee04df031203e5027303b50486066208c8097e0a6f0ad10916098a084b08550866084a08ff078307e8065606ca054805f604e904430527067007e108400a350b8b0b380b320a9508b206d0045903b002d902a103bb04ac052f0663067906ba066c077e08c009140b3c0c160da90ddd0daa0d350d930ce80b540bac0ab3094b086a065f04c3020302530293033405aa06ab0710080408dd07b3079907ae07ef077a088309f70aa60c570e970f1510c80fb90e1f0d600bc5098808c0072f07840685050f046e0255015401c1028105c108810b100d1b0d010ca10aae098409190ae70a690b5f0bb90ab709ae08b407db063e06d105ae050706cb06d307fb08ed09840ade0a0f0b3c0b910bf70b460c620c240c8d0bbb0abb09af08c407f5065606f5059e0524056a044c03f601e2006e00df0049024b04710682086b0a580c760e8910141282125911c50e910ba208be062f067b06e606df061d06e204cd03430366031204d60456057f056505540593052406f406d3076e08a90898084c08fc07df07e707030825081608c7075c07e50683066b06a6063007f607bb0844096109e208cf075c06bc043b0320027c016601e801d70217048805de06e907a008fd08260955099a09ef09330a150a68092e088106b1041c03ef0146011b014101a1013d02f902c4038f042f059405db053306d306d8071109280ab70a6a0a4809a107d705520444038f021102af014e010a010c014901ac01220291020803b803bb040b0670077c08d1084c080b07790513042b03db02f0020603d4024202610186001d006500790130030f058906210791060805160367018e00bd00a201ab02470325036f0299010f011a01b30189024e03d70315041e040004b303270358025201490075ff07ff1dffb3ffa500ca01e302af030d04fb0390030703950247020c02b001f600c9ff43fea2fc47fb90fabffaf3fb1afeee000604d906e308d309910951088506a2040403cc01d400d5ff8ffee6fcfafa29f9daf764f7f6f77ef9b5fb3dfea8009802d4034404f9032f032a022e0170000000d2ffc7ffb3ff71ffeffe32fe67fdd4fcbbfc44fd5ffeb1ffc2002701ab0078ff06fed3fc42fc6afc0bfdbdfd25fe08fe70fda3fceefb9cfbd4fb7cfc58fd1dfe84fe75fe0bfe7afd02fdc4fcb0fc99fc45fc89fb71fa3af937f8c7f71ef82bf9b0fa47fc84fd3efe93fec2fe24ffe4ffcf007a016a014c0035fe9cfb17f93af74cf631f6a3f64df7f4f79cf85ef944fa4bfb43fcdffcf8fc8cfcbafbd4fa26fad3f9e7f93ffa9bfad5fad6fa96fa3bfaecf9bef9cef917fa7bfaeffa62fbc0fb18fc6ffcabfcb7fc77fcccfbc6fa95f96df88ff713f7e3f6e2f6f4f613f76ff735f879f933fb0efd82fe35ffeafea6fdd7fb04fa94f8d3f7b9f7eef723f816f8a9f711f79bf681f6e9f6bcf7b4f899f93cfa8ffac9fa14fb79fbf4fb4cfc29fc70fb2ffaa2f840f765f628f67df612f77bf784f729f78ef618f616f6acf6ecf79df955fbc4fc97fd92fdd0fc88fbf9f983f85cf784f6fbf5abf574f56af5a6f52bf6fdf6f1f7c3f84df978f954f930f93df97ff9f0f951fa4bfad1f9e8f8b0f785f6abf53af557f5f8f5e9f605f816f9e1f957fa77fa4afa02fabaf97ef97af9b9f92cfac9fa51fb68fbe7fac2f91ff882f660f5f2f44ff542f666f77df856f9dbf925fa40fa33fa28fa25fa1afa0cfadbf967f9d7f860f831f887f84ef925fac0fae7fa90fa0efaaff988f989f964f9d7f8fcf718f786f6a2f662f775f899f994fa56fb15fcddfc7afdb9fd54fd28fc82facef866f794f64ef65df6a7f618f7a7f76bf851f927fae3fa76fbdafb30fc68fc4bfcc4fbccfa7ef945f873f71ef73cf78bf7c8f7f7f736f8adf882f992fa84fb1ffc33fcbffb11fb6afaf0f9caf9e0f9f4f9e7f98df9c8f8caf7dbf64df685f6a0f769f98bfb86fdedfeb7ff070011001100f7ff78ff58fe71fce3f92ff7dcf450f3c6f220f30cf450f5b4f619f889f9fbfa53fc8bfd80fe04ff0cff8cfe91fd72fc9ffb76fb36fca5fd21ff0200cfff89fecbfc5bfbc4fa1ffbf1fb78fc37fc19fb7cf912f85ff782f755f871f975fa3afbb7fbf8fb21fc3afc4bfc7cfce0fc80fd69fe86ffa900b9018e02f302c602e2012c00c9fd08fb4bf805f682f4ddf30ef4f0f45cf63df871fac8fc0bffea001f0297025d02a001b000c9ff09ff86fe39fe09feeffddafdb8fd82fd2ffdbdfc3ffcc3fb5cfb29fb39fb92fb34fc05fdd9fd8afe00ff34ff43ff4aff4eff3affe1fe21fe05fdcafbdbfa9ffa41fba9fc85fe5f00cd019b02be0253029f01ea0073005f00a200f400fb006c003affa7fd37fc70fb99fb97fc02fe4cff0b002700daff81ff74ffd7ff8d005e0111028a02da02260390032004b6041c05180585046103db013700bffeb1fd2cfd27fd81fd03fe89fe05ff7bff0900cc00bf01c602b8036204b204c104aa0488046c043f04e0034c039c020402c9010902b4029303460481042c0451032c0210014000edff340004013c02a303d40470053905150445025700e6fe7efe68ff78013b04200789090d0b8d0b0c0bbb09f107f5050a0464020701e7ff06ff62fe18fe53fe17ff5200db01740304059a062e08ad09e10a5c0bd60a62095b07680542043a043d05ea069808bc09110a76090a081b06f5030402c3007000170190025904f4052007c8071c087608f10887090f0a360ace09eb08a90754064e05cf0407050c06a6077909260b310c650ce00bd40a8f0954081307b5054d04fb0225024d029b03e805d0089e0bc80d1b0f7e0f150f1d0ea30cbe0ab108b406220564048d048405050785088b09d8094409ff0787064705a404e304d5052c07a208eb09f70af30bda0c9a0d0f0ee40d000da00b150ad008340823084d086208050839076306e1050d061307a708500aa20b260cbd0ba50a2c09c507e3069a06dd0686073a08c50832097a09b509070a4e0a750a8b0a8c0a9d0afb0a9a0b530cf60c260db80cc70b6f0af2089e078406b0053f0521055905ff05f30618086209970a990b6b0cf90c4b0d8d0dbc0de00df60db60de60c790b71092c07540560049604ea05c30773098e0ae30aba0aa70afe0aca0bc90c5f0d120dd20bcb09810795055504dc032104d304b905c106cd07e0081a0a6a0bc00c080ef40e490ff80ef30d6b0cbc0a15099d076f066b058504da036c0350039f033b040505f205e206cc07ba089509490ad30a190b1d0bfa0aa90a2d0a880996085007da055004f602280207029a02cf035305cf060a08cb080b09f708b40872085d0866087008640817088c07f2066c061b0609060206ca05490579049303f602df0267037b04be05d6068607a3073e079206ce052305bb049304ab040a059d054b06f7065f074807a20689055404800361030804360560060107d706e805920457038f026002b30234039703b60389033603fa02f30224037003a20399035b030c03e702170395033904c4040105e50489041604b1036a032a03d60254029701b600ddff46ff28ff9dff8a00a4017d02ad020502a400eefe6efd94fc95fc62fdb5fe34009801b5027e03fc0337043a0409049903da02be013c0072fea3fc25fb51fa5efa34fb84fcdcfdcafe19ffdcfe51fecdfd91fda6fdf8fd62feb8feeefe08ff06fff4fedafeadfe6efe1afe9dfdfefc53fcc0fb8afbedfbe3fc33fe6bfffbff93ff3bfe43fc3dfab7f8f0f7f3f790f86cf94dfa0ffb96fbf3fb44fc9bfc1cfdd3fd96fe32ff65ffebfec9fd3dfc95fa39f96cf823f841f897f8e8f82df966f97bf960f9fff83af83df762f6fdf56af6bcf798f985fbfbfc85fd1bfdfbfb76fa04f9fef77cf78af708f897f8eef8caf8f8f7a6f62ef5dcf301f3b3f2bcf200f378f31ef426f59ff646f8cef9dafa11fb84fa7af933f80ef73ff6b5f56cf54cf517f5bcf433f468f394f2fbf1bef10bf2d6f2caf3b1f45ff5aaf5b7f5a9f576f52cf5c5f421f46bf3d5f273f276f2e1f277f31ef4baf421f56bf5abf5c8f5cdf5adf53df593f4ccf3ebf21ef27bf1e5f06ef026f002f02df0baf089f19df2e6f333f584f6bdf784f8a5f8ecf73df6faf3b8f1f2ef1def40efe3efa0f025f140f13af15cf1a9f120f292f2b6f2abf2b0f2e6f27af34bf4eaf423f5ecf454f4c3f384f389f3c8f305f4eaf371f3a3f27ef145f043efa9eedaeefbefc3f1d1f387f544f6f2f5d5f458f31df274f136f134f123f1c0f035f0bfef7eefadef56f048f17af2cff306f514f6e0f63ff749f712f793f6f4f541f562f46ef36bf23ff10bf0e5eedbed40ed58ed2deec5efd1f1bbf329f5edf50bf6f5f50ef65ff6d4f611f7a3f695f538f401f385f2f9f209f446f52af653f6e8f545f5b3f480f4a2f4c3f4b8f464f4c3f325f3caf2c3f229f3e5f3b8f490f553f6ddf643f792f7c6f707f85bf8a4f8ddf8f2f8c4f878f831f8f7f7e3f7e0f7b1f750f7c0f617f698f564f561f580f59ef5a7f5d2f557f640f783f8cef9acfaf1faa6fa03fa7df958f98cf900fa6ffa9afa8afa57fa1cfa06fa16fa29fa2afaf1f95cf989f8acf711f723f716f8c5f9d6fbaefdb3feb1fec2fd46fccffac2f943f95af9e1f9a8fa9afb90fc56fdc5fdb3fd0ffd08fce3faf3f990f9dcf9c4fa19fc81fda1fe4fff81ff5bff28ff16ff2cff4eff3cffc3feeefdeefc12fca9fbcefb67fc4dfd4efe54ff69008801930254037d03df028c01d0ff21fef2fc78fca6fc3cfde1fd5afea1fecffe19ffb1ffa300e00144039604ac056d06c706c4067706e30513050304ae02270198ff35fe48fd05fd78fd94fe2300d2015d038a043a05810590059a05d5054f06e6067807d907ed07c5076e07e606320643051604db02cd0123010d01830155025c036c046b0563064d071a08cc084d098a0987093009730862071506be04c3036703d3031305e906f408e30a540c050df90c3e0c040baa096c087507ee06c306d106ff061507e0065b0680057604a4035b03d6033e055d07de09800ced0eee107412491340136412ca10c40ee10c750b900a0a0a5c090d081106a1035401f8ff03008f0171040d08bd0b0f0f95111d13c513a713ff1234126a11a710ee0ffc0eac0d250c8d0a300966082b085508c9084609bf09620a2c0b0d0cfd0cb70d190e500e6f0e9b0efc0e5b0f780f3c0f830e6d0d610c960b3c0b840b480c5c0daf0ef90f0011b211ce113d112b10b00e0a0d9e0b850acf099709b209080aa70a640b1f0cdd0c700ddb0d600e140f10106411b5129d13e4134513ce11e50fce0de10b7e0aac096909b709470add0a6e0bd60b2e0cc20c920d890e8c0f39105f102a10b50f400f160f1a0f270f3b0f2a0ff40ebd0e5e0eb60dcd0c910b340a25098f0896085309850afb0ba50d390f81106811ac115311a910db0f190f850ed80ddb0ca00b430a2f09e9087809a20a090c120d790d6e0d240dee0c0b0d460d630d4c0de10c480cd60b900b6f0b680b340bc30a460ad2099509c509410af40adc0bc80ca20d660ecd0ea50eea0d8b0ccc0a2909ee0757077707f5077d08e208f508d008bd08ce081a09b709730a370bf70b700c770c010cf10a7609fb07cb06340662061b071208050990098c090a090e08dd06dd05490559051d0641076708450990095609e40864080508db07b1076a070d0792061f06e605d805eb0510060c06d1057205f60492048504d40474053d06cc06e30679069f05af041104eb033d04db046305a205990557051205f004d904ac044d04a203ce0214029d018c01e0016402f3027a03e103330479049a0488043a04a103de02230295015d018601e8015702a702ac0272021f02d701be01d301e201b60123011800c8fe85fda0fc63fce2fcf2fd54ffb400c1015f028d0262021102bb016e012f01f100a1003a00b3ff03ff3afe69fdabfc2efc00fc14fc4cfc78fc7cfc72fc80fccdfc63fd0dfe7cfe7cfefefd3cfd92fc43fc64fcdbfc64fdc9fdf6fde0fd92fd1efd84fcd7fb3cfbc9fa91fa93faa5faa8fa8ffa58fa19faecf9c8f9a9f990f979f97ef9b7f918fa8cfaf3fa20fb18fbf9fad7facffadefad4fa93fa15fa5ef9aef846f839f884f8f2f829f9fcf86ef8a5f702f7d4f61ff7c4f775f8cdf8b6f84cf8c0f762f75cf78ef7dbf71cf82af81df811f8f8f7cff772f7acf68ef552f441f3cbf230f351f4ecf58cf7a4f802f9b1f8e4f712f797f680f6c1f618f725f7d7f644f68ff50af5d2f4b0f471f4dbf3c8f285f182f006f04cf028f118f2cef22bf344f391f36cf4c6f569f7cff85cf9ecf8a7f7e8f557f468f327f380f30df43cf4d3f3ccf252f1f7ef34ef29efd6efdaf0a2f1f6f1d0f14ff1e6f0d8f019f1a5f150f2dbf25af3d4f334f48df4cff4d2f4b7f48ef44ef416f4d7f35ef3b5f2e2f1e6f00cf086ef5cefb2ef72f046f105f26ff249f2c4f120f18ef063f0a0f0f7f041f151f119f1f9f042f1fff12af35df403f5eef42df408f325f2e7f13ff2fff2a5f3a9f306f3ebf1a9f0c8ef83efb2ef38f0cdf026f15ef189f1a8f1e4f130f25cf279f285f26ff260f25af23ef22df22ff23cf281f2f9f26cf3d0f304f4e7f3b0f385f364f36cf37af34ef3eef260f2acf120f1dcf0d6f024f1aff143f2e8f284f3eef33cf46df472f46ef458f408f48af3dbf2fff14cf1fbf018f1bbf1aff29df36af4fff454f5a9f512f67af6e7f632f729f7e5f678f6eef585f545f509f5cef46cf4c5f308f367f208f229f2bbf272f321f48cf49af495f4c2f44bf556f6b4f701f901fa79fa4bfaadf9c9f8c2f7dbf62bf6b0f580f58df5baf517f6a1f64ef737f83ef923fac0faddfa61fa86f98af8a4f70df7b7f66ff624f6c7f568f551f5b0f590f6f3f798f927fb6afc27fd47fdf1fc54fca7fb35fb1dfb5afbe3fb81fceffc0afda8fcc0fb87fa3cf928f899f79ff714f8c9f87af901fa70fae2fa6afb18fccafc5bfdc7fd10fe48fe89febefec5fe8ffe1afe87fd1afdf6fc20fd86fdf8fd59feadfefafe43ff80ff83ff27ff6bfe68fd5efc9efb54fb8ffb41fc38fd4bfe5cff4a00030179019b016d010d01a1005e007000d90085014802e50237032a03b902ff0120014300a0ff63ff99ff3a001201d20144024c02f90188013901310186012502e702b0036304e2042a0534050605c70497049104cd043b05b005040604068e05b40497037402a10150018c01470238031604c40436058805f60590064a071208b40814093e093a090f09d1086808c307f5060e062e059004400439047e04ee04710504068106c606d006920631060a0661065f070209e20a7d0c7d0da50d0e0d1a0c0a0b0b0a37096b089807db063f06da05c505db05fc052c065f06a4062607d907ab089c097e0a370bcd0b220c320c240c040cf20b1b0c610c970ca00c440c7f0b960aaf09f8089a0866083208fd07b7078307b1074a0846098c0ab80b840ce80cdb0c8b0c4a0c220c140c220c170ce80bbb0b930b880bba0b010c430c7e0c850c4b0ce70b410b690a9909e6087d0892080709b509860a360bb10b180c660cb10c220d9f0d1a0e9b0ef00e020fe60e8a0e060e940d280db70c3a0c6a0b300abf083e0709069205e405ef068c08450ac50bf50cad0d030e3a0e5d0e820ec20eec0edf0e9f0e0e0e450d880ce30b680b250bdd0a720af90972090809fd0835098d09e709010adb09bb09c4091c0ad80aa90b4e0cb30cb60c780c400c0c0ce10bcc0baa0b880b940bc10b010c470c460ce30b3b0b560a5f099208e10751070607f5063607e207c608b409940a330b980bf60b4a0c930cd20ccb0c6e0cdb0b120b340a6a09a408ea076607180714076e07ea075a08ae08cd08d90815097f09090a980adc0abf0a680af2098a0955091f09bf082e086707a7064d066e060207d9078008b1086a08bc07fb0690069b0622070308d90855095709ca08e507090773064e069e0612075e075b07f1065106d00590059f05ee053606540651062e060706f705e405c305a1057b056d059005c905ff0521061c0606060d063106640687065806c405e504dc03eb024f0212023a02bc0266030e048e04b30481042504ce03b90303047e04ef042005f40493044604340461049b048604ed03dc028a015e00b2ff9fff1700ee00de01c1028003010440043f040004a2034603f702b5026f0205027c01f30092008300d0004d01c6010a02ff01bc0165011201d00091003f00e2ff8eff60ff73ffc3ff3300a200ef000a01fc00ce0087003200d9ff8cff6aff87ffe6ff75000401610170012b01ad002700b9ff71ff46ff16ffc4fe4bfeb0fd11fd92fc45fc33fc5efcb6fc35fdddfda3fe7bff5500040165016001e60010000eff0ffe40fdbafc6bfc3bfc15fceafbcbfbd7fb17fc89fc11fd7afda9fda0fd6efd45fd4bfd7dfdcdfd1efe45fe3efe19fedffda3fd6cfd1cfda8fc12fc58fba4fa24faf0f91ffaadfa6dfb39fce8fc4bfd60fd38fde4fc90fc5ffc4bfc54fc69fc66fc47fc12fcbffb67fb19fbcffa9ffa9cfabdfa06fb67fbadfbc2fba6fb5bfb17fb08fb2afb73fbc2fbdcfbc0fb85fb3bfb0bfbfffaf3fadcfab5fa72fa33fa12fafff9fdf908fa0afa1dfa5bfab7fa2ffba5fbdafbc0fb5cfbb4fa05fa84f93af940f992f905fa92fa27fb9afbe4fbf6fbaefb1afb52fa5ff97af8cdf758f735f763f7bef744f8e7f87ff90efa90faeafa2dfb5efb65fb4ffb24fbd6fa85fa48fa11faedf9d1f996f948f9f6f897f84df821f8f3f7d0f7bdf7b0f7d0f730f8b5f85df90efa8efadafaeafaa6fa2cfa9bf9faf87ef847f842f874f8c3f8f7f812f91bf90ef915f943f979f9b3f9d7f9b5f95ef9e8f85ef8f3f7c2f7aef7b7f7caf7c2f7bbf7d0f701f86bf807f9a0f92bfa94fab6faa5fa6dfafff982f90cf997f83ef800f8b4f765f71bf7d8f6d0f619f791f727f8aff8edf8f1f8daf8b9f8c4f80df96ff9e3f947fa61fa2dfaa8f9cbf8d5f705f77cf66cf6cef658f7e3f742f855f84af84df866f8aaf802f934f93ef924f9e2f8a7f883f85ff843f82ef811f814f84ef8aaf827f99df9cef9baf96bf9e8f86cf80ef8bcf77df743f7f3f6a9f679f65ef676f6c4f627f7a7f737f8b4f82df9a4f90bfa7cfaf4fa46fb61fb28fb81fa9ef9baf8fbf78ef764f73ef706f7b8f663f64ff6a5f649f71cf8d8f836f945f930f91ff953f9d3f96afaf2fa38fb0efb8afac5f9d3f8ecf72df79cf65af66ff6c7f669f73bf809f9bcf92ffa43fa12fac3f976f96af9b2f92dfabcfa24fb29fbd0fa31fa6ef9c9f861f829f81ef82bf836f858f8a0f805f987f907fa59fa80fa89fa81fa8cfaa6faa6fa7bfa1bfa8ef912f9d5f8dff830f9a3f908fa5afa9dfacefafffa29fb35fb31fb26fb19fb1cfb21fb04fbc2fa5efae5f987f958f949f952f95af952f953f973f9b8f930fac7fa60fbf9fb8bfc0bfd7ffdd8fdfffdf3fdacfd29fd80fcbdfbebfa2dfa95f92ef90cf92af979f9fcf9acfa7cfb66fc45fde8fd32fe13fe98fdfafc67fcfcfbc0fb9afb69fb2cfbf1fadafa0ffb98fb59fc2efde2fd57fe96feb0febdfed0fedffed4fea3fe47fecefd58fdf7fcb0fc7dfc47fcfefbabfb61fb3dfb64fbdcfb9efc92fd8dfe6aff110071008c0073003300e1ff91ff49ff09ffd0fe8dfe3cfedffd80fd36fd1bfd35fd82fdeefd59feb7fe07ff59ffc3ff5000ed007701c0019b010501170008ff1dfe93fd82fde4fd8ffe46ffe0ff4c009600e4005301e0017202d602de027f02d001fa003b00afff59ff2eff14fff7fee3fee7fe18ff91ff50003d013d022303c70323043a041a04e2039203190373029b01a600ccff39ff00ff28ff8afffeff80000e01b40185026b033e04e6044c057105790572055a052f05d4043e048a03cf022902b7016b0130010801eb00e40018018a0130020103d303830414057b05bf05fc052b063e063106e90559059c04c703050393028402da028c0361042305b90508061006fb05d505a9058b0560051705ba044604cb03760351036303bc034504e804a80566060b079e070408340841082108d6077b070b078e062506cc0584055a053005f304b204660421040d042c047d040f05c605950685076f083309c409f809c6095409b40803086b07e0065e060106c905c3050d068206fa0662078f0782076c075a075f079507dd0722086a08920885084e08d9073c07b9066e067506df067007f5076608b008ea084209a409f309220a0e0ac1097a093f090b09d208510872076d067705e4040305be05de0631085d09370acd0a0f0b030bd00a700af9099f095f0936092a090d09cb0881082c08e607d707eb0715085f08ac08f8085a09b209eb090a0aed0997093409c7086508380831085108ac081b098009d209df09a30952090009d608fc0849099009c009b1096e0933090809f60806090b09ed08c708910861085e0874089b08dd081b094b097f099b099e09a709a909ae09cc09de09cb099a093109a2082508c0077d076e07690760076e078e07d1075408ed087609df09fb09c90979091409b60885086f087208a308e508230958094d09ee0859089e07f20698069206d0064707bd07190864088a08840863081408a6074d0714070c0740078107b207da07e907f007090817080308d3077b071807e206db06f9062f0745072907f506b00675066206610663067206770672067606690643061306d2058e0568055a0561058a05c00504066506ca061e0751073d07de065c06d105690549055c057f05990580052e05c4045004e703a4037c036d038603ba030104550491049f04890453041e0415043a048904f6045e05aa05d705cf058a0512056a04ac03050388023e0225021a020a02f701df01cf01d601ee0115025802bb024303e8037c04cd04ba0438046a039502ea018701660163015c0149012d011c0127014a017801a601c801e001f9011202280231021c02e10184010d0188000b00a4ff67ff64ffa3ff1a00b3004501a901c301900122019c001f00c2ff89ff6fff6bff75ff87ff97ff97ff79ff3bffe7fe9bfe77fe90fee6fe65ffebff5c00a600bb009c004900c5ff26ff8afe10fed2fdd3fdf8fd20fe2afefefda5fd32fdb5fc4bfc0dfc0bfc5bfc06fdeefdeefec8ff39002d00aeffddfefefd43fdbefc79fc69fc73fc92fcbefce0fcf3fceafcb3fc62fc0cfcc1fb9efba6fbbffbdbfbecfbdffbcafbbdfbbafbd1fb01fc33fc6bfca5fccdfce8fcf0fcd3fca1fc60fc05fc9dfb28fb98fa0bfa9ff961f96df9b5f9fff929fa1bfacdf97af95af984f907facafa8bfb30fca3fcc7fcabfc56fcbafbf9fa31fa6ef9daf882f849f831f82ef826f82df84bf86bf89cf8def81ef970f9d6f92bfa6efa8afa63fa14fabdf962f92af917f905f9f6f8e2f8b1f87cf84cf80af8c4f780f72ef7f4f6edf60ef76af7f1f769f8c7f8fcf8edf8bcf884f83df806f8e7f7c4f7b4f7bff7caf7e8f712f822f821f811f8daf797f756f700f7b5f683f65af657f67af699f6b8f6d1f6cff6dbf610f758f7baf71bf83df827f8e6f77bf71cf7e3f6b3f692f677f63bf6fff5dcf5caf5edf54bf6b9f634f7a4f7d4f7cbf78ff714f791f62ef6e7f5ddf50ef649f68cf6c9f6d5f6c4f69ff652f604f6d2f5b3f5cdf528f694f60bf774f79df79af780f746f714f7f9f6d6f6c2f6c3f6bcf6c0f6c7f69ef64cf6dbf547f5d5f4b7f4e5f46ef535f6f0f68df7fff726f823f80bf8d2f7a0f78bf77cf784f799f78af763f72cf7d7f68bf655f615f6daf5b1f58ff5a8f515f6b3f675f730f89ff8c8f8bff884f844f811f8cef78bf754f719f7fbf607f718f734f757f766f783f7c3f70ff873f8e0f826f948f94bf91ff9e5f8b0f86df82df8f4f7a5f758f720f7f6f6fcf640f79df70ef87ff8c5f8f2f81ef948f991f901fa6afac2faf6fae2faa0fa48fadbf978f92ff9e3f89ef85df809f8b8f782f767f78bf702f8b3f89af99dfa80fb31fca3fcc0fc9efc56fce3fb60fbddfa4efac9f960f90cf9e3f8f0f81df971f9e6f959fac8fa29fb61fb7ffb95fba8fbd4fb23fc77fcbffce1fcbafc58fcd8fb4ffbe9fabcfabafaddfa1bfb58fb9dfbf0fb47fca7fc05fd42fd56fd43fd06fdbcfc83fc5ffc5afc6dfc7dfc87fc8dfc8efc9efccafc08fd57fdabfdeafd0efe18fe05fee6fdcffdc6fdd5fdf8fd1afe2ffe30fe19fef6fdd3fdadfd88fd66fd4bfd51fd8bfdfcfd94fe2bff92ffaeff81ff29ffd3fea4fea9fed9fe23ff6dffadffe0ff02000e00ffffd1ff89ff37fff1fed0fee5fe32ffa7ff25008800af0091003e00d8ff8bff75ff9affe4ff330069007c007c007d009000be00fb00380170019d01c701f601230240023d020902a0011a0193002f0012004000a9003501b6010e02370234021a020e021c0246028b02d10203031f031b03f902cc02990264023f022a02260243027602ae02eb0217032c0341035d038703cd0313043b0440041504ca038d036b036b038e03b103bb03b603a1038d039b03c203f50331045c046b0475047c048504a804d504fc04240537052d051e050a05fa040c0532055c058a059c0580054e050905c504ac04b704d6040c053a05520571059305ba05f7052d064a066006670668068506a906bf06ce06be068c065d062e06fb05db05be05a705be0501066206e3064f0783078e076f0737071407fb06df06d206c306b406c706f0061e075c078d07a707c707dd07dd07d907b9077c074e072e0721073e0764077c079a07b107c207ec0717082f08460849083a083f08480846084b083a081008f307e007d607f00712082b0850086a086c086b0852081b08f107d907dd071c087108b608ec08f108c808a40886086f0875087e088008a208d80819096b0998097c092e09b3082d08dc07ba07b107c307cc07c407d707030841089c08e8080d0926092e0930094d096d0979097e0962091f09d3087208fe07a6076e076407aa0719088a08ed081709fe08d10896085b0840082e081c082408380856089008c508dd08e708cf089e087908570837082c081e080608fb07eb07d207c907c007b507c507e30706083e086d0883088c0875083c08fe07b30761072a070607f9061c0754079007d50705081b0835084d086208810882085008f7077507e10670062406fd0505061d063e067806bd0603074d0779077c0772075c0751076a079307b607cc07b90777071d07a7062106a905460509050e0545059905020657068e06b706cd06d606de06cf06a4066d062b06e905b90588054d051105d004a104a504d7042a058e05db05030612060706ef05d505a70560051305c4048d0482049304ac04be04b1048c046504420429041c040904ed03da03d403e6031504490476049604a0049b048e046c043204e6038e03410317030e031c032b032103fb02ca029b0281028902a702d6020f03420365036e034c030103a0023e02fb01e401f0010d02280230022d02290223021a020202cf018b014d0127012d0158018e01b601bd019b0162011d01d7009b006d004f004f006b009d00d800060116010e01f700e000d400c6009d004d00d0ff3dffbdfe6efe5efe87fec7fefffe29ff41ff56ff7cffabffdbff020010000600f0ffc9ff96ff5cff12ffc0fe77fe34fefbfdccfd98fd62fd3bfd25fd29fd46fd63fd73fd76fd69fd60fd6ffd8efdb6fde0fdf3fdf4fdedfdd6fdb6fd8ffd54fd0dfdccfc8dfc5efc42fc25fc0afcf8fbeefbf8fb1efc47fc69fc7cfc70fc4ffc2cfcfffbcffba1fb65fb2afb03fbeafae8faf9fa00fbfbfaf3fae7faeffa19fb50fb8bfbc1fbd8fbdafbd4fbb9fb8cfb4cfbe5fa69faf5f98cf946f922f902f9e1f8c8f8b7f8d1f82bf9aef94cfaeafa5dfba5fbc8fbb7fb7dfb1bfb7efac1f908f961f8f1f7c1f7b4f7c4f7eaf713f850f8a8f8fef84ef98df9a7f9b2f9c6f9daf9f8f91afa1cfa06fadcf991f93af9daf860f8e3f774f717f7e5f6e6f6faf621f756f789f7d0f735f89bf8fdf84bf969f96ef970f969f96af968f93cf9ecf883f802f890f73cf7f5f6c4f6abf6a3f6c9f629f7a6f731f8abf8e3f8e3f8bcf876f838f813f8f4f7e5f7e1f7cdf7b6f79af765f72ef706f7edf6fef63df788f7dcf72ef869f8a4f8e8f818f933f922f9c9f843f8b6f735f7eef6e8f600f72ff762f77cf792f7a9f7b1f7baf7c4f7c0f7c5f7daf7ecf705f81bf818f80ef805f8f5f7f4f702f808f819f838f857f888f8c3f8e6f8f2f8def89ff855f814f8dcf7c2f7c2f7c2f7caf7d7f7d7f7ddf7e7f7e6f7ecf7fcf70ff839f879f8b2f8e8f80df90ef905f9fff8faf80bf92af93af942f93bf91af9f9f8ddf8b6f895f876f84ff83af83ef850f880f8c6f809f952f994f9b8f9c7f9bdf992f966f949f93af947f961f96bf96af960f94df951f96ff992f9baf9d5f9d5f9d2f9daf9e9f90efa3afa52fa5efa5cfa47fa37fa2cfa1afa0dfa01faedf9e2f9ddf9d4f9daf9f1f914fa56fab1fa0cfb62fb9ffbb2fbadfb97fb70fb4bfb20fbe2faa2fa64fa2cfa17fa24fa49fa8afad8fa22fb6dfbb1fbe1fb08fc25fc38fc56fc80fcaafcd4fce9fcd5fca2fc55fcfcfbb2fb80fb62fb5efb67fb6ffb7afb82fb84fb92fbaffbdefb2cfc91fcfefc70fdd7fd26fe65fe8dfe97fe89fe5dfe12febefd6cfd29fd06fdfdfc00fd09fd0afdf9fce2fcc4fca9fca4fcbafcf1fc50fdc6fd41feb2fe01ff27ff2fff24ff18ff1eff36ff56ff77ff86ff7aff5bff2bfff6fecdfeb2fea7feb0fec5fee3fe0bff32ff4fff5eff55ff35ff0affdefec5fecffefefe50ffbcff2d009800f200300152015e0155013f0127010d01f700e800db00cd00bb009d0076004d002a001c002f005e00a500f5003901690180017d0171016701640174019801c801050247028102b202d202d902c902a3026b0232020402ea01f00110023b026702880291028d0283027802780285029802b902e3020f03420373039603af03b803b103ac03aa03ab03b603c103c303c303bf03b503b303b303b003b203b503b903cc03eb03100440046a0482048c048604700462045c0462048004a904d004f5040a0509050305fb04f5040205150523052f052e0521051e052605370557056f057005620542051d050e051605300561059105b205cd05df05f00517064f068e06d40605070f07fc06c50675062a06e405a205720545051b0508050e0531057e05df054006a006ea061e0752077e07a307cb07e307e507e207d107b207930763071b07ce0679062a06fa05e205db05ec05ff0513063d067606bf0622078307d0070b0821081408ff07e207c907cb07da07ec0704080708ef07d007a80783077a077e078407920791078007790772076d077707760764075107370722072f0755078f07e30733087108a308b408a60890086f084e084908500860087d088a087f0867083708f507bb078307540744074307500776079c07ba07dd07f307ff0718082e0840085c086e0877088d08a408bc08e108f408ea08cd08910845080d08e307cc07d107d607d107cc07ba07a1079a0798079b07b207c807dc07fc0718083008560877089108ad08b3089e087e084a081208f207e107de07ec07ec07d507b40782074b072b07170710072107380755078607b707e8071d08410852085c08500833081408e807b6078f07650737070d07d606970666064106370653068106b406eb06100725073b0748074f075d0760075b075a074e0737071c07ee06b3067e064e062e062806270623061d060906ef05e005d405cc05ce05c805b905ad059c058d058c058a0589058e058c0585058405820585059905b105cc05e805f005e205c2058c0549050905c604860450041c04f003d203b803a4039603840373036f0376038f03bb03ea03180441045b046c04780478046b044e041804d00382033203ef02be02960276025a02390219020102f101ee01fb010f022a0247025b02660264024f022d020302d301a90189016f015b0148012e011301f700db00c700ba00af00a700a1009a009a00a100ad00be00c500b80091004e00f7ffa3ff5fff39ff37ff4bff62ff6dff5cff30fff5feb8fe86fe6bfe61fe68fe7efe99feb5fecffeddfedcfed0feb4fe8ffe6afe3efe10fee7fdbefd9dfd8efd83fd78fd63fd32fdebfca1fc5dfc38fc3efc5ffc8ffcbffcd6fcd3fcbbfc8cfc57fc2efc0cfcfdfb03fc0afc11fc14fc01fce0fbbcfb8dfb5efb37fb0bfbe6fad3fac7facefae5faf6fafdfaf9fadafaaefa83fa54fa31fa23fa1bfa1dfa25fa1cfa05fae8f9b9f98af969f947f92df91ef909f9fbf802f911f932f961f980f98cf984f958f920f9f0f8c0f8a6f8a5f8a1f89ff899f875f841f809f8c6f78ff773f760f762f777f784f796f7b1f7c1f7d5f7eef7f3f7ebf7d8f7a5f769f734f7fef6e2f6e7f6f5f610f72ff733f727f716f7f3f6d8f6cff6c5f6c5f6cef6c2f6b3f6a5f685f668f657f63cf628f61ff60bf6fcf5f4f5def5d2f5d8f5ddf5f2f513f61ff61ff616f6f5f5dbf5d7f5daf5f4f520f63af64af652f639f618f6f7f5c3f592f56af539f515f509f5fef409f52af543f560f577f56af550f539f51cf51cf542f571f5abf5e2f5f4f5f3f5e6f5bef596f574f541f515f5faf4e4f4edf416f53cf568f58ff590f582f56df546f52af523f520f536f565f58bf5b0f5c9f5b9f596f56df537f518f51af525f547f577f596f5b3f5cef5d2f5d5f5dcf5d1f5cdf5d4f5d6f5e9f50cf626f643f65af651f63bf61ef6eef5caf5b9f5abf5b6f5d5f5ebf506f622f62cf637f64af656f66ef693f6b1f6d9f60af72df752f772f773f765f74ff725f707f7fbf6f3f600f71cf731f74ef76ff77df786f788f774f767f76cf77cf7a9f7e9f71bf843f85bf857f853f85af860f876f896f8acf8c8f8e8f8fdf815f92af92bf927f920f90ff90cf918f928f949f973f995f9b7f9d1f9d5f9d0f9c9f9c0f9cef9f8f92ffa74fab3fad7fae9faecfadefad6fad7fad8fae1faeffafafa15fb3dfb6afba1fbd5fbf5fb08fc0bfcfefbf1fbe9fbe9fbfffb27fc53fc81fca4fcb0fcb2fcb2fcb5fccdfcf7fc27fd5bfd88fda4fdbafdc8fdd0fdd9fde0fde5fdf0fdfdfd0bfe20fe35fe46fe5dfe78fe94feb3fecbfedbfeedfe02ff22ff54ff8effc8fffaff140016000a00f6ffe9ffe9fff3ff09002800440058006600690068006a0074008f00be00f60037017801ae01dd0102021902280230022d02290226021f022102270229022c022b02250224022b0239025b028f02ca0212035b039603c703e703ef03f003eb03e003e003e603ec03f9030504090414041b0417041a041e041f04300450047704b304f304260554056f056f056c05620553055605630573059205ad05ba05c605c505b305ab05a505a005b305d205f305250658068106ae06d006e206f406fa06ee06e806df06cf06d606e406f10609071807130712070907fc0607071d07340760078907a107bf07d407db07ed07f707f5070008050801081208260832084b085808530853084a0839083d084308420852085b08570863086c086f0887089e08ac08cb08e408f0080c09200928093d094909430946093e092809220918090909100912090a0915091a091709270936093d09590970097c099609a709aa09bb09c109b809bb09b4099e099909910985099509a509ab09bc09bd09ac09a909a1099609a809b909c109dd09f309fc09120a1a0a100a0f0afd09dd09d209c509b709c609d509da09f009f909ef09ef09e109c909c809c609c209d609e509ed09080a190a190a230a1b0aff09ed09d309b509b409b709b909d109e309e709f809fa09ed09ed09df09c709c409be09b309b909b3099f09980984096909660960095509600968096c0986099a09a409b809bb09ac09a709940978096a0950092c091d090d09fe0808090e0909090b09fb08dd08ce08bc08ad08b808c208c708d908e008d908dc08cf08b608a9089208730864084f08390839083b083e0853085a0852084a082f080508e907cc07b407b207ae07aa07b407b407a907a70797077a0765074b07310728071d0712071607120709070a070007ec06dc06c106a20690067e0672067a067e067b067b066e065706450629060806ee05ce05b305aa05a1059a059d0593057e056b054e0530051d050705f104e504d704ce04d104cf04cb04ca04be04ab049a047f0464044e0434041d0411040504fa03f103db03bb03960368033b031a03fd02ea02e402e202e602f002f302f302ea02ce02ab0288026402470237022c0224021a020b02fc01e901cd01af01930174015b01470136012a011e010d01ff00f000db00c600ae008f00700052003500220013000400faffeaffd7ffc7ffb3ff9cff89ff72ff57ff41ff2cff1bff13ff09fffdfef5fee6fed3fec3feaffe98fe81fe60fe40fe27fe07fee6fdd1fdb8fd9ffd8dfd79fd65fd56fd41fd2efd25fd17fd0ffd0ffd06fdf8fce9fccdfcaefc96fc79fc60fc50fc39fc25fc1bfc0bfcfdfbf6fbe2fbcbfbb7fb97fb7bfb6cfb59fb48fb3cfb21fb05fbf0fad3fabafaadfa98fa88fa83fa75fa6cfa6dfa64fa5cfa58fa48fa3cfa36fa21fa0bfaf9f9d7f9b5f99ef97cf95ff94ff93af92df92cf91ff914f90ff9f7f8dff8cff8b5f8a5f8a4f89cf89bf8a2f896f88af885f86df853f841f822f808f8f9f7e2f7d4f7d3f7c4f7bbf7bcf7aaf79af793f77ff772f773f768f763f767f757f747f73df721f70af703f7f2f6ebf6edf6ddf6cef6c6f6aaf693f68af676f66ff675f66ef670f67ef67af67cf686f67af66df667f651f642f63ff62ef626f62bf61ef616f615f6fdf5e8f5dbf5bbf5a7f5a6f59ef5a4f5baf5bff5c8f5d4f5c9f5c1f5c2f5b2f5abf5b2f5abf5aef5b9f5b2f5aff5b4f5a4f59cf59ef590f588f588f577f56ff575f570f578f58bf58af586f582f56af55df562f55ef568f57df582f58ff5a4f5a5f5adf5bef5b9f5b5f5b7f5aaf5a5f5aaf5a2f5a4f5aff5aaf5aff5bcf5b2f5acf5aef5a2f5a3f5b3f5baf5cef5e7f5edf5fbf511f617f623f634f631f631f636f62df631f641f644f64df65af654f657f664f665f66ff680f682f68cf69df6a1f6adf6c4f6cff6e2f6fbf607f71af72ef72ff732f73bf737f73bf748f74cf75af76ff776f784f798f79df7a9f7b8f7baf7c5f7d8f7e6f702f827f83ff85af872f877f87ef889f889f893f8a6f8aff8bff8d8f8e9f8fdf811f918f924f92ff92df935f944f94cf95df977f98df9abf9cef9e5f9fbf90bfa0efa1afa2efa3efa5bfa80fa9dfabbfad7fae6faf6fa00fbfcfafafaf7faedfaf1fa02fb15fb34fb5afb7afb9cfbbdfbd4fbecfbfefb08fc17fc2bfc3dfc5bfc7cfc95fcabfcbafcbcfcc0fcc4fcc7fcd4fce7fcfafc19fd3cfd5bfd7afd96fda8fdb6fdc0fdc9fddefdf5fd09fe21fe36fe44fe54fe63fe6ffe7efe8bfe97fea8febdfed3fef0fe0dff29ff44ff59ff6aff7fff90ff9dffadffbfffd5fff1ff0a001e00300039003c0042004a00560067007a009000a900bf00d700f100040116012a013d014f016201730185019601a201b201c701d901ec01fd010802170226023102400250025c026b0279027f028b029d02ac02be02cf02dc02ee0201031103250338034403540364036e037d038d039903ab03bc03c403ce03d703d903e203ed03f203fd030904130426043704430458046d047a048b049a04a104ad04b904bd04c804d004d004d904e204e304eb04f304fa040a0517051e052f053e05440553056205670574057f0582058e0599059c05a705af05af05b605ba05ba05c705d705df05f005fc05fd05080610060f0619061f061e062806310636064706530654065a065a0653065b0662066406700678067806860691069506a206a806a306aa06af06ad06b506bb06ba06c206c906cb06db06e506e406ea06e706d706d906de06de06eb06f606fa060407070700070307ff06f306f606fa06fb060a071607190726072c0729073107320728072807220716071c072507280735073b07340735072d071e071b07150707070a070e0711072507330734073d073d072f072a0725071f07230720071507180718071007150716070d070d070707ff0607070b07080710071007040703070107f906f706ee06e106e106df06d706dd06de06d606d906d606cc06d006cf06c406c206bc06b106b406b506b106b306a80694068d06840678067c067f067b067e067d0677067c0679066f066f066706560652064f06460645064106360633062d06240623061606ff05f305e605d905df05e505e505ec05ed05e605e305dd05d205cf05c505b705b705b605b105b305ad059c058b0574055c055005410530052a052505200526052d052f053405300523051e0517050f050d050705fc04f804ef04df04d204bb049c0483046b045a045b045d045c04600460045f04630463045f04590447042f04210416040d040f040c04ff03f003d903be03aa03980386037a036f0367036a036c036a036903610355034f03490344034503400335032b031d030f030703fc02eb02d802c102aa029b028d02810278026a025c0254024d0248024802480246024702450242023e02340229021e020f02fd01f001e401d701c501af019c019001820176016f0167015c01550150014e014c01480143013b01310127011e0113010901ff00f200e800e300dd00d600ca00b800a4008f007e0072006a0062005c00590058005800560052004c0042003200230016000c0007000200fbfff4ffebffdfffd1ffc0ffadff9aff86ff74ff6aff65ff66ff6fff74ff73ff73ff6eff62ff55ff45ff36ff28ff1cff17ff17ff15ff11ff0cff00ffeefeddfeccfebefeb7feb1feaefeaefeabfea5fe9ffe93fe83fe75fe66fe5cfe58fe54fe52fe53fe4ffe4bfe4bfe4afe46fe43fe37fe2afe20fe15fe0cfe0afe04fefafdeffdddfdcafdbbfdaefda6fda4fd9ffd9ffda6fda8fdaafdaefdaafda3fd9dfd92fd89fd87fd83fd7efd79fd71fd6afd65fd5afd50fd49fd39fd29fd23fd1cfd1bfd21fd24fd23fd21fd16fd0efd0bfd04fdfefcfdfcf9fcf6fcfbfcfcfcfdfcfdfcf3fce7fcddfccdfcc0fcb9fcadfca6fca7fca3fca1fca5fca3fca0fc9ffc98fc94fc96fc97fc9efca9fcabfcadfcb2fcadfca4fc9afc86fc6ffc5efc4efc46fc48fc47fc48fc4cfc47fc44fc49fc4cfc54fc5dfc5dfc5efc64fc66fc6dfc78fc78fc6ffc67fc58fc49fc3efc2efc21fc19fc0efc0afc12fc18fc22fc2dfc2cfc2bfc2ffc30fc36fc3ffc3ffc3cfc3bfc37fc3afc43fc44fc42fc3efc2ffc1ffc17fc0ffc0cfc0cfc06fc07fc0ffc15fc1ffc2cfc2dfc28fc27fc22fc23fc29fc2bfc2dfc2ffc2efc31fc39fc39fc3afc38fc2afc1bfc13fc0bfc0dfc17fc1afc21fc2cfc34fc3bfc43fc40fc38fc2ffc22fc1cfc22fc29fc36fc43fc46fc4afc53fc55fc56fc54fc45fc36fc2bfc23fc2bfc41fc54fc65fc71fc70fc6afc62fc51fc40fc32fc26fc2afc3cfc4ffc67fc80fc87fc85fc81fc76fc6efc6bfc64fc60fc63fc6afc7afc8efc99fca1fca3fc94fc81fc77fc72fc74fc7dfc82fc8bfc98fc9ffca9fcb3fcaffca7fca1fc98fc94fc99fca2fcb3fcc5fccffcdbfce9fce9fce3fcdafcc6fcb3fca8fca3fcabfcbdfccbfcd8fce4fce8fcebfceffcebfce9fce8fce5fcecfcfdfc0dfd20fd30fd2ffd24fd17fd06fdfafcf2fce7fce3fceafcf2fc02fd18fd2bfd38fd3cfd34fd2efd30fd30fd35fd3dfd41fd46fd4dfd4dfd4dfd4cfd43fd39fd32fd2efd32fd3afd40fd48fd52fd54fd5afd63fd67fd68fd6afd66fd64fd67fd6afd75fd82fd86fd85fd85fd80fd7ffd80fd7efd7dfd7efd7afd7afd7efd80fd87fd8ffd90fd93fd9afda2fdabfdb6fdbbfdc0fdc7fdcbfdd0fdd5fdd2fdccfdc3fdb5fdaefdb0fdb5fdbffdcbfdd0fdd2fdd7fddafdddfde3fde8fdeefdf5fdfbfd06fe12fe19fe1afe19fe13fe10fe10fe10fe15fe1efe22fe25fe2afe2ffe35fe3cfe3ffe40fe41fe41fe45fe4bfe4ffe54fe5afe5efe62fe65fe67fe6dfe75fe7bfe82fe8dfe97fe9ffea4fea5fea2fe9dfe99fe9bfea4feaefeb7febefec2fec5fecafecdfed1fed4fed4fed5fedefee8fef4fefffe07ff09ff09ff06ff06ff0cff12ff17ff1dff26ff36ff47ff51ff55ff51ff45ff37ff32ff35ff3eff4eff5fff6fff7dff88ff92ff97ff95ff8fff88ff83ff86ff93ffa6ffbcffceffd9ffdfffe2ffdeffd3ffc5ffb8ffafffb0ffbbffd1fff1ff0e002100270026001e0015000f000e0014001d002e00480062007700840087007d006c005e005500500052005c006d0081009400a700b800bd00b500a600970093009e00b200cd00ea0002011501210123011b010e01fc00eb00e200e200ed00000116012a013a0145014a014c0147013f013901380142015b0179019501ac01b701b501ab019901860177016c0168016f0180019901b501cd01de01e601e201da01d601d301d301db01e501f00101021402250231023102270218020502f801f901fe0106021502250236024a025a026402690260025202490246024a0256026502730283028e0295029d029d02940288027a027202760281028e029f02ad02b602c102c802ca02cb02c602ba02b202af02b502c502d602e502f202f402f102ef02e802df02dd02dd02df02e902f80208031a03240328032a0325031d03180312030a03090309030c031a03290334033e033e03370332032c0327032b0333033b034803560362036e036f03640359034a033d033b033e0344034f0357035d036a037303750375036f0362035a0358035c03690374037a03810382037d037c0378036f036e036d036c03710376037a03810383037e037d037b037703770374036e037003730376038303910398039f039f03980391038903810382038403830387038803830381037a036e036603620363036e037a03840393039c039e03a303a20398038f03840377037103700372037d038603870386037e0371036b0365035f0362036a03720383039403990398038f037f03740368035f036203670369036f0373037203730371036703600356034b034b034d034e035803610366036d0370036c03690363035803500347033d033e033f033d03420345033f033a0335032b0325031f03160318031f03260333033c0340034503430337032b031c030903fd02f402ee02f502000306030c030c030303fd02f602ec02e702e302dd02e102e602e802ee02ee02e402dd02d402c402b902b102a802a602a802aa02b302be02c202c502bf02ad029f02930284027e027b0278027d02820285028c028c0281027602670252024202390235023a02450250025b025f025c0259024c02350226021b021102120218021e0225022802210218020802f101de01cb01b801b201b601bf01d201e301ec01ef01e701d501c301b0019d0194019101910198019f019d0197018a017701660155014301380130012c0132013c014701540159015001430132011b010801fa00f200f100f300f500fa00fa00f200ea00da00c300ae009b008b0081007d0080008a009400970096008e0080006f005f0050004700430042004400450041003c00310020000e00fcffe9ffdaffd0ffcaffc7ffc8ffcdffd3ffd6ffd5ffd0ffc5ffb6ffa9ff9eff94ff8cff87ff83ff7dff74ff68ff5dff50ff43ff38ff30ff2bff25ff21ff1fff1eff1dff1dff1dff1aff14ff0afffcfeedfedffed1fec6febdfeb9feb7feb4feb1feaefea5fe98fe8cfe7ffe73fe6bfe69fe6bfe6efe6dfe68fe62fe59fe4ffe48fe3dfe32fe29fe21fe1afe16fe11fe0cfe08fefdfdf1fdeafde2fdd7fdcdfdc3fdbcfdb8fdb5fdb5fdb8fdb6fdb1fdabfda0fd96fd8ffd86fd7ffd79fd70fd68fd65fd5efd55fd4efd46fd3ffd37fd2afd21fd1ffd1cfd1dfd23fd24fd24fd22fd17fd0bfdfffceefce0fcd8fccffccbfccdfccbfcc9fccbfcc7fcc3fcbffcb8fcb6fcb7fcb1fcacfcacfca6fca2fca0fc96fc89fc80fc73fc68fc61fc57fc54fc59fc5bfc60fc68fc66fc62fc5dfc52fc4cfc4efc4cfc4ffc55fc51fc4dfc4cfc42fc37fc30fc23fc18fc13fc0dfc0ffc18fc18fc1afc20fc20fc20fc21fc17fc11fc0ffc06fc02fc07fc0afc10fc18fc17fc14fc11fc03fcf9fbf3fbe9fbe5fbeafbebfbf1fbfcfbfffb02fc06fcfffbfafbfafbf2fbeffbf5fbf5fbfafb00fcfffbfdfbfcfbf1fbe8fbe3fbd8fbd8fbe0fbe0fbe4fbecfbeffbf4fbfcfbfbfbfbfbfcfbf4fbf0fbf1fbecfbedfbf3fbf4fbf9fb02fc03fc05fc05fcfbfbf5fbf3fbebfbedfbfafb01fc08fc0efc0dfc0ffc14fc11fc13fc17fc14fc15fc1afc19fc1cfc25fc28fc2ffc37fc36fc36fc39fc33fc2ffc30fc2ffc34fc3cfc3efc46fc51fc55fc5cfc66fc68fc6cfc71fc6ffc72fc78fc79fc7ffc89fc8cfc94fc9dfc9cfc98fc97fc91fc91fc97fc9efcadfcc0fccbfcd9fce6fce6fce7fceafce9fcecfcf2fcf3fcf8fcfffc02fd09fd14fd19fd21fd28fd28fd2cfd32fd34fd39fd43fd4bfd57fd65fd70fd7cfd85fd83fd81fd82fd81fd86fd91fd9afda5fdb1fdb9fdc4fdcefdd2fdd7fddbfdd8fdd6fdd8fdd9fde0fdeffdfefd11fe23fe2efe35fe37fe33fe32fe36fe3cfe4afe5bfe67fe71fe78fe7bfe7dfe7efe7dfe80fe87fe8cfe95fea2feaffebdfeccfed9fee4feebfeeefef1fef1feeffef1fef8fe00ff09ff15ff1fff27ff2fff35ff3cff44ff4cff56ff5fff67ff6fff78ff81ff8cff98ffa2ffa7ffa9ffa9ffa9ffabffb1ffbaffc6ffd5ffe4fff3ffffff08000e001100130016001c0022002900300037003c0043004b0053005a0062006b007300790080008b0093009b00a500ae00b500bb00c000c200c500cb00d400e100eb00f400fc00fe00ff00020106010b0114011c0124012c012f01310138013e0145014f0156015b0165016c01720178017c01800187018b018e019401970198019e01a201a801b301bb01c001c501c601c801d101da01e501f201f701f801fc01fc01fc010102030206020d0210021202160219021b022302290230023d0246024b0250025002510258025d0263026d02720273027802780276027902780278027e02820285028b028c028b02910294029802a202a802ad02b602bb02bf02c802cd02d202da02db02d802da02da02da02de02df02df02e302e102df02e302e402e602ed02ee02ee02f502fb0201030d03140316031b031d031d0322032303210322031e0319031b031a0317031c031e031f0327032c03310338033b033a033d033c033b033e033d0338033b033d033f0348034b034b034c03460340034203410341034603490349034d03500352035b035f035e035e03590350034c034603420347034d03540360036503640364035f0356035403530352035603570355035903590358035c035c03590358035603540359035c035d03620362035e035e035c0359035a03560350034f034e034d03500352035003510351034f0352035303510352034f03480345033f03360331032f032d03320337033a033e033d033603340331032d032e032d032803260323031e031c031a03150312030c030103fb02f802f602fb020003020305030303fc02f802f302ec02e802e202d902d402d002ca02c702c402be02bb02b802b302b302b002a802a2029e029a029c029f029e029c02940286027b0272026902660265026302620262025d025902520245023a022f0223021e021c021a021b021d021b021a02180211020a020202f601ed01e601dd01d701d201cb01c401be01b401ab01a3019a01950192018d018901870182017e017b0174016e0168015e01530148013a012f0127011e01180112010b0105010001fa00f400ef00e900e200dd00d600d100cf00ca00c100b700a9009b00900086007f007a0072006a0063005a0052004e00490044003f0037002b00200015000e000d000c000b0007000000f5ffe9ffddffd1ffc8ffbdffb2ffa9ffa0ff98ff91ff89ff7fff77ff6fff68ff63ff5eff57ff53ff50ff4eff4dff4bff44ff38ff28ff16ff07fffafeedfee3fedafed0fec8fec4fec2fec4fec7fec6fec3febefeb4feaafea0fe94fe8afe82fe77fe6efe66fe5bfe52fe4bfe43fe3cfe37fe30fe2cfe2afe26fe23fe21fe1afe12fe0afefefdf4fdebfde1fddafdd6fdcffdcbfdc9fdc4fdbffdbbfdb4fdaefdabfda4fd9dfd98fd90fd89fd85fd7dfd75fd6ffd64fd5dfd5bfd58fd58fd5dfd5cfd59fd58fd51fd4bfd48fd41fd3bfd36fd2afd1efd16fd0cfd05fd04fd01fd00fd03fd01fd02fd06fd06fd06fd08fd05fd01fd00fdf9fceffce6fcd6fcc7fcc1fcbcfcbdfcc5fcc9fcccfcd0fccffccefcd3fcd3fcd4fcd6fcd1fccafcc6fcbcfcb3fcaffca7fca2fca2fc9dfc9bfc9efc9ffca4fcaffcb4fcb7fcbbfcb5fcaefcacfca5fca1fca3fc9ffc9dfca0fc9dfc9bfc9dfc99fc97fc9afc9bfca0fcaafcaefcb2fcb8fcb7fcb5fcb6fcb0fca8fca4fc9afc94fc95fc94fc97fca3fcaafcb4fcc1fcc6fccafcd0fccefccdfcd1fccffccffcd3fcd2fcd1fcd5fcd3fcd3fcd7fcd7fcdafce5fcecfcf4fc00fd04fd07fd0efd10fd15fd1cfd1cfd19fd18fd12fd0ffd16fd1efd29fd39fd42fd4afd52fd55fd58fd60fd62fd64fd69fd68fd68fd6ffd75fd7efd8cfd91fd95fd9afd9afd9cfda5fdaafdaffdb7fdbafdbffdc9fdd1fddbfde9fdf1fdf9fd03fe07fe09fe0cfe08fe05fe07fe0afe12fe21fe2dfe3afe48fe50fe57fe5ffe62fe63fe66fe64fe63fe67fe69fe71fe7ffe8efe9ffeb3fec1feccfed4fed3fed0fecdfec6fec2fec4fec6fecdfed7fedffee7fef1fefbfe09ff1cff2bff38ff41ff43ff43ff45ff44ff44ff44ff40ff3cff3cff3eff46ff55ff65ff76ff89ff97ffa2ffaaffadffadffadffadffaeffb0ffb0ffb0ffb0ffb0ffb5ffbeffc9ffd5ffe1ffebfff4ffffff0b00170022002b003200360039003900370033002c00260021001f001e002100290036004a00610079008e009e00a900af00b000ae00a900a000940088007d00750076007e008d00a000b400c400d200db00e000e300e200dd00d600cf00c900c700ca00cd00d400db00e200ee00fb000901170122012601270125011d0114010801f900ef00ea00ec00f9000a011c012e013c014401480146013c01320126011b0119011d012601350143014c0150014c0140013401280120012201280131013e014b01560163016d0170016f016701570148013c0131012e012c012b01300136013f014d015c01680174017c017d017d01750165015501430130012601220121012b013b0150016a018201900196018f017b01660150013c0132012c0129012e01370140014e015b0164016e01750178017b017b0174016c0160014e013f012e011d0115011301170127013c014f0162016f017401790179017601760173016a01620158014b0144013b012e01220112010001f500f100f60008011f013901590176018e01a201aa01a2018f017001490125010201e000c800b600ad00b600cc00eb0014013b015d017d0192019a0198018501610136010701dd00c200b500b400c300d800f0000c01250137014501490141013601270116010e010a010701090109010601070109010e0116011c011a011701100108010301ff00f600ef00e700e200ea00fa000e012301300132012f01260117010701f300dd00d100d400e7000b01330150015c01530137011101e600bb009a00850082009800c200f9003401640180018a018101670144011c01f000cc00b200a600ac00bf00d800f4000b011a0125012b012c012c012a0124011f011a0113010e010a010301000100010501140129013f0153015e015c014f0138011801f800d800bd00ae00ae00bd00dd0005012d0152016c0179017f017d01740169015d014f014101330120010c01f700e000d000c800c800d300e500f900130130014c016b0187019b01aa01b301b401b101a7019101700143010b01d400a70087007e008b00aa00dc001b016101a901e90115022c0228020b02df01a80169012d01f500c600ab00a800ba00e000100142017401a301cc01ed01fd01f301d1019c015e012b010b01ff000a012301450170019d01c101d901da01c1019b0170014a0135012c012b0136014801610181019e01ae01b201a80197018f018f0194019b0199018c017d01710169016a016c016a0168016501620167016a016701610155014a014d015f017b01a201c701e101f201f301df01ba0182013a01f400bd00a000ac00d9001c016b01b201e70108020e02f701cb0189013e010001d800cd00e1000501290148015c01660171017a017d017e0178016e016a0166015a0143011701dd00a9008a008b00b300f20038017d01b301d601e601d701a4015601f400940054003b0049007700af00e2000e01290131012b010f01e500c000aa00b300e40029016e01a201af0193015601fc0090002000b3ff5aff2bff2fff68ffd3ff5300d20042019401c401d801c90197014e01ee0087002b00d9ff96ff65ff42ff33ff45ff74ffbeff19006c00ac00d800ec00ef00e700ca009a005e001700d5ffa8ff8aff7aff75ff71ff72ff81ff99ffb9ffdefff6ff00000300fcfff1ffe7ffd4ffbaffa0ff83ff6fff69ff69ff6aff6bff62ff56ff4dff46ff44ff4aff4fff58ff68ff77ff84ff8bff7dff59ff26ffe6feadfe87fe76fe7efe9cfec7fefefe3cff73ff9affa5ff86ff45ffeffe96fe51fe2dfe25fe36fe55fe74fe90fea7feb1feaefea0fe88fe74fe6ffe77fe89fe9afe9cfe8efe77fe5bfe44fe35fe25fe16fe0afe04fe0efe27fe41fe55fe57fe41fe1efef5fdc8fd9cfd71fd4afd32fd36fd59fd9ffdf9fd56feaafee9fe0aff0affe1fe88fe07fe6bfdcbfc45fcebfbc5fbd2fb07fc5bfccbfc51fde2fd71fee2fe21ff23ffe9fe81fe03fe83fd10fdbafc85fc74fc83fca3fcbffcc5fca7fc69fc24fcf1fbeefb2bfca2fc41fdf2fd96fe15ff5bff51fff2fe46fe61fd6cfc93fbf4faa3faa0fad8fa3cfbbdfb48fcd2fc51fdb4fdf5fd15fe14fefcfdd7fda1fd60fd16fdc4fc75fc32fcf9fbcefbaffb99fb95fbacfbdffb30fc94fcf2fc3bfd65fd68fd52fd30fd05fddefcbcfc9cfc83fc74fc69fc64fc5ffc4ffc38fc1efc05fcfafb02fc15fc35fc5ffc89fcbafcecfc10fd23fd1cfdf2fcb3fc6ffc2bfcfafbe2fbdefbf7fb2dfc75fccbfc19fd3ffd35fdf5fc86fc0bfca1fb57fb45fb6dfbc3fb42fcd3fc54fdb2fdd5fdb0fd55fdddfc5dfcf8fbb8fb9bfba4fbcbfb01fc47fc8efcc3fce5fceefcdafcc0fca9fc96fc95fca0fcadfcc0fcd3fcd8fcd3fcbdfc8cfc53fc1efcfafb02fc3afc93fc02fd69fda8fdb8fd94fd39fdc2fc42fccafb7bfb67fb90fbfcfb9afc43fde5fd5dfe94fe8efe4efedcfd53fdc5fc3cfcd3fb93fb7efb9efbecfb54fcd4fc56fdc1fd0efe2dfe12feccfd68fdf9fca5fc80fc91fce0fc59fddbfd54fea3feaefe74fef4fd36fd61fc98fbfffac4faf9fa96fb91fcbffde9fee8ff9100c3007e00c9ffb9fe84fd5afc69fbe0facffa29fbddfbbefc9afd55fed4fe0cff10fff4fecbfeb3feb1feb9fec6febffe8efe38fec0fd33fdb4fc5bfc38fc5cfcc2fc51fdf9fd9afe16ff6cff9affa3ff9eff8fff75ff54ff24ffdafe81fe19fea9fd45fdf7fcc4fcbbfcdafc1dfd86fd11feb4fe6eff3000e3007501ca01c4015d0195007cff3efe0bfd13fc87fb80fb00fcf6fc38fe8bffb9009001eb01c7013901650086ffd0fe61fe4cfe88fef8fe7dfff5ff43005a003300d3ff50ffc4fe4bfe06fe0afe5bfef5fec3ffa0006d0107024e023902c8010f0132005effbcfe70fe89fef9fea4ff5a00e600250104018900d8ff22ff99fe6afeaffe63ff6f00a501cb02ab031b04020464035f022101e3ffdffe3cfe12fe5bfefafec4ff8c00290185019f018501530127011a013b018a01f8016c02c902f202d6027402db0127017b00faffb8ffc2ff10008c001a019f0107024b026f027a0278026d0259023e021e02fc01e401e101f601230262029d02c402c302890218027c01cd003000cdffc2ff2600fb0028028303d004ca053c060d0640050404a1025f0181002f0065000a01eb01ca027603ce03c2036103ca0220029101410142019e014d023003230401059d05de05bd053c0575049003b002fd0196017e01ae0111027b02ce02f602ec02c2029b029302cb025503260425052b06f8065d073a0781064905ca033a02e100fcffa7ffefffc300ef013b036f045605dd050f06fd05cb05a00583057d058805860561050805660482037d027d01ba006d00ad008101d70275041e0693079008ee08a908c7077806ff0491036502a40152016f01f301bb02af03b804ab056c06e706fb06a406f305f904e603fa0263024d02d402e3035105e506450825095209a70836074905360373016e005a003f01ee02f504da063508b208400814077a05de03af0226025c024703a5042d06a007b1083909320998088b074006e004a303c302580275021f032b046f05be06da079a08ee08c2081e082607f605c104c8032903fe0251030104e704e405c4066b07d407f407d7079e0756071407ec06cf06b3069906730648062f062a063a0665068b0696067d062b06ac052405af047704a2042b05fa05f006ce076808b308a8085f080708b20772074f072e07fe06be0665060206b60589058405b105ff056406e0065807b607ed07de07850700076f060206ed053806d906b1077f0806092109ab08af0765060b05f3036a038c035504a6053a07c808150adc0af20a520a0c096107b8056904bc03d103810487059b067107e407f507b1073c07c7066b06410655069306e406330760075e073407e4067e061e06d005a405a805ce05ff0526062006e1057e051205ca04d2043305e205c306a4075a08ca08db088608d607d806a90579047203bc02730290020103aa0364041405a9050e0636061e06cb055305db047f0454045b047f04a904c904d804db04dd04dd04d504bc0480041b049003e9023e02b10166017d010302e80203041405d9052006d305fc04bf034d02da0098ffaefe37fe42fec9feb6ffe2001b023103fd0367046a0413047903bd02060270011101ef00f200f800d8006f00bdffe1fe0bfe7bfd58fda3fd42fefefe93ffd4ffabff1bff50fe86fdf7fcddfc52fd42fe86ffde00f901a102aa02f7019700b5fe93fc9dfa37f99af8daf8c3f9ecfafafbacfceffcf2fcf4fc1bfd80fd08fe6efe7dfe04fee8fc4efb7bf9bff785f613f670f687f70df99dfaf2fbe0fc49fd42fde3fc3bfc75fbb4fa06fa88f934f9e1f876f8dbf705f725f678f526f55bf50ff608f713f8f7f877f98df93bf983f893f79cf6bff53ef53bf5a6f56ef65af713f86ff850f8a5f799f65cf513f403f35ff234f29df28af3b7f4eef5e6f64cf70ff732f6c8f429f3b3f1acf073f02ff1b9f2d6f40cf7b5f866f9d7f8f6f624f4f2f0f0edd2eb08eba5eb93ed62f058f3dcf562f785f768f668f409f204f0deeec1eeb2ef5af123f3a0f46bf53af52af473f25ef06eee0aed60ec9eeca7ed1befb3f015f2ecf237f303f362f29cf1def02bf0a4ef44efe3ee8dee42eefaedeaed36eedaeeebef47f196f2a6f333f401f431f3f6f187f052ef94ee4cee7beeefee4fef83ef75ef11ef8bee07ee8bed42ed38ed5aedc8ed85ee7aefb1f006f22cf3fdf345f4d9f3ebf2baf17ef094ef1deffaee22ef6cefa7efe3ef23f048f05df049f0eaef67efe9ee91eea8ee3fef2af052f175f241f3a1f383f3d9f2e6f1ebf01cf0ccef0af09ff05cf1f3f11ef2f4f19ff148f137f17ff102f2c1f2a5f382f44ef5d9f5daf54bf539f4d9f2a4f1f2f0ccf027f1aff105f21df20af2f1f11ff2a5f267f35ef471f584f6a0f7a9f859f98af913f9e9f756f6a5f411f3e0f12df1faf073f1a5f27af4cef635f921fb3efc5efc8bfb26fa86f8e4f683f580f4ecf3f9f3b0f4e9f570f7def8d2f938fa26fad3f998f9a0f9e4f95ffaecfa60fbaffbb4fb40fb57fa14f9c5f7f0f6f8f6f2f7b2f9b5fb6afd8cfe11ff22ff09ffdafe73febbfd9cfc30fbd3f9dbf87af8c5f897f9b9fa0cfc6bfdb6fed5ffa5000d012001fa00bd0086004c00edff5bff92feabfdddfc4dfc11fc3efcdffc00feaeffc501eb03a6056f06ff05740442020b0066fe9bfdaafd65fe8affe8005f02bc03bb04110583041e0339015bff18fed8fdb6fe8d000803b6052908fb09da0aaa0a8009a8079405af0339025401fc002b01e9012f03d0047c06ba072408a2076b06f304c0031703f3022d0394031d04f3043706e107be09620b6a0cb60c4c0c580b1b0aac08160783052704540367036e0432064d082c0a610bcc0b730b830a4c09fe07cc060206c7052e0635078b08ce09c20a390b3f0b140bd30a870a460a040ad509f2095e0af90a8b0ba50b0c0bed09a108ad0793075f08ce09830bf80cd20d030e780d460cb70a09099e07f40633074708ed098b0ba80c270d0a0d930c290cdf0bb50bb20bb20bb90bf00b470ca60c020d160dca0c420c890bc50a300ac7099109b8092e0aed0af70b010dd00d5b0e840e5e0e2b0ee10d790d010d5d0ca50b290bf10af50a200b0c0b8e0ae50959096709810a780cd30e0611571275129311f00ffe0d4b0c020b4e0a640a1a0b420caa0dc50e2f0fd20e9f0de90b570a4d092709250af30b170e1e105511601164109e0ea80c490bc70a290b450c7c0d640ef50e240f250f470f660f590f1c0f8d0edc0d840d9f0d290ef70e6d0f230f2a0ea70c220b4d0a570a3c0bd60c960e10102211861137117310450feb0dd60c210cf10b740c6f0db70e3d109c118a12e6125c12ef100c0f090d690bb10acb0a7b0b890c800d440e150ff40fee10fd11ac12ac120412b810240fd50de90c660c4e0c4d0c4a0c7b0cdc0c890da50ee40f11112212d9122d134313f31235123011d50f4d0ef70ce20b390b390bc90be40c8f0e5e10e611d712b8128211ac0fac0d270cb40b490ca10d620fed10ea1163124c12d5114c11a910ed0f310f4c0e480d680cc10b8a0b090c1b0d920e4510c211ca125f135613b812a7110f100b0ef90b1e0af008e908010afc0b6a0e8310b811e8110f11970f230e0c0d990cef0cc10dc30eb60f2f1004104f0f210ecb0cbe0b210b160ba70b8a0c790d410e7f0e080eef0c480b790915087307c8071009d40aaa0c540ea00f9f10791105120b1255119e0fff0ce609bc06fe030a02e9009f003301870289041e07e7098e0cd40e73106411c3119111da10ac0ff40dbb0b24093a062f034b00d2fd2ffcd5fbeafc5affbb024a065a09820b990cd30c7f0cb70b830ae008d906c7042a0356025f02fc029503ba034e038002bd0158014c0165015f011e01d600e10078019a02f203ff046305fa04da035002a7001bffe5fd2ffd0efd86fd66fe54fffeff2500c9ff25ff7dfe00febdfd9afd7dfd6cfd79fdbdfd3bfec2fe10fff6fe5ffe68fd50fc3ffb52fa95f902f9a7f89af8cff829f97af989f956f91af915f981f956fa32fbabfb84fbbbfab1f9e0f87af87af892f858f8a7f7a3f686f5a3f425f4ecf3def3e8f3f5f31ff479f4f0f489f54bf61ff709f8e5f854f916f911f856f660f4aef269f189f0c2efb0ee6bed6bec38ec55edbbefb4f271f53ff7c3f756f78bf6b2f5f3f41af4c1f2f1f003ef66eda9ecf3ecd4edd2ee6bef3cef75ee76ed88ec14ec4aec08ed4deeeaef76f1c0f294f3bcf363f3b1f292f114f025eeafeb2ae940e772e62fe742e9c2ebe1ed0aef11ef9dee6deecbeec3efd0f026f184f008ef01ed18ebafe9ade815e8cfe7b8e70fe8f5e834eab4eb2bed2ceebeeeefeeaeee37eea0edcfecffeb57ebc5ea6fea4aea0ceac8e98fe953e954e995e9c7e9e7e9ede9cce9eee995ea9eebefec20ee99ee55ee7aed31ecfaea0cea37e986e8f1e75de71fe767e710e821e968ea85eb83ec62edf2ed4dee66eef8ed2bed1eeccbea89e986e8afe741e74de79fe749e829e9ece9aaea72eb2eec1ded38ee1cefb1efc7ef1feffeed98ecefea51e9e2e79be6dfe5f1e5c5e672e8b2eae8ecddee5df02ef18df186f1d9f099efc7ed6deb29e98ce7d6e657e7dce8c5eac4ec85eeb4ef82f002f113f1e5f07df0bcefddeef4eddbeccbebe2ea26eafbe984ea83ebdbec2eee0def9fef21f0b5f0b2f101f320f4cff4c6f4cbf32af21cf0afed42eb1ee97ae7f2e6dbe713ea69ed3df1abf450f7ecf861f90cf927f8acf6daf4caf27ff061eeb8ec9ceb5deb01ec43ed09eff6f085f290f304f4e3f3aff3ccf350f457f592f673f7caf779f77df640f5fff3bff2b7f1faf08bf0c0f0b5f131f3fef49cf679f78af7f5f6fef535f5daf4d1f410f55df575f575f570f565f58df5f2f57af636f701f88ff8d0f8b2f83af8cef7bcf714f8e0f8cff962fa71fae9f9d4f88cf73ff6f6f4e8f341f32bf305f4e8f595f8b4fba2feb800b2017a01280022febdfb35f9e8f610f5cbf352f3aef3c5f499f602f9bcfb8bfeff009a0227039b0239019aff38fe41fda9fc08fcf4fa68f9aaf739f6a6f520f675f753f957fb4dfd4bff5b015203df048105d804fe025d00a5fd8ffb7efa7bfa55fba4fc00fe20ffc1ffc6ff50ff9ffe17fe1dfed1fe080062016002b8027102c40102016400e2ff64ffdcfe59fe19fe5afe2fff7800ec0134032704c7041f053e050f0561041f0361017afff4fd46fda3fdfffefa001403ea043c06f30631071a07d00679061a069d05f7041004e702bc01d4007400c900aa01ba02a90338046e04a5042a0524068e0716095d0a390b8d0b570bb30a9109e507dd05b803e501f1001601420230044a060a083b09c409c30990095b0947098609040aa50a5b0be10b030cbe0bfb0ac4095b08d80667055704ca03e803e904af06fd089c0b1a0e2410ac119512de12ac12e0116710690ef60b4d09e706f904a903280355032104a805cb07680a680d5e10e712db14fa153816cf15c01424133d11130fce0cc50a0c09c10727073207e70766096f0bba0d1310fa1121139c136d13cc1225128211e9107610f90f690fff0eb00e8b0ec00e250fa60f5b100e11a1111f12461204129311fb1071104d106e10a010c7108610d60f260fc00e0e0f70109f12231594174919ef19a51964185e16fc135411a10e620cc50a080a760ad40be00d751017137f15af175f19721afb1ac01ab4191b18fd159f138711df0fdc0ec20e500f421076117a121e138f13cb13021488143815f015b0162a174d1755172c17cf1650166315f3134e1297102d0f890e950e250f251038115512c81389158c17b7196b1b2c1ce01b611af5173b157b120710400e120d800cb20c710da20e55103d122d142416c517e018791955197718261760154b133e11420f950da90c8e0c570d070f161104138e14551565152715c01458141414a713e612f411d210ca0f4c0f560fd20fa8106511c811de118b11ef105610bd0f3b0f0e0f260f860f48102111d7114c1222123f11de0f200e6c0c570b180bca0b650d5c0f291180120913d41244127e11ad10f20f100fec0dab0c5a0b3a0aa5099209f209b80a900b500c030d850dd30d070ef80da40d2e0d920cf20b930b740b980b060c7c0ccd0cf20cc20c460cb00b000b4b0ab2092209a30864086608bc0879095a0a1b0b880b560b800a4b09e907a006b4052305ec042505be05bf062e08c509310b270c4e0c990b440a9308ee06b5050105cf040d057105c305e805bf055905ea0491047404aa0412058a05f50527061206bf052c056f04ad0300038e027802ac020b036e039b037f032d03c80287029902ff02a3035a04e6041f05ff048d04eb0334036c0289017c003effecfdcafc1ffc30fc11fd98fe730039028d033e044904ce030403190227013a004dff62fe84fdc1fc2bfcd3fbb3fbc6fb09fc7dfc35fd3ffe90ff04015c023a035f03b402510187ffb6fd24fcfcfa38faa7f92af9baf868f86cf8f3f8f5f94cfba5fc9cfd02fed9fd42fd8dfcf8fb8dfb51fb36fb1ffb1bfb39fb6ffbbdfb03fc09fcc3fb3bfb78faacf9fbf861f8e8f78ef737f7f8f6dff6e1f611f770f7e0f765f8f0f856f990f990f93cf9b4f81cf880f711f7e3f6daf6fdf647f796f7f3f74df865f82ff89ff7b0f6b1f5f4f49bf4cbf462f5fcf565f677f61af68ef511f5abf479f46df450f425f4f2f3abf386f39cf3cff32af495f4d3f4edf4eef4c5f4a3f499f488f487f49af4a4f4caf40df52bf507f56bf41bf356f183ef07ee7bed21eeb5efe2f116f49df53af6eaf5c6f459f319f234f1eef03af1b6f13af28af260f2dbf118f118f020ef5aeebeed8fedeaedb3eefcef9ff131f38bf476f5aff55df5a3f47ef333f2dff06def15eefdec24eccdeb0eecafecaaedcdeeb1ef4ff09af073f01af0c1ef6def67efc2ef49f0fbf0acf103f208f2bdf10af130f052ef60ee94ed0bedb5eccfec66ed3dee4fef68f026f18af18ff11af166f090ef83ee7beda2ecfaebd1eb45ec1ced42ee6bef22f064f03cf0b1ef27efdaeebaeeedee69eff5efa5f06bf1fbf14ef23bf282f151f0e3ee62ed45ecd0ebebeb9beca2ed8eee49efc1efdeefeeef23f06cf0ddf04ef163f11ff188f0a6efe0ee7eee7deef8eec6ef82f014f161f149f10ef1dcf0a6f08cf07ef042f0f8efc5efb4ef0cf0d4f0bdf19ef235f33ef3edf27cf2fef1b0f189f142f1d9f049f093ef0cefecee2cefdcefd3f0b3f167f2def207f329f373f3dff37ff42ef593f5a2f557f5b4f40af48bf330f30ff314f30ef319f341f374f3c9f325f445f425f4c4f327f399f24bf242f299f23ef3f7f3c2f48cf52ef6b4f611f726f70ef7dcf699f685f6c2f647f71af80ef9d0f934fa09fa2df9d2f73bf6a4f469f3b8f286f2e1f2bef308f5caf6e4f8f8faa6fc73fd00fd6afb1df9b2f6e6f42ef499f402f608f833fa45fc06fe43ffeffff7ff49ff02fe4cfc5dfa90f82ff769f668f61ef74bf8a6f9d8faa4fb15fc5afcb0fc50fd32fe10ff99ff85ffc4fe9efd78fcaffb75fbb2fb1afc73fc9efcb0fceffc89fd7cfe97ff8100f100d9005900beff5dff66ffd6ff8600320198018c0101011a001bff4cfee7fdf4fd48fea2fed3fedffe08ff9dffc800680211043c0599052b0548046903db0299026b02040248017400f4ff2a004a0124033d050e071e08350873071e0690042f033202ab019601ce012d02a9023603cf0381043305c5052a065506550660069406f3067007ca07cd077e07f70676064e0691062007cb0742085b083008dd07870756073007ef0692061606a0057e05c8057a06840792085f09da09f909db09c809d309f8092f0a380aec096c09d90879089e084109220afc0a650b340ba30af4097b098009de09460a8a0a6d0afa098209360934098f090a0a730ad70a370bae0b710c550d100e620ef00dab0cf40a3409e80788070a082709930ace0b940cfe0c1a0d160d380d710da60dd60dcd0d7a0d090d7a0cdb0b560bd70a5f0a210a230a760a3f0b400c2a0dce0de40d730dde0c610c340c7d0cea0c1d0df60c4c0c490b630ad109bf09530a500b770cb10db60e610fc70fcf0f810f0c0f690ea20de90c340c930b350b020be40ae60ada0abc0abe0adb0a1a0b900bfb0b300c3d0c160cdd0bde0b170c7d0c140d9d0dfe0d580e970ebf0ee80ee00e850ee70dec0cac0b770a6909ae088708da088a098a0a7f0b2f0c960c970c4c0cff0bb90b870b880b8f0b8a0b980baf0bdd0b430cb30c080d3c0d180d8f0ccf0bd40abc09cb081208c0071608fd084f0adc0b2f0dff0d4f0e150e7d0dc80ce80bd00a92092b08d7060a06ee059106d90747096a0a190b380bfb0ac60aaf0ac30a010b2b0b250b0c0bdc0aa60a830a460ad3093c097808b107320705073007b6075908ef087409c109da09e509d909c209b0097609f7083e08420739067d0535057d0551065f0762083d09c509f809ef099709fe085208b5076707a5074b080f099609740992083b07ca05b1043f045304ad041005410550058105f605c206ce07ba08390929097d086b0750065c05b8047b048e04e60489055a064a073908d708eb085e082d0799050b04d5023f026002f702b60352048c0472044b045904d704c305cb068c07c20752078006b1052505ec04cf04680483033902e20005000700e5005802eb032605e5054a068d06e8065707950750074f06890453023300a5fe07fe67fe7dffe400310218039503cc03e90311043c043e04f4035b039702fb01ca011202a8022a033303a00294016b0093ff4aff86ff0d009200e70021017101fd01c70292030304d603f3028a010400c1fefbfdbafdd0fdfffd2afe4bfe82fe01ffd3ffde00e901a002c50253026a0156006affd3fe98fe9cfea7fe96fe69fe28fef0fdd8fdd1fdc3fd99fd42fdd9fc93fc97fc01fdcefdc7feb4ff6600ba00b6006e00e2ff18ff15fed7fc80fb4dfa6cf90cf93ef9d8f9b7fab6fbadfc8cfd48febcfed4fe87fecbfdc7fcaefbabfaf2f9a3f9b5f928fae9fac0fb83fc0afd2dfdf5fc82fce9fb55fbd7fa59faddf969f901f9c5f8c4f8e0f800f9fff8b9f847f8dcf7a5f7daf78cf893f9c9faf9fbe2fc6ffd96fd48fda0fcb5fb89fa3ef9e8f78af646f53ef48cf366f3e5f3f5f47af636f8c7f9f7faa3fbb5fb4efb8ffa82f94af8fbf6a0f572f4aff379f3fff339f5e2f6b8f864fa8ffb24fc1ffc7dfb68fafcf844f772f5bff356f27ff15df1e1f1faf26ff4e6f52ef720f895f8a1f860f8e5f76bf714f7dff6ddf602f729f749f754f72af7d3f64af685f5abf4e5f34ff323f371f319f404f5fdf5c4f651f79ef7a4f783f73ff7ccf63ff6a9f517f5bcf4b9f403f595f53df6b2f6daf6aaf624f681f5eff47df445f448f474f4dbf478f52cf6e6f677f7a6f778f707f776f60cf6e2f5e0f5eff5eaf5b5f577f55df57cf5ebf58af610f758f744f7d3f63df6b3f54bf525f53bf56bf5b4f50ff671f6f0f687f713f886f8b7f87af8daf7faf606f653f513f54df5fbf5e7f6c9f785f808f94af965f95cf917f992f8c3f7adf68cf5a2f41ef434f4e1f4f4f546f7a0f8cdf9c0fa68fbb0fba1fb3cfb88fab5f9e6f82ef8a6f74bf709f7ecf6fdf645f7ddf7b6f89bf95efacbfac0fa5afac5f931f9d6f8cbf805f980f923facbfa66fbcffbdffb95fbfdfa31fa70f9e9f8b4f8e9f880f95ffa6ffb85fc5bfdbffd85fda7fc64fb15fa17f9baf80ff9e7f901fb14fce7fc70fdb4fdbefda5fd71fd23fdcffc87fc5cfc69fcb0fc19fd86fdc7fdaefd2ffd5bfc5dfb83fa10fa24fac7fad8fb1efd6afe92ff7e002b0190019e015601b900caffa6fe70fd4efc6cfbe6facafa24fbe6fbf0fc22fe51ff52000c01730185015101ec006500d1ff44ffcffe86fe70fe84feaefed2fedcfecffec4feddfe3affdbff9d004e01c201df01b0015301e4007700060086fff8fe6ffe0bfef1fd37fedcfecbffdd00e401ba0242036e034203d8024e02c1013f01c5004600bbff2dffbafe88feaafe1effc3ff6d00f200450175019901c8010c025f02b302f902260338032503e3026c02cc0118017200f3ffa2ff71ff4bff24ff08ff21ff92ff7000a601f5021004b904ca04500470035c0242014a008eff23ff1eff83ff440043014a022803b403d60399031c038302f0017c012701e500a5005500f4ff96ff4eff39ff6effedffa90083015002f1025d039403b203d8030a043b044604f6032c03f401790006ffe9fd50fd4dfdd2fdb2fec5fff10015021c03f3037f04ad047604d903f002e901f1003900e6fffbff6500ff009601050243024d0234020c02d80198014b01eb0086003800180039009f002d01be0134027302800277026a026402600244020402ac015401260142019b010c02690283025002e7016101dd0073002000e6ffd0ffe3ff2a00ad005c012a020803db038c0405051f05c004e803a5022b01c7ffb7fe2dfe3ffed6feccfff50014020203ad0303040404c1034503a70208027a011501ef0000013a018f01e30124024f025b02510245023c02410262029102ba02ce02b0025e02f3018f015b017001bf01220277029802850261024b0257028b02c602ef02070313032e037003c603ff03eb035f0366024c01660004005600370158026503160452043e040404d503d003e503f903fc03db03a003710360037203a103c503bd037e030a0381021c02fc013002b50266031604af0419055605770578054b05ee0458049603da025602360297025e03570457052906b90610072a0700079006c905b20477034b02680105012c01d501f3025e04ec057107aa085c096a09ce08ab0753060b0505046b0339036303de0385043605dc054e0678066e063f060106cf05a70582056a0565058105d7055c06f1067707c207b9076f07f3066106de057805350525053e057805d5054406b40622077c07ae07b1076f07e9064306a0052d051a0569050206c5067e070608570866083008c40726076506b20531050b055e051206ee06b70727081a08a407ea06240697055b057205d4055b06e10656079f07b307a70781074b071807dc0689062806be05660550058405ef057106cc06dc06b306740650066d06b406f106fc06bb063e06c405730555055e055c053105ea04a3048604bc043a05de058c061907680774073307a906f60535058d042404f703eb03ee03ed03ee0315047104f7048905eb05f605b5054105c50469042a04f703cf03b603c50319049e042005660538059304b103dc02530235026302ab02f3022a035f03b30326049d04f204f4049104e50317035b02ea01d10106027302ea02410366034e030503ae025d021c02ef01c10189015a0148017001dd017102f8023f031d039f0202028101440153018601a901a00167011d01ed00e400f5000c010e01f900e400e600090143016e016a013401dc0086005200450050005b004f002800f7ffcdffb8ffc2ffe5ff1900530080008d0071002900ccff7cff53ff58ff7fffa7ffb7ffadff9cff9fffbbffd7ffd0ff89fffdfe50febafd65fd5dfd8afdccfd0ffe57feaffe22ffa6ff170050003d00e6ff6affe6fe6efe03fe98fd24fdabfc36fcdafbaffbcbfb40fc11fd29fe57ff5700e000ce002f0036ff2afe44fd8efcf7fb64fbcffa5bfa45fab4faacfbf4fc29fef1fe1fffb9fefdfd38fd99fc35fcfffbdbfbc0fbb8fbd1fb1bfc94fc19fd87fdc3fdb9fd73fd09fd8bfc10fca7fb4efb0cfbe2fac0faa3fa8ffa86faa1faf7fa84fb34fcdafc39fd35fdd5fc39fca4fb4dfb40fb75fbcffb1dfc45fc3efcfafb88fbf7fa55faccf982f97ff9c8f94dfae2fa72fbf3fb56fca0fcc5fca1fc2afc6ffb89fabbf942f930f97ff90bfa95fa07fb5bfb8dfbb1fbc9fbbdfb8afb38fbcafa65fa28fa0ffa20fa50fa81fab5faedfa0ffb1dfb0ffbd3fa79fa1bfac1f990f998f9c7f91bfa8afaf3fa50fb94fba1fb80fb36fbbbfa2cfaaaf939f9f6f8f2f822f98ff92cfacbfa5efbcefbf7fbe5fbaafb45fbd4fa66faedf97af91bf9ccf8b3f8e4f84cf9e4f990fa12fb56fb59fb18fbbefa6cfa22faeff9d0f9a3f978f963f965f997f9fef970faddfa2afb2efbf9faa2fa31fad7f9aef9a5f9c0f9e6f9e9f9d3f9b8f9a1f9b9f906fa5bfa9afaa2fa56fae8f993f96df994f9f4f945fa6ffa6afa32faf7f9d5f9b9f9a9f99df97ef96bf977f98ff9b7f9e1f9eef9f2f9fef909fa23fa43fa45fa37fa2ffa27fa37fa55fa4dfa15faacf91af9a7f884f8abf819f9a3f904fa2efa26faecf9adf986f971f989f9d3f934faa9fa15fb37fb06fb82fab2f9def843f8f0f7f9f751f8c7f85bf907fab5fa68fb02fc40fc0ffc6bfb61fa3ef948f89bf75af77df7dbf772f838f90bfae2fa9bfbfcfb00fcabfb09fb59fac8f95ff939f955f998f905fa8afaf6fa36fb30fbcdfa31fa8bf9fcf8bdf8dcf838f9c6f965fae9fa50fb92fba1fb94fb7bfb53fb32fb16fbe5faa4fa56fafbf9c3f9c6f9f6f94efaaefaecfa0cfb20fb3afb80fbedfb55fc9efcabfc66fcf4fb7efb20fb00fb1bfb51fb8efbb8fbb3fb91fb68fb4cfb63fbb1fb16fc78fcb0fc9efc5bfc0ffcdafbe6fb2efc88fcdafc0dfd1cfd26fd3efd5cfd78fd72fd30fdc9fc61fc20fc2cfc87fc0bfd98fd06fe37fe38fe1bfeeffdcffdc4fdcdfdedfd10fe20fe15feedfdadfd79fd70fd9dfdfbfd65feb3fed0febbfe8ffe7efea2fef7fe6bffd2ff0f001d000700e0ffb9ff8bff4eff03ffb6fe80fe7dfeaffe05ff5fff9dffb4ffb7ffbfffe3ff2d008c00ec003901620166014101ec007100e6ff6eff39ff65ffeaffa8005f01d401f401cb017c0139011e012b015e01a201e901330275029602850232029e01ea003e00c4ffa1ffd1ff4200e900b001840261032e04c4040705db04410464037602ab0136011a014701b1013602bd024703bf030e042f040d04a803230396022202ef0101024c02cc026103ec036804bb04db04db04c1049504720450041f04e60390032003bd027a026e02b9024703ff03d5049805270684069b066406fb056605bc042b04be0382038d03c003010451049204be04f20429055f05a705e50509061c061306f305de05c705aa0598057a054b052d05220534057e05e8055c06d9063b0771078a076d0715079e0602065605d70494049b0401059c054406ec066607a507c907cf07c307cf07e507fb0716080808b90740079c06f20595059c051106f106f107c70855096b0911098c08f4076d0726070607fd061a073f076507a607ea07230865089608b408e008020914092c092f091a0910090009e108c0087f081708b507640741077507d7074708c5082a097b09e2094b0a9a0abf0a820ade091a096208f5070d087d0804097c09a20972092309c60877085c085208480852085b0867089808de083809c2095f0a000ba40b080cfe0b860b8f0a3f09f507df062806fa052c069f064d071108e108cc099f0a350b860b670bdc0a210a4b097908dd0766070e07e806e106fc065007c2074a08f5089b09270a9c0acc0a9c0a1a0a41093708430780060606ed050c0645069c06f8065d07df075b08b208e008c2086108f7079f0776079007bb07cd07b6075b07ce064806dd05a305b205e8052d068606d2060807390757075f07600744070507af0632069a0511059e04570456048504cf0432059205e70540068e06cd06fc06f606ae0633068305bc0411049103490343036a03b3032404ab043b05c60520062a06e10546058204d303550316031a033d0366038d03a403ad03b003a3038a0375036a037903af03f503330451042f04cf035003d1027402520263028e02bb02ce02c202a5027a0250022d020502d901b801aa01bb01f5014c02ad0202033b03540349030f03a302070244017c00dbff83ff80ffc2ff25008300c700ee0006011d013b0163018e01ba01ea011d0242023e02f10148014b0019fff1fd13fda6fcb8fc3dfd12fe15ff28002901fc01810292021d022d01e6ff88fe53fd6efceffbd0fbfafb66fc15fdf6fdf9fefcffc2001c01f5004f0054ff37fe1ffd39fc98fb39fb21fb51fbadfb25fca8fc18fd71fdaffdc5fdb8fd85fd20fda2fc29fcc9fba6fbc2fbf3fb18fc0dfcb5fb2dfbabfa5bfa64fac3fa40fbb5fbf9fbf4fbc9fb9efb7bfb67fb4afbf5fa66fab2f9f1f85ff822f82ff87df8eef859f9bef91dfa69fab1faf3fa10fb0dfbe1fa71fac8f9f8f807f82bf796f665f6b7f67df774f86ef92dfa72fa4afad5f927f974f8dbf74ef7ddf68ff662f67bf6e6f680f72df8b1f8bdf853f88ff79cf6dcf59af5def5aaf6d0f7f9f8f0f983fa81fafff91cf9eaf7aef693f59bf4e8f38af378f3d2f3a5f4c5f516f756f826f971f939f997f8e2f759f7fdf6d8f6c7f68ff63df6f1f5bdf5d9f552f6e7f666f792f734f773f689f5acf432f441f4baf498f5bcf6e3f7faf8def94cfa3bfaa7f98ef830f7c6f56df461f3baf26af28df224f305f431f596f6fff765f9b0faa7fb2efc17fc2bfb87f962f7fdf4dcf260f1a9f0d7f0d5f155f32cf525f7edf868fa73fbddfbb8fb13fbf8f9a4f848f7f6f5e9f444f4fef330f4cef496f565f60af747f728f7d3f670f659f6bcf682f795f8aff96cfab0fa77fac4f9d8f8ebf709f75bf6f7f5cef5f6f564f6eaf674f7d6f7ddf7a6f759f70ef708f761f7eef791f81bf95af960f949f928f929f94bf95ef953f90ff975f8a7f7d2f612f6a9f5c3f55ff680f7fef882fad1fbb1fcecfc98fcd2fbabfa5ff911f8cdf6cbf537f51df59bf5acf61df8c6f96efbccfcbdfd1bfebcfdb1fc1efb38f974f73ff6ddf57ef604f800fafcfb82fd36fe14fe48fd19fce7faebf92ef9c4f8a7f8bff816f9aef96afa3efb16fcd3fc72fde3fd06fecffd2bfd15fcc8fa8df9a6f85df8ccf8d0f940fbe1fc70fec1ffa700f30095008dfff8fd29fc7dfa3ff9b6f8f4f8d7f934fbd0fc68fecfffe00075017a01e100aeff0ffe47fca7fa90f944f9d4f92ffb10fd0dffcb00010280025602b301d90008005dffd4fe55febbfdfefc4bfce9fb15fcf2fc67fe1b00a201a302f502a702eb01fe00120041ff96fe23fef2fd0afe6dfe11ffd7ffa2005901ea01460261023a02d2013a0193000600aeff96ffb9ff01005500ab000a017b01fd018802090363037b034703c402f801f900e4ffe3fe2cfeeefd48fe3dffb0006c022f04aa059e06dd064506dd04e302b900d8feb4fd8ffd66fef0ffb40142034d04b8049f044904ed03b403b103c803ca0393030d0345026d01c4008200c1006301340201039703ea031604280424040b04c3033a038302c5013e012d01ac01b60223049905be06580735075706f6045103b8017f00d1ffc4ff5c007601df026704c705c606420715074306040591033c0263012d0193016e026b034304d604150517050705e704ba049004600438043c046804ad04fd043405430534050605be046804fa03880348034e03a4033804b404c6046104a303ee02c5026103af045406ae074b080f081507bf058f04c7037b039f03ee032a043c040f04bc038903a50337044a059e06e207d0081e09c208e707a40611054f0369019aff5ffe33fe77ff3b02ed05a109630c690d900c5e0a990712055d0379021b02f901da01d5013e024b03fe0419070109220a300a12091e07fe04460364028c027a03af04a805ef056d057304740300038403ed04d606b408df09f209f1081707da04cd024d019900d600e8019b03b005ba075e09680aa20a060ac70808070105100380019f00ae0098011003ab04e0056d0674063e063906bb06a3078f081509c9089107c305cf03330255014501df01e9020404f804c3056406f906ab075b08c808b608e9076d06a9041e034802660234033404ef040a0596040b04d5033f045305b206e00782085d08760713067e040e031b02ca0129022503630480053b0669061a069d052a05e104cb04c604c104da042c05d305c3069b07e6075207c50592036a01eeff83ff4300d701bd038805e206ac07f007ad07f706f205b40470037402ec01f501a102ca03280565061607f60607068e0419034b0271027003d004d205ed051705af0354029f01b601540204035e034c031603100377034c043205c805e1058005e00457040704e603d3039a0325038a02f1018b017e01ca01560201039003dd03ec03d203b803d3032a049304ce049204c4038702270105006bff64ffdbffc000f90175032305b906c207ca0790063c046d01f6fe97fdabfdf7fed7009402a403e703ae03640352038403b5038403bd0276011b003fff4cff55000c02cb03e604ff0419049c0222012600d5ff07005b007a00510011001700b300e5015a038d04fc04720428039e016700eaff2b00d30064017501e200deffd4fe3efe6ffe6fff0401cb025104340547058e0432037e01c5ff55fe66fd14fd5efd29fe3eff60005401f0012a021c02f501e001f201210243022602ad01e70001003affc7fec2fe21ffb9ff5a00de0025012201d9005c00c6ff41fff5fefefe62ff0e00d8008b01f101e5015a015f0027fffffd38fd10fd99fdaefefaff2401e8012e020e02be0166011a01cc006400d1ff11ff37fe6bfdcefc78fc7afcd7fc77fd39fef5fe83ffdeff1b006200d8007b011c02720235024701d4ff37fecffcebfba4fbd7fb4efcd8fc5cfde1fd75fe1effd7ff8300f7001601d10023002cff1afe1cfd67fc20fc47fccdfc85fd35feb1fedbfeaafe36fea8fd2afdf2fc1cfda0fd64fe2dffafffbaff47ff73fe89fdd3fc79fc7dfcacfcb7fc72fcd7fb14fb8efaa8fa92fb49fd7cff9a0118038e03d00209019efe0bfcccf92af83af702f772f76ff8f0f9d7fbd6fd8dff9b00bd001000fcfe06fea1fde1fd67fea9fe27feb3fca8fab1f874f75ff772f83dfa36fce9fd09ff96ffadff66ffdffe2afe54fd83fcd7fb58fb0ffbf1fad9fac2fab1faaafac3fa0dfb80fb16fcb7fc37fd77fd60fdedfc55fcddfbbefb28fc04fdedfd7dfe64fe84fd15fc81fa2cf968f847f8aef88df9c9fa3cfccafd2efff4ffc8ff87fe5dfce9f9fef745f714f82afab8fccdfe98ffc2feb2fc42fa62f8d5f7ccf8cdfa1bfdf2fec9ff95ff9ffe44fde6fbb6fac1f925f9fef851f924fa3dfb2cfc98fc53fc71fb65fab9f9c5f9a1fa09fc74fd65fe89fecefd80fc04fbb4f9e8f8c0f814f9bdf98bfa49fbeefb82fc04fd7bfdcefdcbfd62fd90fc6afb3dfa52f9c9f8baf814f9a8f967fa49fb3bfc2ffdf4fd3bfed4fdb2fc07fb5af939f8f7f7acf80afa74fb6efcb6fc53fca1fb0dfbd1fafafa52fb7cfb47fba9fabef9e5f878f8acf8a0f934fb05fdaffec4ffebff17ff77fd5bfb37f967f71cf67df58cf533f673f73bf94dfb69fd3aff5e00a300ffff90feb1fcc3fa18f900f89bf7d0f77cf860f92ffad1fa46fb9dfb00fc80fc00fd5bfd5cfdd8fce6fbb2fa73f977f8eef7e3f76af882f90dfbe2fcacfef1ff49006cff5cfd8dfaabf76bf571f402f5eef6c3f9d5fc6fff1b01a0010801abfff6fd42fcdafad9f92ef9cbf89ef89bf8dcf86df944fa5efba3fce5fd03ffd3ff2300d4ffd0fe22fd17fb1af999f7faf65cf788f822fab8fbeefcb4fd30fe98fe1bffb7ff33004a00c1ff8dfeeffc47fbf0f93cf942f9dcf9d6faf5fbfafcc5fd44fe70fe55fe01fe85fd0afdabfc79fc8bfcdffc57fdd9fd43fe79fe80fe70fe65fe79fea5fec5feaffe4afea8fd10fdccfc07fdbdfda3fe44ff52ffc6fee0fd16fdd4fc46fd44fe66ff39007f0038009eff0affb2fe94fe8cfe64fef7fd5dfdd8fcb3fc1bfd06fe32ff4000da00e50089000c00b6ffb5fffeff5500850078003b000100f9ff33008900b4007700c6ffccfee9fd8bfdecfdf9fe6000a4015a025702bd01e4003100edff2c00c5007101f0011602cf01210129000afff0fd20fde7fc84fd0cff5501f2034206ad07d407ad068604f20184ff9ffd6dfce0fbcefb1cfcd1fc13fefeff73021d057207d408de089a0772050a030b01d5ff62ff62ff74ff60ff36ff36ffabffb60025029f03cf047a059a055a05de042f044a032902e200baff01ff00ffcbff2c01c9024404410590053b055304020389012b002cffcafe1dff1b0099014c03f1045a065c07e507f30776076f0602055803ab01450059ff04ff4eff23006701fc02a30423064707d407b3070407f705cb04c503fa026502f60198014e0139016201d1017e023703df038404340507060707f90782085108390762054b037f017a0073003201530279034c04bc04f104080511051505f904b7046c043b045504e204c805d306c3073d0812084a07fd056804e602b6010a0105019a01ac0218049705f9062008e20832092309b008ec070307070610053b048103d8024102b30150015401db01f50295045e06eb07020977095c09ee084b087e0788065305ff03e40252029202b4035105e306ff075608f90742078106e70584053405e604b004ab040505dd05f8060508b608b508f407b70654053304af03d1036c043505c305e905c5058b0590051306e2069d07e2075c071d06a90493034c03f70332056b06240715076e06af0537053d05c0055f06bd06c4067d0626060f064306a006e306b60605060b052104c2034d04a8056a070c09e6099d0955087906a90477031b0380035e044505fe058c06ed062f0759073b07b506db05d404e803610350039a0316048504d7041d0554058505b505c405b105a905c3051206920606072207bd06d605ae04b203310365035204a705fe0600085408dd07cf06770538047203340357039803b303a803bc0334044105bf061a08ab08210889067404b802eb012902160308047f046304ef039d03d1038604760542068d063d067e0586049303db0275026902b9024803f0038a04f0042505450559055d053c05c204df03c702d3016801c601d00226044f05e805df056d05db0464041e04e8039d033503b9024a020b02fb01010207020202fd0113025002b60232039b03d303d50399031f036f028f019800b9ff2cff25ffbcffd1001b024203f9032804ea0377030f03d502bc0294022a025f0143001bff47fe23fed8fe48001102ad03a004aa04e1039f025d018000300052009d00be008000deff02ff2efea4fd93fd05fed9fed5ffb7004901770151010101b0006b001c00a3ffedfefffd0afd48fce1fbdafb17fc7afc05fdd3fdfdfe82001d024d039203a402a60026fee5fb84fa54fa2bfb83fcc4fd7afe78fef4fd53fd00fd57fd69fefaff9b01c202ee02e501bfffe0fcebf97df707f6cef5cdf6bbf83ffbe0fd12006901a301ba000cff21fd83fb8ffa45fa47fa2cfaaaf9c3f8e7f7a2f759f82cfac1fc5aff4101ee01300152ffe3fc83fac3f8e1f7d1f76af866f97ffa9ffbb9fcaafd56fe8ffe24fe1ffdb2fb2bfaeff83cf810f851f8c4f833f9a6f92efacefa94fb60fce6fcfbfc89fc96fb60fa2cf930f897f75bf74ff759f759f740f744f7a4f787f807faf6fbd5fd22ff6dff7cfe8bfc15faa9f7d2f5cff48ff4f7f4d1f5e9f645f8dbf97bfbf7fc0efe77fe26fe32fdcffb54fa04f905f881f775f7b4f71df871f868f803f86bf7e3f6d9f690f7f0f8acfa3efc17fdfcfcedfb25fa28f861f60ff574f49ff46bf5b6f63ef89cf987facffa65fa88f985f89bf710f7f5f62bf7aef768f833f90bfad7fa60fb93fb67fbd7fa12fa40f96bf8a7f7edf62df698f564f5bdf5daf6a9f8c0faa7fcdffd04fe21fd85fba0f902f800f79df6c1f61ff758f751f70bf79df659f67ff61df735f892f9cdfa9bfbc3fb2efb17fad2f8acf701f7f3f65df71df8f2f88af9cef9b1f934f989f8e9f77ff78ff733f84af9a8faf9fbd5fc16fdbbfce4fbebfa17fa7ff92ff908f9d2f880f815f89cf750f760f7ddf7ddf849fadafb4afd43fe73fec5fd4cfc3afafcf7faf582f4e1f332f456f521f741f947fbe2fcd4fdf9fd6dfd61fc11fbd2f9e3f861f867f8e7f8a9f985fa48fbc2fbf7fbfbfbe1fbcdfbd2fbe6fb07fc23fc1ffcfefbb7fb41fbb9fa43fafbf917fab3fab6fbf5fc23fee6fe0eff8ffe83fd35fce8faccf90cf9b2f8aef803f9a7f97ffa75fb6afc36fdc7fd1afe38fe37fe1cfed7fd61fda6fca7fb94faaff932f959f931fa89fb19fd88fe87fff6ffe0ff74fff9fe9cfe66fe46fe0cfe89fdc5fcf0fb58fb56fb1bfc8ffd59fffa00fa0117025301f5ff6afe0efd1bfca8fb9ffbdbfb45fccdfc68fd11fec4fe75ff17009600df00d900690088ff4ffef2fcbefb0afb14fbeafb6cfd53ff3b01be0291039103ca027e011500f8fe6afe77feeefe73ffb8ffa0ff50ff17ff41fff2ff150156025a03e303dd035f039b02bc01dd00120067ffe9feabfeb3fefbfe73ff03009a003601cd015202b902e302ba0247029c01d80022008eff29ff04ff2bffb3ffa900ee013b034204ab04560470034e025d01f5001f01ac015802d9020a030003da02bb02c102e1020e034b038f03dc033e04a104ea040805e4047904e5033d03a402430222023d028b02e5022b035703590340033103360357039d03f0033b047c04a504b804c804cb04bb0499044704b503f7021f026101100159014e02de03a9053e074b08940824084c075b0699053705170510050705da048c044d0437046004d8047e0522069f06bd066d06da053405c504d9046a05450620078f075c07ad06bd05e50478047404aa04e704f004c30494048604bc044505ee058a060f077407cf074908d608500989093309260888069a04d702cf01d201f20202056a0790090b0b960b4d0b9f0ae8096b093a090b098c089407180666040b036d02ce022f0424062508bb09790a410a5009ef0783067605f004f3046b051206b5064307a607e90731086b088408700807084407520656058b0432045404e904e60514074e088809980a6f0b060c2f0ccf0bee0a8709be07e505400411039202c3029403eb0488063b08e309420b2a0c850c290c0f0b6209490715053403ee017a01e90102037404ec051307d10749089308d308210950092d09a208a60765062e053a04b403ab03f8037e043205f805cb06ab077008f808330906097508a307a7069e05b004f10383038203e7039f048a055d06e9062d072a07ff06d706ae066e06fa053205270416033e02e50135020a032c0455053406a0069e0632067905a104c40303037f0242025302ab022b03c2036704fa046e05ba05bf057305e8043a049a033603180331035c036a035003280311033303950306044c043b04be03f7022d029a0164018a01e4014c02a502da02f002f002cf028d022f02bd0153010e01f000f5000301fb00d900af009800b4000d018201ea011502e2015c01a600eeff65ff2dff52ffdaffbb00ce01e602be030f04b803c4026801feffd8fe22fee3fdfbfd44feb3fe4bff12000a011302ed025b03340376024a01ebff99fe8afdddfca0fcdbfc80fd72fe85ff7c0016012e01ba00d4ffb9feacfdeefca2fccafc4ffd0bfec8fe5dffbaffd7ffb8ff78ff2affdefe9afe5afe15fec5fd65fd05fdc2fcaefce3fc6bfd33fe1dff0900c90038013f01ce00eaffa9fe35fdd2fbc2fa31fa3cfad7fac1fbbbfc93fd22fe69fe83fe88fe81fe6bfe2cfebdfd26fd80fcfcfbbcfbbdfbebfb21fc30fc17fcfdfb0dfc72fc36fd28fef8fe53fffefe04fea8fc4dfb66fa44fae8fa27fcaafdf4feabffa4ffe8febafd79fc79fbf3faeafa2cfb89fbd3fbf3fb00fc21fc63fccdfc4efdbafdf4fdf3fdb5fd4efdcefc3bfca3fb0dfb77faf6f99bf965f968f9b4f946fa1bfb24fc31fd15fea8fecffe99fe1dfe70fdaffce2fb06fb35fa94f944f970f921fa30fb66fc80fd3cfe82fe56feccfd19fd69fcdbfb90fb89fba4fbc6fbcffbacfb7bfb6ffbadfb4ffc34fd09fe7afe47fe61fd0ffcb3faaaf93ff979f925fa0efb00fcd7fc98fd43fec3fe02ffd8fe24fefafc8ffb2afa29f9c4f8fef8c3f9d8faf2fbebfcabfd25fe71fe9dfea7fe94fe50fec1fdebfcdffbc5fae6f97cf99ef94afa45fb3afcf8fc65fd88fd95fdb5fde9fd1ffe1ffebafdf5fcf6fbfffa6bfa69faeffad7fbd0fc87fdd9fdbefd45fda8fc18fcacfb7cfb85fbb4fb01fc5afcaffc04fd50fd84fda2fd9dfd6afd1cfdc6fc7bfc5cfc73fca9fce6fc04fde8fca1fc4dfc18fc38fcb4fc70fd43feeafe2cff00ff75feaffdeefc63fc23fc33fc74fcbcfcf0fcf4fcc1fc76fc2bfcf1fbe1fbfefb41fcaefc37fdc9fd5dfed1fefdfed3fe4cfe7afd89fca2fbeffa98faa2fa05fbbafb9ffc7dfd2dfe82fe6efe0bfe8afd24fd0dfd3efd8bfdc6fdbbfd62fdebfc8ffc7afcc2fc41fdbefd0afe07febbfd51fdedfcb0fcb4fcf2fc56fdd0fd34fe61fe50fe00fe87fd16fdccfcb5fcd1fc05fd38fd66fd8dfdadfdcbfdd6fdc0fd8dfd43fdfefce4fcfcfc36fd82fdc7fdf3fd13fe35fe66fea5fed4fed5fe9bfe1bfe6bfdbafc2dfcdffbebfb4afce9fcb6fd8bfe42ffc5fffcffe1ff7effdffe1cfe54fd9dfc14fcd9fbeffb4bfcdffc88fd28feb2fe21ff72ffa2ff9aff47ffa4fec2fdd4fc24fcdffb15fcb6fc85fd4cfef1fe6dffc8ff0f0035002800d5ff35ff66fe94fde2fc6ffc4ffc7bfce9fc94fd6afe4eff1b00a600dc00be005900d1ff46ffbffe3ffed1fd7cfd57fd73fdc5fd35fea0fee8fe0eff2fff6fffe2ff7500ee001201bd00f2fff0fe0bfe7dfd5cfd9bfd09fe79fed9fe2aff77ffc6ff070022000700acff2cffb1fe5ffe53fe95fe0bff93ff0f005c00710057001f00e0ffadff87ff64ff3afffdfeb6fe82fe7afeb6fe38ffe7ff9a002b017a01820157011001c900950071004f002400e3ff8fff35ffebfec7fedafe26ffa4ff4900fe00b1014902ac02c3027e02d701e500d5ffe3fe4dfe3cfeb6fe97ff9d00820118024f023602ec018f012901b9003b00bcff5cff44ff92ff4e005c0181027d0313041f04a203b002740129000eff58fe24fe70fe28ff2700380138021403bc031e043004e703420353023e01370072ff13ff2bffaeff750057012a02c3020e031103da027f021d02c801880162015b017801ba011b028a02ee0223031703d60273021002d601d50100023b026302660245021102ec01f30130029e022903b00310043004fc037b03ca020e0272011501000129017901da014602bf023d03b6031404360406048e03ee025a020102f7013b02ae0227038503b1039f035303d9024202ae0148012c016901fc01c00286031c0463045f042204c50369031e03e302bb02a802a902c202f1022203440343031503c80277023f023a027102d5025903e5036204c8040c051805e1046704ae03d302050272013f017401f901a9025903df0333045e04680463045a0440041304d1037203020395023402f201de01f9014602c1025103e5036904c104de04be045e04d2033703a70241021a0223024b027b029d02b402dc022f03c2038e045e05f1050a067e056004f40291018f002b0062000e01f201cd027e0305046704b104e604eb04ac042d048103d60263023d025c029d02cc02cb02a102680251027f02eb02790300044c044a040a04a5033f03fb02e202f1021c034b036f03830382037b0377036e035d033a03f00285021802c801b90101028d023403c1030604ff03c80383035403490343032303d1024702a4011701c000b600ff0084012e02e80298032e049a04c304a5044c04c30324038b020002930149011d01130130016501ab01fd015102aa020b036803b903f5030304d8037603df022d028201f700af00c3002701c1016b02ef022d031c03c8025702f301ae019201a001c501fa013e028402c302f302fe02d902850202026701d500630030005c00df009f0178022f03950399034003af02180294012b01d9008e004d002b004000a100490105029802d5029f02060244019b003a0033007500dd0049019801c401d501d001bf01a801860158012301de008b003500e6ffaaff94ffb2ff0c0099004501fc019f0207031703c2020402f300c4ffb1fef6fdbafd00feb2fea3ff9c00740115027402920279022d02b80127018100d1ff29ff96fe2afef8fd14fe88fe49ff35002401e50148023d02d1011e014b0089fff4fe9afe76fe79fe92feb4fed8fe0dff5fffcdff4f00d10028013001dd0032004dff59fe86fdfbfccdfc02fd95fd6dfe63ff55002501b301e801b9011e011f00dafe81fd56fca1fb8afb1afc2ffd88fed7ffe0008001b0017901eb00160013fffefdfdfc3dfce2fbfcfb81fc54fd47fe25ffc2ff0300e9ff8dff11ffa0fe5afe3ffe3afe2efe05feb9fd5dfd19fd0cfd45fdb4fd38fea7fee5feebfec7fe8dfe4ffe19feeafdbafd88fd5afd33fd23fd32fd61fda9fdfefd4efe8cfeacfea4fe77fe2bfec3fd50fde2fc83fc44fc31fc54fcb3fc3efdd4fd57fea8feacfe68fef2fd67fde6fc86fc51fc4efc7cfcc8fc26fd83fdc4fddefdd2fda7fd79fd5dfd56fd64fd7dfd89fd87fd78fd57fd2efd08fdeafcdafcdffcf9fc24fd4cfd5afd52fd3bfd20fd19fd3bfd77fdb7fde0fdd2fd89fd18fd97fc2bfcf3fbf8fb39fca4fc19fd82fdccfde4fdd3fdb0fd8afd75fd75fd75fd60fd22fdb3fc2efcbcfb83fb9ffb0bfca4fc47fdcefd1bfe2ffe1cfeeefdb9fd8dfd6cfd58fd42fd13fdc9fc63fceffb96fb80fbb9fb3ffcebfc81fddcfdebfdb8fd6cfd2efd14fd29fd57fd83fda4fdb0fd98fd66fd23fdcdfc72fc25fcf2fbeefb1bfc6dfcdefc5bfdcbfd2afe64fe63fe2afec2fd3efdccfc91fc97fcd9fc32fd69fd67fd29fdc1fc63fc36fc49fc9afc0afd76fdd2fd17fe3afe4cfe54fe44fe1bfedafd76fd00fd8cfc2cfc05fc22fc6ffcd6fc33fd5efd56fd30fd09fd0efd50fdb8fd2ffe8efeadfe8cfe39fec4fd4dfde6fc8bfc44fc15fcf5fbeefb0bfc4dfcbdfc55fdfbfd99fe13ff46ff30ffdafe51feb8fd2bfdb3fc61fc39fc2ffc45fc79fcc3fc1cfd79fdc8fd0afe42fe77febafe09ff4aff63ff35ffaafed5fde3fc08fc79fb55fb91fb1dfcd3fc8bfd34febefe18ff40ff34fff3fe96fe2bfebcfd5bfd0efdd7fcc2fcd5fc0efd6afdd3fd24fe4ffe4afe19fedafdaffdadfde2fd3cfe99feddfee8feabfe3dfebcfd45fdfffcf6fc1ffd67fdb6fdf8fd32fe68fe9cfed2fef8fef4febffe59fedafd72fd44fd5bfdb6fd2efe8dfeb4fe9bfe4efef8fdbdfdb0fdd8fd1afe4efe61fe4afe15feebfdedfd29fe9dfe26ff95ffcbffbdff73ff14ffbffe81fe56fe2efef4fdaafd5ffd2cfd37fd90fd2bfef0feb8ff5300a2009b004800ccff48ffd0fe70fe25fedefd9efd71fd6bfda2fd1afebefe6dff00005c00790060002400d8ff84ff2dffd9fe8dfe4bfe18fefffd05fe2ffe7ffef1fe73ffedff4800710064002f00e2ff8bff3bfffffed6fec4fed4fe0cff69ffd8ff3f00870098006a000e009eff2fffdbfeb0feb2fee1fe3affadff29009800e3000001ec00b10066002000e2ffb0ff8aff6eff63ff74ffa4fff2ff5000a900f300220130012101f500ac005200f8ffadff86ff8affb9ff0a006800bf0008013a01500150013c011701ee00c700a50091008c009200a500c600ed00170136014501430132011a010c010d011a013701590172017b016d014a011d01f100d000cb00e5001a015f019f01cb01df01d501ba01a5019b019d01a601a901a401a001a301b201d501f601fd01e0019f0151011b0113014301a80120028e02e90225033e033b031303c4025d02e6017901370129014e01a10109027402dd0233036f038b0370031b03a0020e02850130011c014501a20113028202ea0242038903c803ef03f303d503890313038e020502920158016201b1014102e7027803da03f703d903a80378035b03580355033c031203de02b602b502d602070334033a031203d902a902a102dd024d03cc03340455041c04a6031b03ae029102c5023503b90312041d04e5037b030303ae0289028a02a702c502e1020a034d03b8035004f5048205d305c20546057704710364028701fa00d7002f01e901e302f703ea049205e205d2057305e4043a0492030903a4026702570267029002d7022d038f03fd0359048e04960468041104b203610335033c0361039603d403030419041604e6038f032b03cb028e029702e2025b03e203420460044004ec038d0358035e039c03fd03470455041d049e030103880255027902e5025f03b703db03c5039103710377039b03cb03e203d603b303850361035a0357033c030703b702680245025f02b10228039403d103d903b00370033f032a033303520368035a032303c2025002fc01db01f8015202c6022a036b037e037203640364037a03a003b4039d035803e7025b02d9017d0158017301bd0121028a02dd020c031e0316030003ed02dd02d102c802b20288024c02fb01a4015b012b01250150019c01f1013c026702700268025d0261027b029902a4028a024702ef019e016601540160016d0169015901470146016601a001e1011a023e0251025e0266026a025c022602ca015901e10075002900fdfff0ff0a004e00c0005201e40155028c0279022702b5013801bf0058000a00ddffdaff02005000b10006013d0154014b0130011201f300cd00a40080006b006e008800ab00c300c300ad0090007a00770087009b00a200900062001d00d6ff9fff84ff8fffc2ff10006500ac00d500d200a3005a000d00c8ff91ff6dff5eff5dff66ff7cff97ffa8ffa8ff99ff85ff80ff94ffc6ff0a00450057003700e9ff82ff24ffe9fedafef4fe28ff62ff98ffbfffd0ffcfffbcff95ff64ff33ff05ffe6fedafedcfef0fe13ff37ff59ff77ff89ff8bff7bff5aff32ff02ffc6fe82fe3bfef5fdc6fdc1fdebfd47fec2fe38ff92ffc2ffbbff83ff2cffc1fe51fee8fd90fd59fd4bfd60fd9bfdf3fd4ffea5feedfe17ff21ff11ffedfec3fe9dfe79fe5cfe3ffe15fee5fdb9fd97fd89fd93fda8fdc8fdf0fd1bfe4dfe83feabfeb7fe9dfe57fef6fd94fd41fd10fd05fd14fd38fd67fd95fdc0fdddfdddfdc0fd88fd3cfdf9fcd3fccdfceefc29fd65fd98fdc0fdd7fde4fdeefdedfddffdb5fd64fdf8fc7afcfefbabfb9ffbddfb65fc1cfdd3fd6afec4fed0fea1fe4afeddfd6ffd07fd9efc3cfcddfb84fb4cfb46fb71fbd8fb6cfc07fd8efde3fdeffdc3fd73fd0efdb2fc69fc27fceefbc1fb9efb97fbb4fbe7fb28fc5dfc67fc4dfc1ffcf3fbeefb21fc71fccafc0dfd1cfdfefcc7fc82fc4bfc29fc12fc0cfc18fc27fc39fc40fc25fcf2fbb8fb8afb8dfbcdfb2efc92fcd8fce0fcb7fc7cfc41fc1ffc17fc13fc0afcf2fbbcfb74fb1ffbbdfa6dfa4dfa69fad1fa7bfb38fcddfc42fd4afd0afda5fc32fcd3fb92fb5efb30fbfdfabdfa85fa69fa73fab8fa3cfbe4fb95fc2afd79fd7dfd3cfdc3fc41fcd3fb82fb58fb4bfb41fb36fb23fb09fb00fb15fb45fb9afb03fc63fca8fcc4fcaafc69fc16fcc3fb8cfb75fb6ffb6ffb65fb40fb0efbdcfabdfacdfa09fb57fbb1fb06fc44fc76fc9ffcb4fcb5fc95fc49fce5fb7bfb1cfbeafaeefa17fb64fbc5fb20fc70fca9fcc0fcc7fcc5fcbffccafcddfcdbfcb8fc6cfcfdfb95fb5afb5bfb9ffb0afc6bfcaafcb9fc9dfc76fc55fc43fc4bfc65fc7afc8bfc91fc82fc69fc4afc28fc12fc11fc1bfc32fc4ffc68fc83fc9bfcacfcbcfcc2fcb7fca7fc9dfc9cfcb5fce6fc20fd61fd9efdcbfdebfdf6fde0fda7fd4ffde4fc8efc6ffc94fcfbfc83fdfcfd45fe50fe25feebfdc4fdbefddcfd09fe26fe1efee6fd89fd23fdcffca3fcb3fcf8fc5afdc5fd1bfe47fe4ffe3efe25fe16fe1afe2afe40fe4dfe49fe39fe20fe08fefbfdfbfd03fe12fe2afe56fea3fe0aff78ffd9ff0a00fcffbfff6dff25ff00fffbfe02ff02ffecfec7feadfeb2fee8fe52ffd5ff5200af00d100a8004100b2ff17ff98fe4cfe3afe61feb3fe1eff96ff0c007200bc00da00cb009b0054000000aeff62ff2cff24ff51ffb3ff3600b30009012a011a01f700e700f800290166019001970178013b01f800c600ac00af00d100010133015b0175018d01b101ea013b028f02bf02b0025802bb01040169001500250090003101db016002a202a8028a026402480236021e02f501b4016601300127015601bb013a02b4021b0364038c039a038f036b033203e5028e0248021c0219025202bf024c03e7036b04b304b5046f04f80378030c03cd02d10204034c039a03cc03d103b803880354033f0350038003cb0314043b043d041404c703770336030b030603230353039303d4030b043904510455045704590467049004c204ea0406050605e304ae04710436041404100436048d04fb046405bb05e405dc05bd05980574055d0541050e05cf0488044604210416041e043a045f048e04d6042e058805dd050e060606c5054805a104fc0379033c036203da037d042705a705e605f305dd05bb05ab05a705a405a20591056a053c050c05ea04f4042905870505067906c406dc06b0064a06ca054005cb048d048604b6041d059205f5054006600652062606d6056805f2047d042204060421046204b804fd0422053a05470557057c059d05ab05af05970563052905e0048d04570448046d04cf044805b005f405ff05d705a6057d056c058105a205c005dc05e205cc05aa0573052a05e10497045a04400445046c04bd04160563059805980564051b05c604760440041204e103b4037e034f0345036103a7031e04a60422057f0597056005f1045a04bf034d03100312035503bb032d049d04ec0413051f050b05df04ac0468041a04d4039b0380039403c203f60321042a041304f303d703d303e903f403d9039203180388021902eb0114028d022603b3030504f9039a030f037602ff01cd01d6010b025302870297028902680258027402b102fd023c0340030603a9024702070201022302570287029e02a2029e0290027e0270025b02400224020102db01bd01a5019d01b101d101eb01f301d60196014a010401d800cf00d900e800f200ec00d300b0008600670063007a00a900d900e800cc009100470012000f00330069009b00b000a7009000780069006e0081009800a700a100890066003f0028002e0044005a005a003800fdffc0ff92ff86ff94ffa4ffa0ff84ff58ff2bff0afffbfefefe08ff0cff08fff3fec6fe8cfe51fe29fe25fe48fe7efeb0fec9febefe9dfe77fe5bfe4efe46fe3efe35fe2bfe2bfe42fe65fe88fea2fea8fe9afe82fe66fe50fe49fe48fe49fe47fe32fe09fedcfdaffd8efd8afd9cfdb8fdd7fdeafdebfdd6fda8fd65fd16fdbbfc6cfc41fc40fc6efcbffc0efd43fd53fd32fdeffca5fc60fc2ffc15fc02fcf3fbecfbe9fbfefb35fc86fce1fc2afd40fd22fddafc77fc20fcedfbd6fbd8fbe9fbf2fbf7fb03fc14fc39fc73fca9fcccfccdfc9afc47fcebfb94fb60fb57fb64fb81fb9dfb9ffb8ffb79fb5dfb4dfb52fb61fb76fb81fb6ffb49fb12fbccfa97fa7ffa77fa84faa1fabdfae1fa0afb24fb30fb26fbf8fabffa93fa74fa72fa89faa0fab7facbfad6fae3faf0faeffaf2faf6faedfae9fae8fad8fac4fab6faa7faa4faabfaabfaabfaa5fa96fa9afaabfaaafa9cfa7ffa46fa14fa02fa09fa27fa47fa45fa29fa01fad1f9b7f9bcf9c7f9d7f9e6f9e5f9e2f9e7f9eaf9fbf919fa35fa4ffa58fa3afa04fac8f996f991f9c1f90bfa5ffaa1fab5faaffa9efa86fa7ffa85fa7efa6dfa51fa1cfae7f9c6f9bcf9dcf922fa6bfaacfacefabbfa88fa4ffa18fafdf9fdf901fa07fa02fae6f9cef9c1f9b6f9c0f9e3f909fa35fa5efa64fa4efa27faf6f9dbf9e1f9f8f91cfa3dfa4afa52fa5bfa62fa79fa97faa6fab8facafac9fac0fab6faa0fa90fa8bfa8efaa8facafadbfae7faf2faf8fa0efb33fb4afb4efb30fbebfaa3fa76fa6bfa90facffa07fb32fb42fb2ffb19fb0bfbfcfafbfa02fb00fb01fb03fbfdfa00fb0cfb16fb2cfb47fb58fb6afb76fb70fb70fb7cfb88fb9efbaefba6fb96fb8dfb8ffbb3fbf5fb3afc71fc8bfc7efc5efc38fc13fc02fc08fc1afc37fc57fc71fc87fc8ffc8cfc92fc9dfca4fcacfcaafc91fc75fc61fc55fc5ffc79fc96fcb4fccbfcd6fcdffce0fcd7fccffccffcd7fceefc0efd2bfd3ffd45fd41fd42fd4cfd5efd7bfd98fda9fdb1fdacfd9bfd8dfd94fdb4fdf0fd38fe71fe86fe6bfe2efef7fde5fd01fe45fe8ffebffec3fea1fe73fe56fe55fe72fea2fecffeedfef7feeafeccfeabfe96fe95feadfed6fe03ff26ff38ff3eff44ff4aff4fff4cff3aff21ff0fff15ff3dff82ffd0ff1100340033001b00f8ffd5ffc2ffc5ffdafffcff22004300610081009f00bd00d900eb00e900d600bd00ac00a900b800d500f3000701110116011d012e014301580169017001710175017c0185019201940187017901700170018401a501c701eb010502130220022c0238024e02660271026c02520227020102f60115026702d10230036e037603510322030003f80210032e033f03430335032103210337036203a703e90310041c04ff03c00383035c0357037c03b203e003fe03050400040704130421043504370422040f04fd03f6030b04300459048f04b804cf04e104e404d904d604d104c104b504a50493049704af04db041e0558057f059d05a305960590057c054f052405fa04d804de0409054c05a305ee051a062d061806e405b10581055c055805640576059605b105c405e105f705050612061006030601060106040617061d060d06f705cf05a4059b05ab05d10511064d0678069c06a806a2069d068a066d065a063d061606fd05ee05ee05120647067d06b106c806bc06a6068b067b068a06a106b006b106880641060206d805d70512066906c00605071007e1069e06530618061006280646065d064f062006f505dd05e70520066c06ae06db06d706ac06760638060606f805fe050d062c06410646064c064a064506520660066e067f067b06600644061d06f105d905c805bc05c505d405e405ff05120617061b061306fe05ed05d305af05930573055205450541054a056e059605b405ce05d105b6058c05570524050905ff040705260541054e0556054c053505270519050a050505fb04ec04e604db04ce04cb04c004b704c004ca04ce04d804d204bb04a4048604630449042d0413040b040c0416042f043f04400440043a04310429041204ea03ba038303540342034303540375039403ad03c003bf03a80389035e0333031603ff02ef02e102cc02be02c802e002040330034b0348032f03fd02c0028802580237022c022f023c0249025002590264026c0273027602650245021b02eb01c101a2018001640151014401470161018401a701c001bf01a5017c014a011901f000cc00b200a20099009c00aa00c300e200000111010f01f300bd007c003d00100001000d0026003e004c004c0045003c003b004200450038001800deff96ff58ff32ff2eff4fff82ffafffcbffccffaeff7bff42ff11fff5feebfeebfeeffeebfed8fec0feaafea3feb0fec2fecdfecffec3feadfe98fe81fe62fe3bfe0bfedffdcafdd3fdf8fd2bfe57fe6efe6cfe4dfe25fe02fee2fdc9fdb8fda7fd94fd87fd7dfd7cfd8bfda2fdbdfdd6fddcfdcbfda8fd75fd3ffd14fdf3fcddfcd3fccffcd3fcdbfce0fce6fceefceefcf0fcf6fcebfccefca6fc71fc3dfc1cfc0afc0efc27fc44fc64fc8dfcacfcbcfcbcfc9efc6cfc3afc0efcf3fbeefbf1fbf3fbf4fbf1fbfbfb18fc39fc5dfc7afc78fc5bfc2dfce8fb9ffb65fb3ffb3ffb67fb96fbbffbd3fbc2fba6fb94fb85fb84fb90fb8cfb7bfb69fb4dfb34fb27fb17fb0afb08fb08fb19fb40fb66fb89fba0fb95fb7bfb5ffb39fb1afb0dfb00fbf7faf8faf6fafafa07fb0ffb20fb41fb5cfb70fb77fb5bfb2afbf2fab8fa98fa98faa1fab7fad5fae5faf2fa06fb16fb31fb4ffb58fb4efb2ffbeefaa8fa77fa5cfa6efaa7fae9fa29fb57fb5ffb55fb48fb34fb25fb17fbf9fad7fab1fa83fa66fa66fa71fa93facbfafffa2efb51fb5afb57fb4bfb26fbfbfacffa9ffa84fa89fa9ffacdfa08fb33fb56fb74fb80fb88fb8dfb81fb6ffb58fb34fb12fbfdfaf2fafffa26fb52fb7cfb98fb96fb83fb6dfb5afb57fb5bfb55fb4efb3cfb14fbf3fae5fae5fa06fb43fb80fbb6fbdbfbd7fbb7fb90fb67fb50fb4efb51fb5efb71fb82fba4fbd8fb08fc35fc5cfc6bfc6dfc67fc50fc2dfcfffbc6fb9cfb90fb9bfbc7fb09fc42fc71fc98fca5fc9efc84fc55fc22fcfbfbdffbd4fbd4fbcdfbcffbe0fbfefb36fc7ffcbbfce4fcf3fce3fcc5fca8fc8bfc79fc71fc6bfc72fc8afca7fccefc01fd33fd67fd92fda4fd9cfd75fd32fdf2fcc4fca5fca4fcbbfcd8fcfffc30fd5efd8bfdb0fdbcfdb3fd97fd67fd37fd14fd02fd0bfd27fd41fd5afd6dfd7afd96fdc5fdfefd3cfe6cfe78fe67fe3ffe02fec7fda2fd95fda5fdccfdfbfd2afe4cfe63fe7dfe9bfeb6fec9fec6fea6fe73fe36fefefde0fddafde8fd0afe35fe62fe96fec7feedfe0eff24ff26ff1cff02ffd7feacfe8cfe85fea1fed8fe19ff5bff92ffbaffd4ffe1ffe0ffd2ffb2ff85ff55ff28ff09ff02ff0fff2eff5aff8affb5ffd9fff2ff01000800ffffe3ffb6ff7aff42ff22ff24ff4aff8effdfff2f007200a300c000c400ae0087005900340029003700520073008f00a200b700d500f900210142015401550144011f01ed00b600830063005e007500a600de000c012b01390135012a0121011a0114010b01fd00ee00e600f00018015c01af01ff01340241022c020102d401bb01b701c301d901ed01f601fd01050215023a026a029602af02a40271022802dc01a2018c019501b101de010e023b0268028d02a302ad02a80295028202700257024202350233024a027a02b802fa0235035c037003720368035a0341031b03f302cc02ac02a202af02d00200032d034e036a0375036a035d034a0329030603e402c502b602c002e002160351038503ad03bf03c103c703c603bb03b0039c037b0361035203500363038303af03ea031c043a044b04440425040304dd03b0038803620344033e034b0361038303a303bd03e103060421042f042004f003b90388036803640373038a03b303e9032a047204a504b0049b046a0436041b040d040404fe03ee03dd03e50302042c045c04760472045d0434040004d703b4039903920392039803a903b803c703e40307042a044b04550445042704f603c003a3039a03a203c103eb0318044b0478049904b104b2049d047b0449041004dc03ac038d038c039803af03d303f5031204310446044e0447042404ec03ad036a03320317031303250352038d03cd03100443045f046c04630443041104cc037d0338030d030e033e037f03be03f1030b0418042c04390432040b04b8034903e602a3028d02a602d102010337036d03a103d703f803f203cc038a033803ee02b302880276028102b00202036103b303ea03f603de03b9038d035d032603df0290024d0221021d0246028702cf0212033a03420330030403cc0296025e022d020d02f601e901ed01fd011f0259029902d30200030803ed02c3029502700258023f021e02f801d401cd01f0012d026f02a002a8028f026c0246022002fa01c60185014a0123011c01340158017e019b01a901b201b701b1019f0185015f0138011301f200e000e700fd00230155018301ab01cb01da01d301af016f012701ec00c900c100c700c700c100be00cb00f0001a012b011801de008b0043001700fefff7fff9fffaff070024004500620075007b0079007200610042001600e9ffd2ffdcff030031004a004500320025002b004500550042000900baff74ff4cff41ff45ff49ff42ff3bff46ff5dff78ff90ff96ff85ff67ff3dff0affd6fea5fe84fe80fe9afecdfe10ff51ff86ffa9ffb5ffadff93ff6fff49ff24fffcfed1fea3fe74fe57fe60fe89fec5fefbfe10ff03ffe5fec3fea7fe8bfe59fe0ffebcfd75fd59fd6efda0fddafd0bfe2cfe48fe60fe6afe61fe48fe25fe08fef9fdeafddafdc9fdc3fddefd22fe6dfe9ffeaafe8efe69fe58fe5afe5cfe3ffef1fd8dfd41fd29fd46fd78fd91fd86fd66fd4afd4ffd6ffd84fd73fd3efdf9fcc5fcb8fcc6fcdafce3fce0fce5fc04fd39fd76fda4fdb4fdaefda2fd96fd8ffd8ffd8bfd7bfd60fd41fd2bfd26fd39fd67fd97fda5fd89fd4dfd07fde3fcecfc03fd0afde9fc9dfc4cfc21fc24fc4bfc78fc86fc7dfc76fc7afc8efcaafcb4fcacfca3fca3fcb9fcd9fce8fce5fce3fcebfc0afd33fd45fd38fd15fdf0fcecfc09fd21fd1dfdfefccffcb3fcb7fcc3fcbffc9cfc5bfc28fc1dfc2cfc40fc3bfc0efcdbfbc6fbd8fb0ffc4dfc6dfc6efc68fc6afc87fcb0fcc8fcc4fca6fc79fc61fc76fcaefcf7fc30fd43fd3bfd28fd18fd23fd3efd47fd2dfde9fc84fc2efc05fc07fc27fc44fc3bfc19fc00fc04fc2efc62fc72fc51fc0dfcc9fbaffbc1fbdffbf4fbf0fbe1fbfafb4cfcb6fc16fd4dfd4dfd35fd29fd33fd47fd41fd0ffdccfc9cfc94fcbcfcf8fc20fd2cfd24fd18fd1cfd26fd18fde9fc97fc36fcecfbbffba1fb96fb97fba1fbc8fb0efc59fc98fcbcfcbafca8fc99fc8efc8bfc85fc71fc5bfc52fc5efc8dfce0fc44fda5fdeefd0afefefddefdbefdaefda3fd80fd3cfde3fc93fc78fc9ffce6fc1efd21fdeefcb0fc97fcaefcddfcecfcb4fc4dfceefbc8fbf4fb52fca1fcc1fcbbfcb5fcdbfc37fd9dfdd9fdcefd8dfd53fd4cfd79fdbbfde4fddafdb8fda7fdc3fd0afe4ffe5ffe33fee0fd8afd5efd5cfd64fd62fd4afd1bfdf4fceafcf6fc0efd22fd25fd25fd27fd26fd27fd2afd27fd29fd39fd54fd7afda5fdcafdedfd15fe40fe70fe9dfeb5feb9feadfe95fe82fe7dfe81fe8dfe9afe9cfe91fe7efe67fe56fe4dfe44fe32fe10fee0fdb4fd98fd8efd94fd9cfd99fd98fda9fdd8fd1efe5efe77fe64fe39fe1afe2afe64fea0febefeb2fe97fea3fef4fe75fff1ff2c001300cbff92ff8fffb8ffd4ffb2ff4effd7fe8efe9afee5fe31ff47ff1dffe1fed0fefbfe40ff65ff3affc4fe47fe07fe1efe71fec4fee7fedbfec7fedcfe31ffacff1c0058005a003b0024002d004d00680064003e001000fdff18005900a000c800c10098006e005f006a0076005f001700b3ff62ff4eff7fffccff0000faffc8ff99ff9bffdbff36006c005a001900e7fff5ff4600ac00e800e100bc00b300ed005a01b901ce0194013c010e012f017c01ac0193013701d600bf0003016e01b2019b013201bf008c00ad00f80025010801b5006600560099000301540169014d0127012a016301b501f201fc01d601a901a201d20126026e027d0250020b02e801070253029702a0025f02f701b201ba0103024d0258021502b30173018101d0011c022102db01800158018a01f4014c025f022b02ed01ee013f02b4020603ff02b2026e026f02bc0224035a033b03ee02b302bc020803580367032c03ca0286029502df021e031f03d3026a0236025402a502ed02eb029a023d0218024402ae0207030f03d3028a027c02d0025a03c203cf037e031203e50218038403dd03de038703270308034703c40322041b04c3035c032d035503a303c60395031d03a8028a02cf023f038e0381032803d602cc0218039203e103d1037a031b03f90232039503de03ea03bb0384037f03b103fa0330042704ea03ae039603ab03d903ef03d503a20373036a039303c603d503b70376033e033c0364039303a8038b03550340036103a803f2030a04e303a7037d038103ba03f7030904ee03b8038c039703cb0300041a040604d503b703b703cb03df03d1039a035c033503340359037d0383037103550345035603790394039a03800351033303330350038403b103c103ba03a6039b03ac03ce03ee03fa03dd03a1036703430340035d03780379035f03380324033f037103970394035603f402a8028b02a102ce02dd02bd028d0270028702dd023f037d03830356031c0304030f0324032c030d03d402ac02a802ce020d033a033f032c031103060314031a03fb02b9025e020f02f30107022f024a023602fc01cf01d2010a025e02930282023a02e601ba01d50118024f0258022e02f601e701090243026b02650240022802340257026e024f02fe01b0019701c30109021c02d2014601c500a300f3006e01af017d01f20070005300a7002b017a015301d60067005900bb004801960176011001bb00ca003d01bf01f001ab011901a4009900f100590173011701820021003800b70040015c01e40017006cff45ffa1ff19003800d3ff22ffa0feb3fe53ff170082005500c6ff51ff54ffcbff5a008d0038009fff34ff48ffccff5f0099005f00f0ffb5ffe8ff6300bf00a7001b0070ff0cff1aff68ff92ff57ffcdfe50fe35fe83fef2fe20ffe2fe60fefefd08fe72fee8fe09ffb3fe25fec5fdd6fd4dfed9fe1cfffcfea8fe71fe90fefbfe69ff93ff65ff0affccfedafe1eff58ff51fff8fe81fe35fe3afe7cfeb3fe99fe27fe99fd40fd4ffdaefd0afe0ffeadfd1cfdbefcd5fc4cfdcdfdfcfdb8fd38fde2fcfbfc7bfd13fe64fe4bfef5fdb5fdcafd2bfe8ffeaefe74fe0dfec3fdc0fdf6fd32fe42fe1dfee6fdc2fdbbfdc0fdb2fd83fd45fd0efdedfcdffcd0fcadfc80fc5bfc4dfc5bfc7cfca1fccafcf0fc09fd14fd0dfdfbfcf4fc09fd32fd61fd7bfd6efd51fd42fd57fd99fde7fd12fe0bfee4fdb6fda2fda6fda3fd88fd4efd00fdbdfc93fc75fc5afc42fc32fc3efc62fc85fc92fc81fc5cfc45fc4bfc5ffc6cfc62fc42fc2cfc36fc60fc9bfccffceffc07fd26fd50fd85fdb5fdd2fddcfdd4fdbefda0fd7afd51fd2ffd17fdfffce3fcc1fca2fc99fca8fcbefcc7fcaefc76fc45fc3bfc5afc81fc7efc38fcd1fb85fb87fbe0fb58fca3fcabfc8efc8dfcdbfc60fdcdfde1fd94fd27fdfdfc38fda5fdf0fdd2fd5cfdeefce3fc50fdf6fd5efe37fe9dfdf4fca1fccafc2dfd59fd0ffd61fcaefb6cfbbdfb60fcebfc07fdb1fc49fc34fc91fc29fd8cfd6bfde2fc5ffc54fce4fcbafd49fe3afeaefd28fd31fde3fdd1fe59ff14ff2dfe4dfd0dfd89fd4dfeabfe41fe55fd92fc8afc45fd32fe8ffe0dfe04fd2efc21fccdfc98fdd6fd51fd76fc05fc69fc6cfd5ffea0fe14fe48fdf1fc67fd62fe2eff3dff97feccfd87fd0ffe0dffd0ffd7ff28ff51fef5fd4efe07ff81ff42ff5efe69fdfcfc56fd27fec7febffe24fe79fd50fdd4fd9dfe03ffa7feb9fdddfcb5fc5bfd55fef4fed6fe37fec4fd0dfe0dff3200c1006c008bffd8fed9fe7bff200029007cff99fe37feb0feb2ff7e008000c1ffddfe85fee9fe94ffd5ff4dff46fe76fd6bfd1cfef6fe53ff00ff63fe20fe8efe76ff36004c00b9ff01ffbffe2dfff6ff84007800f0ff71ff7aff1e00f5006d013c019600fcffd8ff3400ae00cf006d00c5ff48ff4bffbdff35004c00e3ff3effd0fee4fe5fffe0ff0100aaff22ffd7fe0cffa6ff40007c004c00f9ffedff570006018b018f011c0199007700de008701f301cc012d0187005000ab00440192014a019600efffc9ff3700d2000f01af00eaff48ff3effcbff8100d7008e00e7ff73ffa1ff64003e019a014101890010004d0035013602a60243025f01b200ce00a5019f0208038c028401b100a50057012e026b02c901af00d7ffd1ff8c006201a00112011f0081ffb3ff870052017901e2001200c0ff3f00420117022e029001d800b4005c0166021c030a03530295016601e1019b02f902af02f70165016001d8015c027202f9014401cf00d800340173013e01aa001c00f9ff5700ee0047012801c0007900a9004601f10143021a02ae016901940117029c02cd02950239021c026102e4024b034503d4024502ef01fa01410267023202b1012801ea000e015b01850162010101ae00ac00f3004a0167012901c0008400a60019019d01e501d801af01bc012702c80246035a030a03a0027502a8020a03410314039a0229020f025102a602b7026102d10166016001a401d601a00100014d00fdff4100e20060015901df006a007d0039013102c6029502ca0110010e01dd01f7029b035e038302cc01dc01c002d9035504d803bd02d601ca018702530364037a021401230042003901370260027e01350077ffcbffee00f90113022d01feff7aff1f008d01c702ff022b020e01a3005b01c002de03f7031003ed017d01180246031c04f303e502be014f01d201c5024703d2029e0176001600a600910100028901730086ff71ff39003901a6012b012b0078ffacffb800ef017f0220024701bb000801150230039f0329033c029e01d201b1028f03bb030803ed0124012a01dd0192029d02d301a300caffc4ff6b0022014901b400c7ff2fff5aff260000014c01df00130083ffa3ff6a005901e401d1015701f4001301bc018802fd02da024202a9017c01d2015f02b5028602e0012501c100de005101ab019101f80029008fff6dffaeff01000e00b6ff30ffdefe00ff91ff4300b200b3006c0028002c008900090163016a013101f800fa004101ae01080224020402d101b701c201d601c2016e01e90060000100dcffe5ffefffd7ffa0ff68ff4eff60ff87ff9fff90ff5bff1afff7fe07ff38ff6eff93ffa7ffc1fffcff5a00c6001f0150015b0158015f01740188017e014801f400a5007d008700b000cc00b80071001800d6ffc1ffc7ffbaff73fff9fe81fe46fe5ffeaefee9fed9fe8cfe46fe54fed5fe91ff1f003600deff73ff63ffd0ff7a00f400ea00760010002700ce00a0010302a901d0000c00ddff4d00de00ee003e0025ff50fe39fec7fe65ff73ffcffeeefd74fdbefd91fe40ff3aff88febffd88fd1efe1cffceffc8ff3affcafe02ffe4ffde003f01cf00faff7bffc5ffa5006a017501bc00d1ff6cffd1ff9b00090199007aff68fe15fe9cfe66ffa1ffe9fea5fdb1fcbbfcb6fddbfe4affb1fe95fdeefc58fd94fec4ff0b003cff13fe9ffd63fe01006e01b601cc0088fffdfeb1ff250136020502a40002ff43fed6fe21000201ab0042ffc5fd3cfdf1fd3bff0500a4ff57fe07fd92fc23fd22feaffe60fe85fddffc06fdf1fd0bffaaff90ff0dffb8feeefe94ff3d00880068001d00010030007d00a80093005a003100310044003b00f3ff7dff0affc2fea1fe87fe51fe00febefdacfdcafdf3fdf7fdc4fd77fd50fd7ffdf6fd74febbfeb5fe89fe84fed2fe66ff05005d004a00faffb8ffbfff1d009d00ef00e90094002800e8fff1ff27004e002d00bdff2fffbcfe88fe90fe9ffe80fe2afec1fd7dfd84fdcbfd1afe3bfe1efee2fdbefdd8fd2bfe8afec5fed5fee0fe18ff8eff22008f00a4006f0034003d00a3002a01690125017e00d4ff8effcdff3c006100fbff36ff91fe7afeedfe73ff78ffc1fea7fddcfce4fcacfd8cfecbfe39fe57fdf4fc8efde1fe110053008eff84fe35fe12ff9c00c301b10180002cffd2fed5ff8801a7025c02e6005effecfed6ff4301ed01220148ff9afd33fd32feacff5d00aeff1efed9fcc2fcd3fd21ffa2ff00ffcefd0efd64fd96fec2ff1f0093ffc2fe82fe31ff70007601aa0112014a00040074003b01bf019d01ed003300e8ff22009a00df00ae00220084ff13ffe3fedbfed3feb8fe8cfe59fe2bfe04fef3fd0dfe54feb0fef8fe08ffe9fed4fe02ff7bff0e0064004b00e4ff97ffc2ff6e004101c201a9011d0199008500e20055016801ee002f00a8ffa6ff0600570032008dffc3fe54fe77fef0fe4aff2fffa2fe04fec3fdfcfd7dfeebfe07ffe3fec8fef4fe6dff0000690086006d00560064009300ce00f9000d0112011901240126011401f300d100b200900062001a00c1ff6cff29ff00ffeefee4fed8fec9feb5fea3fe9efea7fec6fef7fe23ff33ff1affe4febffedbfe45ffe0ff6b00ae009f006f006300aa002901900198013d01be0076009500fc0051013b01af00fcff8dff99fff8ff470028008effc7fe3ffe37fe93fef3fefefea9fe3dfe19fe6efe15ffaaffd6ff8fff21fff3fe3dffe4ff9000ed00e300a1007a00a00006016f019d0179011f01c8009c009d00ac00a10068001200baff79ff5fff69ff85ffa1ffa2ff71ff12ffa5fe59fe59fea5fe0aff43ff23ffc3fe7dfea0fe3aff05008d008a001900a8ffacff48002101a7018101d3002a001000a3007f01ff01bd01e6001500d7ff4200e1000d0176005dff69fe25fe9dfe59ffb7ff69ffb0fe1bfe1dfebafe7cffdaffa2ff11ffa0febcfe65ff3000a60095002900ceffdcff5f0015019c01b6016c01fc00a9009700b600da00dc00a7004e00fdffd8ffebff1d003b001c00bdff47fffbfe01ff47ff8dff8dff31ffaffe5cfe73feebfe73ffb2ff8fff41ff25ff7aff2500c100f000a0002800fdff5d002101d101f5018001d200670085000201630143019e00ceff52ff70fff2ff61005d00d8ff22ffaffebdfe2effa0ffb7ff5cffd3fe81fea1fe20ffacfff2ffd6ff8eff75ffc0ff5b00f0002901ec0071001c002f00a30025015c012a01c10076008600e4003f014401da003c00c5ffb1fff5ff4a005d000d0084ff0effe6fe14ff61ff8aff6eff20ffd9fed0fe12ff7dffd2ffe3ffbdff97ffaaff1400b3003501590115019e004f006200c5002a014401fa008b0056008d000501570126017600acff4eff91ff2a008900470074ff9cfe5afedbfec0ff62005100aafffcfed4fe53ff10007000280073ffe7fe01ffc5ffb70047013501ba005d007800f70074017f010601620001001b008c00f000fa00ae0051002e005a009800a1005400cbff48ff01fff8fe0aff0ffffdfeedfe02ff44ffa1fff7ff2b00460059006b0072005e002a00edffcdfff0ff5400c80011011201da00a700a900e600330150010d017f00f0ffa6ffbeff100048002e00caff61ff47ffa0ff3800a6009100f1ff1dff95fea1fe2bffc8ff0d00d6ff64ff26ff6bff1d00d0001401c3002200b0ffc3ff52000001540119018b0022003d00db009601eb019301ba00dbff73ff9fff0d003f00e9ff2aff7cfe5dfef3fee5ff9900a3000d004affe3fe1affbbff49005600dcff46ff0dff6aff3300f500420106018400220024007900cd00dc0098002e00ebffffff5700b400e600df00b80097008d0083005300f2ff7dff1dfff6fe08ff30ff4eff5fff70ff9bffe1ff210033000d00c0ff78ff5cff72ff9cffbcffcbffdfff15007200de0030015201500148014d0153012c01bc00160079ff2fff55ffc1ff27004b002600ebffd8fffaff2d003700efff6affeefebcfee4fe43ff99ffbcffb0ff9effb1fff7ff530092008e005000ffffc7ffbfffdfff0800270043006900af001401710196016b01fe007e002100fdfffdfff3ffbdff5eff09ff02ff5efff0ff67007d001f0089ff1aff08ff46ff91ff9aff46ffd2fe98fed6fe85ff5500e6000a01dc00a0009500c60002010a01c5005000e8ffc2ffeaff43009a00cf00d700bd008e0053001200d6ffabff96ff8fff80ff5aff2dff18ff32ff7affccfff8ffe6ffb0ff88ff92ffc0ffdbffb3ff4effebfee2fe61ff3b00fb0041010901a5008500e0007b01d401810192008dff19ff77ff5200fa00e3000d0017ffc3fe5fff83005d013e012400c3fefffd43fe38ff080004002cff34feeafda5feffff170145019600b8ff6fff01000001a2016a01820096ff51ffdbffba003a01fc003e00a1ffacff600033017e010301100048ff27ffa7ff49007700f6ff0fff5dfe5afefffed8ff520020006dffbefe92fe0dffddff7a00880015008aff5fffc5ff860026014501e00056001c006900070178015801aa00d9ff6effa8ff4d00d900dc00480089ff29ff64fff9ff5f002f0074ffa2fe44fe97fe5bfffeff0a0087ffecfec5fe4cff420016014801c700faff6eff7aff0700a300e0009f001e00d0ff000097003601790136019d000f00dcff090054006f003a00d0ff76ff66ffa0fff0ff1400ecff8eff35ff0bff17ff3dff4cff32ff09ff01ff3bffb0ff3900a200ca00b6008f0082009800bf00d100ac005200efffbbffddff4b00ca0019011701d20086006a007e0092006a00edff46ffc4fea6feeefe58ff92ff84ff53ff48ff93ff16007c007e0018008eff40ff58ffb3ff08001800eeffd1ff03008500130158012c01b2003d00170045008a00a700860044001c002f006f00ac00b80087003800ebffabff75ff40ff07ffd5febafec3fef1fe3cff9cff0d007600b600b9007e002800e7ffd2ffe2fff5ffecffc8ffb2ffd5ff4000cf0041016b014e011401ed00e400d6009c00270095ff26ff10ff4effb6ff090020000400ddffceffdffffcff0000d9ff8cff3bff0aff0eff48ffa2fff8ff350054005e006a008900ab00b50090003b00dfffb9ffe3ff4b00ba00ed00d0008f006e009900fa0040011f018300a9fffffed0fe15ff83ffb9ff93ff3fff16ff5bff0400b000f500a900fbff53ff19ff5cffd5ff23000a00a6ff54ff6afffbffc700620180012f01ba007b009200d400f000ad001e0099ff6effb2ff2f0089007d001a00a6ff73ffa0fffaff2f001100aeff47ff29ff67ffd1ff25002e00f1ffadff9dffd2ff2800660063002400d5ffb1ffd9ff38009e00da00da00b70096009200b000d400cc008d002e00d1ff9effa5ffc7ffdfffd8ffb8ffa3ffb5ffe6ff19002b000c00d1ffa1ff9bffb5ffcdffc9ffacff8dff90ffc9ff1d005f0074006000420041006600a300d300d400a7006a00370024003600570069005e002c00e5ffa6ff8aff9bffd0ff09001f000500d0ffa9ffaeffe2ff210034000300a7ff5dff59ffa2ff0a004b004000fbffb9ffbcff12008c00e600ed00a6004a001700290069009e009c0061001400e8fff3ff210048003a00eeff90ff5cff6dffbaff10002e000000a9ff5fff61ffbbff33007e006a00feff7fff44ff78fffcff770099005700efffc2ff05009e0036016c0113016800daffb5fffeff68008b003d00a6ff24ff11ff79ff11007b007c001f00b2ff7fffa0fff0ff2a001b00cbff72ff4bff6effbdff01001300f8ffd7ffddff0e0054008f009e0085006600590067008100910090007f006200410021000200e4ffcfffc4ffbeffb6ffabffa3ffb0ffd7ff06001400efffabff6eff5fff89ffc7ffe3ffc1ff74ff3bff5affd7ff6f00d300d7008d0043003f008400da00f600ad002600bbffb2ff05007200a20074000f00c3ffc4ff02003c003200d7ff62ff22ff3aff8effdaffe2ffa7ff67ff62ffa8ff0a003f001c00b7ff56ff40ff81ffeaff390049002d001e0045009f00ff002f011701d00082004f0039002a001100e8ffbaffa2ffabffc8ffecff07000c00ffffe7ffc6ff9fff78ff56ff38ff28ff2bff40ff5eff80ff9fffb9ffdbff0d004a008500a1008d0058002200110038007b00ac00ae0080004500300053009000b2008a001d00a7ff6bff85ffd4ff11000600b5ff53ff2dff63ffcaff16001000b3ff38ffe9feedfe36ff87ffaaff96ff72ff78ffc6ff4600c30009010101c300820069008500af00b4007f002200d4ffc9ffffff510088007d003c00f3ffd2ffeaff14001200d0ff65ff02ffdbfefbfe3aff67ff67ff49ff3aff55ff97ffe2ff100015000a0009001c003900450038002a00340060009c00c000ac006c00390041008000c500d3008900050099ff81ffbcff11003100f8ff87ff2dff26ff6fffcbfff0ffb9ff45ffdefec2fef8fe58ffa9ffcaffc4ffb6ffc1fff4ff43009500d000e400ca00860037000e001e0057008e008d004800f2ffd9ff2200a8000701f2006300aaff3eff5affc9ff1600e2ff35ff86fe57fecdfe9cff34003000abff1eff03ff80ff3c00ab007b00d4ff38ff23ffafff82001301120199001200ebff4100cf00270107017e00e6ff9dffbeff2000750080004100e9ffadffa9ffc9ffe1ffcbff86ff2ffff3fef0fe21ff5dff7fff88ff8effa6ffdeff260059005a002f00fffff2ff09002f0046003800120005002d008100db000601e60094004100190024003a003100ffffb7ff7eff72ff8fffbaffd4ffcfffb3ff98ff8cff8eff8dff80ff6fff6aff7bff9affbdffdefffaff17003f0067007c007a0067004c003a002e00220022003000450062007e0086007d006a005900540052003c000700b9ff6eff45ff4bff6fff92ffa4ffa4ff9dffa4ffc3ffe8fffcfffdffebffd4ffc8ffc7ffc8ffd0ffe3ff0a003e00690079006f005900570077009a009e007a003500f8ffefff1a0050006a0055001900e2ffd5ffecfffbffe5ffb0ff78ff5cff6dff96ffb6ffb9ffb0ffbaffefff380066005d002400e3ffc3ffd7ff08002c002100f6ffdefffeff4f00ab00de00ce009600650059006800720054000c00baff89ff8dffb4ffdcffecffe1ffd5ffe8ff1300330032000700c2ff8fff8affaaffd1ffe1ffd2ffbaffbeffefff3f008b00b000a10074004a003a00430055005900440022000900090023004a0068006b00550032001000fafff0ffe1ffc5ffa3ff88ff85ffa4ffd3fff8ff0a000e001100220043005b004d001a00ddffbdffd1ff0a003e004b003100110017005400ac00e800e000990041000b000a002e0043002100d8ff9bff98ffd5ff2700550048000e00d6ffcefff7ff25002900f5ffa8ff7bff94ffe1ff30005500410019000e0034007a00b300b3007b003100ffff010032006a00820070004500220021003d005b0063004a001500dbffb2ffaaffc2ffe2fff6fff5ffe6ffddffecff170046005d0050002b000600f3fff6ff00000200fdfff9ff080036006b008b008e007e00760085009f00a60083003d00f6ffdafff2ff220042003300ffffd0ffd0ff0a0050006a004100eeffa8ffa0ffd2ff0c001d00f2ffb0ff99ffcaff2a0083009a0069002100030029007700af00a4005c000700e6ff11006600aa00b00077002600f6ff020038006a0069002e00dbff9eff95ffc1ff0800390039001700edffd5ffe5ff120037003c001c00e6ffbaffbaffe8ff29005b0064004c003100310054008700ab00aa007e0047002a0031004c00600053002800fefff2ff0b00390053003f000b00d7ffc1ffd8ff080025001700e8ffbaffb1ffd4ff0c003b0043002500ffffedfffeff2a005600630051003300240033005a008100900080005b0037002200260037003d002d001200fdfff6ff02001a002e002c001f0013000800fffff8ffebffdbffd1ffcfffd8ffe9fff4fff8fffbff03001600330048004d00490041003b003d0046004a00450038002e0030003d00490049003f00320026002400250021001300faffe2ffddffecfffeff0700fdffe4ffcfffd1ffe6ff040019001400f6ffd2ffc0ffd2fffdff2c004900440023000300feff1c004e0072006b003b000100deffe7ff150049005e0047001a00f4fff0ff15004400550039000300d0ffb8ffc6ffe7fffaffeeffcdffb0ffaeffcbfff4ff14001c000b00f3ffebfff2ff00000c000f000c000700020006001500250035004000400033001d000900050010001d001d000500dfffcdffd9ffffff300048002d00f2ffc3ffbeffdfff0a001800f2ffa8ff6fff6fffaaff0300430042001000ddffcaffe6ff1c0041003a000300bcff95ffa0ffccff0600300039002c001c00160024003b00460041002500ecffafff89ff85ffa6ffd8fffbfffeffe8ffceffcdfff2ff220032001600dbff9bff7cff93ffc4ffe4ffdeffbbff9fffb0ffeaff2c0050003f00feffbbffa8ffccffffff17000100c8ff9bffa5ffe5ff340062004e000800c4ffabffc6fff8ff0f00f3ffb4ff78ff68ff93ffd8ff0e001800f5ffc9ffb5ffbfffd7ffe5ffd3ffabff8aff82ff96ffbaffd6ffdfffe1ffe9fffdff1b002e002000f5ffc6ffaeffb6ffd0ffe5ffe1ffc5ffabffb2ffdeff140035002a00f6ffbcffa4ffb6ffd5ffe0ffc5ff93ff6cff72ffa2ffdbfff8ffebffc4ffa8ffb1ffd2ffe5ffd4ffa4ff74ff6aff97ffdaff04000000d9ffb4ffb9ffefff2e0049002900d8ff8aff74ff9cffe4ff19001000d6ff9aff88ffb2ff01003e003900efff8dff4fff53ff8affccffe7ffc2ff7cff50ff61ffa9ff000028000400b7ff79ff74ffabfff1ff0700dcff92ff63ff79ffccff220041001200beff89ff98ffe0ff2a0039000000acff75ff7bffb9fffcff1100f2ffb7ff87ff7aff8fffb5ffd1ffceffb4ff96ff80ff7dff90ffacffc7ffd9ffd2ffb0ff8dff84ff9effcdfff9ff0100deffaaff92ffa8ffe0ff17002100f5ffb9ff96ffa5ffdbff06000300d7ffa2ff8bffa6ffd6fff2ffe7ffbbff8fff86ffa5ffcdffd9ffc0ff97ff7cff85ffb1ffdcffe3ffc5ff9eff8bff9affbfffdeffe3ffccffb0ffaaffbbffd6ffecffefffe4ffdeffe3ffebfff2fff0ffdeffc9ffc3ffcaffd0ffd0ffc6ffb6ffacffb0ffbcffcdffdaffd4ffbcffa4ff97ff9dffb3ffccffd7ffcdffb6ffa1ffa0ffbaffe1fffeff0000e5ffbeffa7ffafffd4fffbff0700f7ffd8ffbfffc3ffe2ff03000f000400e7ffcaffbeffc7ffd7ffe2ffdfffd1ffc3ffc0ffcbffd9ffe0ffdaffc9ffbbffb7ffb8ffbbffc1ffc4ffc2ffc2ffc8ffd6ffe5ffeffff4ffefffe3ffe0ffecfff7fffcfff8ffe8ffdaffd7ffddffefff03000800fffff0ffdeffd1ffd2ffddffe6ffe9ffe5ffdeffd7ffd3ffd5ffdfffeffffafffbfff2ffdfffcbffc5ffceffdfffeefff2ffedffe3ffddffe6fffeff110016000e00faffe7ffe1ffe2ffe8fff3fffafffbfffeff03000400000002000c00170019000e00f6ffd8ffc8ffcfffeaff070012000500efffe3fff2ff14002f0031001b00f6ffdfffecff0900190017000400eefff4ff1600380042002b00ffffe1ffebff100030002a00ffffccffbbffdfff2400590057002500ecffdafffcff38005f0051001400d9ffcaffecff2500490041001e00030006002c0058005f003d001100f8ff03002800410037001300eeffebff12004500630056002400f7fff2ff10003b0054003f000d00e6ffe0ffffff31005300550042002a0021002f004400510051004400350031003100300034003a003e0044004d004c004000310026002000260032003500290019000e000c0019003200470050004c00400032002d0032003e0049004900400032002b00330048005c00680068005e0059005f00660067005c00450032003200410055005e004e0030001f0029004a0070007a005d002900fdfff8ff230059006e0054002400000007003e008300a800990066002f00220049008300a7009d006a0038002a0046007d00a700a100780053004600560075007f006700400020001b003b0061006b0054002f001a002c005a008000840061002c000f00230055008200890067003f0032004c008300b300b900990071005c0064007f00970098007d0061005b0069007a00850078005f005300550060006d0066004600290021002f004e0069006d005a003c002e003e00610085009600860060004300410060009000b100b00092006b00570067008f00b200b4009400660049004d006a0087008d00760052003e0048005f006b00600043002c002e0044005d0061004b0031002a0044007200930091006e0046003c005d008c00aa00a2007b00560056007900a600bc00aa007c005800590074008d008c006b0042003100450069007c0069003b001700190040006e007c0058001c00f5fffeff36007c009e0086004c00200024005a009a00ba00a4006800330029004f008a00af00a500750042002f0044006e0089007e0055002900110016003100430039001c000500010012002d003c002d000c00f6fff9ff16003e004d0037000f00f4fffcff2c0061007b006c003c0011000c002d005c007d0075004a001900010011003c005d005e003c000900edfff9ff170030002d000a00e5ffd6ffdffffbff150016000200ebffe3fff4ff130024001b000000e7ffe7ff0100240038002e001000f5fff3ff0c002c003a0030001500f5ffe6fff0ff08001b001a000800f3ffe5ffe7fff5ff0700150018000b00f7ffebffebfff7ff0e002700300026001400050009001f0039004b004d003e002a002100280038004c00570051004000300025001d001f002b0032002c00200011000100fbff060019002700230011000000f9ff01001800290028001d000f000f002500410051005400430034003f0058006c0071005e003e0031003c0056007000730057002f0016001c003a005300550037000500deffd9ffedff080013000200e3ffc8ffbcffc8ffe0fff3fff7ffebffd6ffc9ffc7ffd2ffe8fffbff01000000fdfff5fff2fffcff0d001d0026002900230016000c000e0016001e0029002e0028001e0016000e000d001900220021001a000c00fbfff7fffbfffdfffdfff9ffeeffe5ffe2ffdfffdaffcfffc3ffbdffbcffbdffbaffacff94ff7bff72ff7fff92ff96ff87ff69ff4cff43ff53ff6dff7cff73ff59ff42ff3fff54ff75ff8dff92ff88ff7dff80ff95ffb0ffc4ffcdffd0ffd5ffe0fff3ff0600100015001f0029003600430044003e00380035003d004800430037002b001b001000110012000d000100eeffdbffccffc0ffbcffbdffb8ffb2ffaaffa0ff97ff90ff8aff8aff91ff99ff9dff95ff83ff75ff74ff7dff8eff9eff9eff8dff76ff69ff6bff76ff7fff7eff6eff4eff2eff1fff21ff2cff2eff1dff00ffe2fec9fec0fec5fec2feb4fea3fe8dfe7afe76fe77fe75fe74fe72fe72fe79fe82fe8dfe93fe8cfe88fe92fea5febdfed4fedafed6fed5fed9feeafe07ff21ff2fff2dff1eff15ff19ff27ff3cff4aff47ff3fff34ff28ff29ff32ff34ff32ff2aff19ff06fff9fef2feeefeebfee5fedcfecffec5febffeb9feb5feb4feb1feaefeaefea9fe9efe95fe8ffe90fe9ffeb7fec4fec1feb6feaffeb8fed4fefafe18ff21ff19ff15ff1fff3fff70ff9affabffb1ffbaffcbffefff2000440054005d00650079009800b700c800c700c200cb00df00f200fe00f700df00cb00c400ca00d100c900ad008a00690054004d00470039001b00f3ffcfffb8ffaaffa0ff93ff80ff6cff57ff42ff36ff33ff31ff31ff32ff34ff30ff29ff24ff21ff26ff35ff43ff4aff4cff47ff40ff47ff57ff65ff6bff66ff59ff4aff3aff33ff36ff32ff27ff1aff00ffe1fed0fec4feb7feaafe92fe71fe50fe2ffe19fe08feedfdcffdb0fd8dfd75fd66fd4dfd34fd1afdf5fcd9fccafcb8fca5fc8cfc64fc3afc1ffc14fc18fc17fc00fcdbfbb3fb91fb8cfb9efbadfbacfb96fb71fb54fb50fb66fb8afba4fbabfba7fba3fbaffbd7fb0afc39fc5efc75fc8afcb0fce5fc22fd64fd99fdbefde8fd1cfe5cfeaafef1fe23ff4bff73ffa1ffdfff23005b0081009500a700cb00fb002c0154016701670163016b018201a101b701b701a30188017f018a019901a10197017e0168015b015c0168016b015f01540149014001480156015d016401690172018901a301ba01d501eb0100022602520277029d02c102de0207033a036a03a103d80304042d0456048104b704eb0416053e055a0568058005a005bb05d705ec05ef05ed05ee05f205fd050206f605e505cb05b005a905a705960584056f0555054a054b054f055c055e0555055e0576059605ca05fb0518063a0663069806ee0649079707e7072b086508ba081d097b09d909230a570a900acc0a080b500b8a0ba80bc00bc80bc60bd30bdb0bce0bb70b8b0b4d0b110bd10a8d0a4c0afe09a5094c09ed0893084208ea0794074007e4068f064406fb05b80576053205f604c40498047e046b044a042e041004ed03de03d703c803b80391035a0332030503cd02a20264020902b0014d01dd007900050077ffe9fe4afea0fd07fd61fca5fbeefa31fa6df9bff812f85ef7b4f601f648f5adf421f498f31ef3a5f228f2bff169f129f1fff0d5f0aef095f07df074f089f0a2f0bff0e0f0f0f00bf13af163f199f1d2f1eaf106f22cf235f250f27df27ff27af275f242f220f217f2e4f1b6f18cf12bf1d3f097f03cf0f5efc0ef54efeeeea2ee35eee2edb8ed6bed1eede7ec98ec5fec51ec3bec32ec3dec2fec2bec4bec6feca6ecf6ec34ed6aedb4edfced4eeebfee30ef94eff9ef54f0aff01af18af1fef172f2cbf21cf377f3bff319f479f4b7f4f5f42ef554f581f5c2f5e8f509f63af646f64df67cf698f6aff6d9f6daf6d3f6f2f6fcf60ef73af735f724f72df713f707f71ff70af7e7f6d1f68af647f621f6d6f584f52ff5a4f417f496f3f7f258f2aff1d9f000f022ef33ee52ed66ec65eb68ea5ae956e878e794e6c2e50be53fe494e321e3abe26ce26ae25ae280e2e8e24ce305e413e51de67ae726e9c2eab3ecfdee3df1cff3acf66ef974fcbaffdd024106e0094f0de610a1141e18bb1b711fdd225226c729e22cf52ff932a0353538a43aa63c8c3e46409f41e642fb43a8443c45954593458f455745cd4440447643674274415140f43ec23d643cd53a8339183894365e350f34ab329e318530622fa92eea2d1f2db92c472cce2bbc2ba32b7d2bb32bdd2bf72b5e2cb22cf32c792dea2d3b2ebc2e242f6a2fc82f013014302f301830d62f892f022f542e972d962c692b252a9f28f9263f2543232e21011f8f1c0f1a8117b414df11050ff20be708e505af028fff95fc7ef984f6c4f3faf056eefbebafe996e7d4e52ae4b0e292e197e0cbdf5fdf27df18df66dff4dface0b7e105e374e428e623e82fea5fecc6ee34f1abf33af6b8f826fb9efdf8ff2a025a0463062d08e709760bb50cdb0dd50e6c0fd90f2210fe0fa30f2b0f510e420d230ca90aff085b07740573038e0177ff51fd5afb46f934f75ef578f39df102f061eed9ec95eb4dea2be93fe859e79ae614e6a1e54ee535e51be516e53ee560e599e5f3e52ee666e6a7e6c0e6d3e6efe6e3e6c9e6a9e65ee60ce6bce552e5ebe483e4fbe375e3fae270e2ede171e1dde04ce0c7df38dfb9de5adef3dd99dd69dd44dd43dd7fddcadd34decdde5fdf08e0e6e0b0e17ee26be32ee4f1e4d6e58ee64ee736e8e7e8a3e991ea46eb0fec06edaeed5cee29ef99ef16f0b0f0daf011f166f142f134f157f107f1d5f0ddf075f028f00ff07eeffbeea5eed2edf8ec39ecf1ea8ce938e866e66fe484e221e087ddf4da07d8ecd4e1d19ece27cbacc710c455c0a9bc06b950b59bb106ae74aafea6eba314a16a9e439c7d9a01994a983c989398c499b49bfd9d22a128a587a9a5ae93b4afba5dc1dcc884d0a7d893e18ceac1f39cfd6e075311ad1bb925702f3b396a42fa4a6353025bbb610068586db771907582787e7add7b597ceb7bdc7a0a79747633733c6faa6a7a65c05fb55934535b4c7e45603e35377730d1296c23bf1d5d186d13670fd20bd408d8064b0545042d0477043f05e106e508600b8c0efc11cb151b1a8b1e3c232728f52cc7316c36ab3ab23e2c42fb445f47e3487d499649a948c04664440541a83ce7374132ba2bfa247f1d3915c90cb803f5f951f0ade6efdcb4d3cccaebc18db9adb1f8a9cea25b9c4296c790488c63882f852283c881fb80538171820c84cd86608a4c8e44931699339f52a654ae7db662bf03c9a1d2bcdc6ae7d0f138fcd006d110771a1724072d5c35733dbd44474b8a512157fc5b7e604b6436679d694d6b1b6c5c6ce86b856a7768c66559626f5e2b5a805585505d4b1c46d940bf3be7363332b62d9829ab250322e51e101c7b196e179e1510143013b8129d123f134b14a815b2171d1ad21c1a208623eb26782acf2de930f6338e36b338823aa03b373c763c073c283bf239f9378f35d5325b2f7f2b5e277222161d73171011550a81031afc8ef439edb0e556de94d709d1ffcaedc575c1b9bd1abb2eb9eab7bdb74db869b97abb3abe5bc156c519ca52cf63d544dc7de356ebebf3c4fc0606bc0f4b19a422e02b8f34b13c6d44524b41516c56995ac65d49600a62e162f9625662dd60be5e1a5cb3587e54a74f064a9c43ca3c7a35862d4c25d51c1614a10b9b03cffba4f42dee24e8f0e2b9de25db66d882d611d53dd424d485d47cd515d714d993dba8de3de261e606eb17f08df538fb16011d07f60c9812f317941c8d20f7235f26ed27d02893287927e2255a231b208e1c39184a133a0e7d081c0289fb47f45cec50e4bfdbacd2c3c9f0c020b8b7afa7a7f59f0499d192588dd8885785ce824981b380f6800182cf836686a2897b8d059210979a9ce0a2aea9f9b00cb98cc141ca8ad307dd49e6b2efddf830011a09561043167a1be91fdf220c259226c1265f26aa25d1238721121f7e1b791760132d0e7808ad02c5fb67f426ed18e5eddc45d53ccd7bc5a8beebb7e2b11aada8a802a593a272a0009f859e1c9e169ea79e079f9b9fa6a08da1a3a20fa453a5d0a6a7a875aa78ac94ae61b009b26ab347b4ccb4c3b4feb39cb280b0d5add8aa68a7c1a30da0209c77984d95629225909f8e4f8dbb8c0f8dbd8d358f8091e293dc96b39ada9ee8a318aaadb033b802c17fca5ad5cae167ee13fbf707fe13421f2e2aec33a33cde440f4c95520f59e15e25643b69916d637124755178f47a317d7b7ef87eed7e117e887c4a7a0a7704734e6e0569a063f55dfd572252324c69465a419c3c30386e34b5302a2d592aae27442572238121af1f8b1e981d271d931d2c1e2e1fee20ea226d259128ae2be42e2a320635c5374e3a323cb73da83ec53e8a3ece3d673cc53aa338ea351b33ea2f382c6c2817240f1fca19f413660d960642ff3ef715efcce643def6d5f6cd05c68cbec7b770b1c4ab01a7b3a2e49eef9b6b99579726965d95d3941f95eb9517975799629ce19f6fa4d5a9b0af90b642be2ec6a5ce7fd721e0d0e89af1f9f913020e0a6f115f18461fce25fa2b2e320238473d72423b47584b2f4f6f52b1545e5655574a57b35680555f53bf50b44d1e4a6946af42c63ee63a1e375b33bb2f482ced2890252922c61e4c1bcc177d143511040e3c0bae087906fd04e90341035703c3037d04d2054307b7086d0af00b480dbe0ef10fec10e2117d12f3128513f3136214e014221557159215a015a2156c15ab148a13ff11f20fa70d0a0be7077504cd000cfd8ef95ff658f383f0e3ed77eb69e9d0e775e620e5d1e378e228e134e090df05dfbddea3deb1de68dfd0e0a1e205e5c4e79ceaf5edd2f1dbf523fa5bfe2502ce056f09e20c45106f1321169418ff1a791d1520b92231255a274d29272bcd2c2e2e292f612fed2e182ecd2c352b752932278824db21141f651c041a8e17f0146212c40f360de70a8608f3054603690088fddcfa44f8aef531f3c8f097eeddec9aeba9ea08eaa7e972e981e9d7e942eaa8eaf6ea14eb25eb3beb48eb57eb56eb40eb51eb85ebd0eb51eccbec1fed84edcdedf3ed1feef5ed60eda1ec84eb2ceae6e859e791e5d4e3e0e1f6df66dedbdc6adb2bdacfd893d79dd6a1d5c5d4fdd3fad20ed24fd19bd03fd021d009d04dd0e5d0bbd124d3ecd4d4d60cd964dbc2dd6be02be3d2e58de829eb88edf8ef62f296f4c6f6dcf8a1fa5cfc1afe85ffcd000002b60228038b036603ee025a021d0182ffeafdcafb73f943f795f4c5f148ef7aecc0e976e7d6e441e217e0a0dd4edb71d93cd71dd563d363d19dcf50cecccc76cb7aca47c94ec8aec7e4c633c69dc5c4c4f7c33fc35ec27cc179c038bfe0bd65bcdcba56b9a5b7e6b51eb431b277b0f1ae63ad19acfaaacaa903a9aba877a8c2a877a93eaa92ab91adedaf02b3ceb6d8ba6ebfbec462ca9ed096d7aede07e6f1edf0f535fe22070b10dc18fa21c92a4f33123c6344104c8953335a0e60b0659f6ad06ea4729375b07766795a7aa67a747a507970770075d171436e4e6ab765e260aa5b1256b450404bae458240383bec355c31fe2cf128ca25c2220320331e941c611b221bf61a0d1be71bd81c2e1e4d20842208250d280e2b532ee4314835b738ff3bc73e6741a0434045a74673477c473247384687448e42e13f7a3ccb386934572f0b2a2824a61df916d60f1b083c0020f88cefebe658de8dd5efccc9c4b9bc09b536aec7a7e6a1219ddd9819957b926590bd8e448e628ee58e9890f792c895de99c49e1aa491aac9b150b9bac1cccaf9d3a4ddade783f168fb7605260f8918e021ad2ae432f13a73424249e14ff6552a5b0460436487675d6a846c886de96d876d0c6c056a6267d763dc5f7c5b8a566751244ca9462441a83b2d36c030782b64265721691cd3175313010f330b8a0722046701eefeddfca1fbb0fa22fa5bfac6fa7efbdbfc35fea0ff6c01020387044906ba07fe084b0a3a0b0e0cee0c7e0df00d460e3f0e1b0edd0d560db10cc60b690ad208f106bf046402bfffcafcb6f990f67bf39ef0efed6eeb2ae934e7a0e564e487e3e9e25ae2fee1dee1dee136e2d8e280e372e4bfe53de73be9a8eb2eee02f114f428f782fa0efe7a01e3043808490b460e2a11c51321163118e719671bc51c021e0e1fe71f982017218221eb211622fa21a321dc20cb1fa71e341d831bc119bf17af15d313fb113910a90e080d780b230ad10896077b063d05f803da02ba01a800b5ffa6fe85fd7afc6efb6dfa95f9bdf8e0f726f77bf6dcf56bf5fbf466f4c6f3fcf2f7f1e6f0a2ef0dee5dec84ea88e8b4e6e7e409e34ee18bdfbcdd24dc93daf0d866d7bad5e5d330d280d0d4ce50cdc9cb48caf7c8cac7e4c650c6ebc5d3c50ac681c667c79fc80dcad2cbbacdb1cffad161d4ccd684d94cdc09df17e247e573e8f0eb7eefe1f26cf6f4f939fd8900c10387062b09a20b8f0d3e0fb7108b1105124912e7112e115710f10e510dbe0bb3097d076605d002040054fd21fab8f67af3c6eff6eb75e8aee409e1ebddb5dabed75dd5f3d2ced031cf7fcd06cc04cbf3c918c99fc809c88dc749c7dcc67ec640c6cbc549c5c7c41dc47cc3efc25bc2c7c11ec158c076bf5fbe2dbdc9bb08ba28b830b610b42eb287b0dcae8cad98accbab93abefab74ac78ad01afb7b018b34fb6ebb93cbe4fc394c864ce00d5cedb03e3d1ea90f288fa3003f20bfa149f1e212888313b3b90447d4d0056215d3063ee68cc6de471b675bc78077bf67c287ed07e1e7fa17e767d9f7bde789275bb713b6d74682e63695db957d451c94b1f464740593a0635ca2fe02af5264e230920cd1de61b7f1a1e1aea19f319a61a501b3e1ce81dad1fc2216b242427372ad72d8a316d355c39e53c3a403743a045bb472e49ce49f9496749194880462a4403417d3d3b394c34392f9e295c23e31ce315480e9806a6fe39f6b1edf9e4d9dbd3d216ca58c1f8b83cb1c4a9e1a20d9dce974093e18f1f8df38afd89b189de89228bfa8c218f4f923596819ad89ff3a56aacccb3fbbb7ec4b7cd8ad758e14feb7bf54dffd6084612181b4423352b92323739a73f8f459f4a664faf5317572b5ab25c2e5e225f735faf5e635d8d5bb45849555a519a4c80473b42933cd8363631872bf725b920c21b0b17a2127a0e670a7d06d90241ffd3fbccf8e4f542f348f1acef92ee4cee60eed0eee7ef2bf1a2f292f476f643f830fad6fb51fde8fe3f006501750221039a0307043204490454041a04cb037a030903990209022101f0ff63fe78fc58faf6f74ff58cf2c0ef1cedd8ea0be9b9e7d0e643e611e625e68de632e7cde764e802e991e968eaa8eb12edceeeddf001f38ef59bf8d3fb54ff00038006180ae10d93114815de18fc1bcd1e6621a423a025482769282a29b929392acb2a632bea2b492c6c2c6a2c342ca62bbe2a4c294027e3244022631f931cbc19d8163714d111a20fda0d370c850af6087007ed05a20462030802b8005fff03fedcfcd3fbd1faf4f92bf979f817f8fef711f855f8b3f811f981f9ebf92cfa3dfaf7f949f95df835f7d0f55ff4d3f226f19bef31eed3ecb0eb9bea61e928e8d6e649e5b0e3e4e1c8df94dd3fdbd3d895d676d475d2ccd067cf52ceb7cd69cd64cdb4cd2bced6cebccfb2d0cdd1fdd223d47ad5fad691d887dab0dce6de83e15fe449e7a0ea21ee7ff117f5abf8e4fb22ff2d029d04d706cb08290a5e0b6e0cfd0c680dcd0dd00dc30dc30d520d9f0ccc0b5b0a7b086d06bb03980060fda5f9a5f5dbf1d7edc5e920e65ee2a3de67db1dd8e2d427d262cfbdcca2ca84c88fc615c587c324c235c12dc060bf0abfa8be9bbe18bfa3bf96c003c261c3f0c49dc6e8c70cc9f1c945ca57ca2ccaadc932c9aec80ec880c7dfc631c68fc5b9c4bbc392c2ffc04cbf95bdb6bb19bac8b87db7a0b631b6dab5fab58ab62bb752b821ba51bc57bf49c3adc7c7ccb1d2e3d88fdfcbe6eded14f587fcd403470b5f139b1b1324222d2036063f2648b8508258cb5ff3650e6bb46f847398765f796c7be17c1f7eba7eae7e027e487cab7951762d72a96db8684763ce5d21585352ef4c7447c441523c82368630272be225f820161d87198716bb14591382129512a512d7129a1346142f15b3163c181d1a9d1c581fa1226a26282aee2d7131613410373e39c73afb3b803c5a3cf63bfd3a7f39cd376b3561320b2ffa2a3c262c216e1b0c15750e7c071d00b0f80ef100e9d6e0aed854d01fc85bc0b1b864b1edaae8a47d9f389b8397519438929b905b8f278f778f2a9001929394af970a9c42a103a7dead8bb599bd61c6adcff6d876e235ecc9f553ff05096b12701b6b24f02cc6346e3c8b43c549b74f1a557a597c5ddf602063ec6418661d669a656364f361d85e135b58563751d04bf145fc3f063af833ff2d35289b22241dd317ba129d0d8808c30303ff71fa82f6d8f29bef55ed8ceb4eea17ea45ead3ea27ec96ed1cef25f115f3fdf447f77bf9b6fb4efecb002d03a905de07dd09d90b8a0dfe0e491044111412e012a4136c14131568155315b914a1131a122310db0d5f0bd708870694040e03fa012d01a10050000700c0ff55ff7efe65fd25fcd9fa04fabbf9cbf968fa62fb7afc09feeaffd301f303fc05bb07a409a30b9a0dd80f14121e1447166418541a3c1cd11df31ee91fc120aa21db2225246d25ab26bf27bf289b291e2a392abc29a22836278725b82307224d20921e191dc81ba51ac619ce189b175116c7140c135d11850f720d5d0b3c092007430579039f01deff2cfe8cfc48fb4ffa64f99af8d9f7f9f629f659f546f406f385f19aef94ed91eb77e984e7c6e520e4cee2cfe1e5e017e03cdf1fdee4dc9cdb40daefd89cd734d6d0d488d374d2a2d104d198d04ad01cd041d0b7d07ad1b0d22bd4d2d5d2d7efd9f7db17de05e098e132e3bae41fe6dce7d4e9d8eb5bee30f1fef312f71efaa1fcf9fe09017202b203ce045705ca05390633062b063406bf0528058e046f03340216019dff26fee9fc69fbeaf987f8a5f660f4e9f1ccee6beb28e8b7e470e192dec9db70d9aed71cd6e7d4fed3dad2a0d15ed0c9ce2ecdb8cb2ecae2c803c853c70ac72bc74cc78bc7fac750c8d4c8aec98bca9ccbf2cc2ece84cffdd01cd2fbd294d37dd305d354d23ad121d028cf23ce75cd0fcdb2cc8dcc42cc7ecb65caa9c851c6bbc3bac0aabdf7ba54b824b6a5b449b375b24cb228b285b27fb369b4e6b51cb878bac1bd10c2a5c61ccc64d291d823df2ae6eaecf0f38bfb4603a00be1148f1ec1282833be3c9e45424e1056c95ccc62c867b56b376f3972bc74487793796f7b3d7d897e087f067f117efe7b357982750771246cb7660c61485b38554a4f5c492343313d48373d31e62bde260322331ecd1ab417c3151c149812f311231134100510b90fa40f9a10ba115b130e16ec18431c3f20f923c827962bb32e9e3116349c35c9364a37f8369336b4355034ef32e1303d2e962b49289224dd206e1c69171d12020c60057dfe03f734ef4de741df4fd7a2cf52c85cc1c8bae5b492afb9aacca66da35ea02e9e6f9cf99a849a809ab19ad79b6b9d559f70a246a6b6aa5bb0aab674bd35c584cd1fd62fdf4de822f1b3f9fd01e8097111d8180220ae26482dad3377392e3f974428498b4d7f516a54f656d35865596d59b858e056ae54ed513e4e3c4ac045a940983b8e369131dc2c4528d3236e1ff61aa7164012b40d70091005a100b5fcd3f82bf55ff2f6ef18ee4fedfdec16ed11ee3bef9df0b7f2dff40ef79bf9e3fbf9fd52008e02c50439078809bd0b200e9a1049134a166919821c6e1f0e2257243426a7279528dc28ab281a2827270c26cc244f23d7218420621f8d1ecb1dc51c561b701948171515e012b010450e6c0b5e08300513026dff12fdecfa3cf9c3f787f6e5f582f544f577f5c4f51ff6cdf659f79bf7d2f7cbf7c1f739f826f98ffa80fcaafe1101c803b806e609200d2410e2122415fa169618d619e81afb1bc21c6d1d211e691e6f1e681eee1d481db51cb51b6c1a0f1934171a1500136610510de009a805e4000cfc07f71cf2a6ed6ee97ce50ee2e8def2db45d996d6bcd3e1d0e5cdb7ca83c769c474c1f8be38bd1abca5bbb0bbe7bb38bcabbc52bd56bebebf77c166c368c580c7aec9dccb24ce67d06fd26ad44fd6fcd7d5d9e8db12deb1e0aee3a6e6c6e9b7ecf3eebef004f28cf2e3f21af3f8f2fff22df337f38af30ef454f49cf4bdf44bf4a9f3eaf2c6f1a1f094ef5bee46ed65ec65eb7eeab0e992e858e71fe6a4e43ae31ee214e171e064e086e0e8e07be1aee199e15ae1a5e0e1df46df77dec5dd53ddcedcacdc15dd96dd6fde7fdf18e07de0b2e043e0addf12df1fde6cdd0edd8bdc49dc33dcbadb5ddb39dbe5dadcda12dbf9daf2da02dbc7dac8da12db24db41db55dbf3da84da2bda9fd93ad90ad9c8d8bbd8dcd8dfd8e9d8cfd841d882d78bd654d533d4ffd2aad162d0f6ce7acd1bcc8bcae1c840c75cc59ec35bc239c19cc0a9c0bbc036c150c264c3d1c4a0c60cc895c98ecb90cd67d06bd4fad886de16e5e0eb2bf3ecfa6102cb093f113f18351f6626812dd334853c2a44da4b9a53dc5a7e618667926ca1700874ad76b0786b7ab47b8a7c247d2f7d7c7c1f7bcb787c757371a26c4967a961bc5be1552e50824a2945f13f9c3a83355b30102b2f2645214f1c091803146e10240e770c590b4c0b560b710b480c150d130ed70f86115913c115f017391af01c5a1fcd216b249e26c528be2a042cf32c532df52c6a2c6c2bd029f7275c25f921511e071a40157b10470ba705ecffcdf956f3c9ec2fe678dfd6d883d24fcc49c6abc03bbbe0b519b1b6ac91a84da59ea243a0009f7e9e759eb69fc6a12ea4aba7bbabe5afe8b459bab7bfacc5fbcb4dd24ad9dde093e8abf00ff94a017309b511b6194e21be28b82f0336203cd241af46354b254f045286549b56be578c58e25833582157b955a8536951e44ec34b51487c442a40923ba4366f31052c80264121281c26179812150e9409ba052402cdfe54fc10faedf79af670f56ef446f43cf44df430f53af65af713f9bbfa5ffcaefe60019904b108010d3d1166150d193b1c251fa621c52391250e277228e129672b042d8b2ef62f46314f32fa320a3320324430c12ded2a3628d4259a234321b71ef41b0a193816731389107a0d600a4a0774041e0204000bfe5cfcb3fa12f9bbf74af699f4fdf260f10cf0a8ef01f0ecf08bf265f44cf680f8b0faacfc80fedfffe400f8013503cc04cc06ec08210b610d9c0fec111614e81563174618b41806190919de18c5185c18c41737171f16781473129f0f510c2109d2059e02c5ffbefca0f9aef68af350f032edcae91de65ae24bde19da11d63dd2ddce32cc3ccae6c806c85fc7c2c62ac6b9c57ec57cc5bcc515c66ec6f5c6bac7c1c828cadacbb3cdbacfe6d12dd496d61cd9b2db52de08e1d7e396e635e98eeb62edddee24f01ff120f23ff333f449f597f6cbf737f9cffaf2fbd8fc89fd9dfd9efdc1fda3fda2fdb3fd5efd1cfdfbfca0fc77fc64fcecfb68fbd9fa07fa6bf918f9e4f820f9aaf924fa95fab3fa3ffa72f956f803f7c8f5b0f4b4f3f5f271f218f2fcf120f251f26af261f2f7f10df1d0ef40ee87ec17ebf7e92ae9dde8a1e829e891e790e64ae53ae431e344e2b2e110e18ae085e0a6e01ce100e29fe2fde222e392e2bee1f1e0dcdf20df03df31df1fe0b5e146e3f4e483e670e730e8bfe8bce880e8ede7c4e680e547e420e35fe2d6e14de1bde0e9dfe9dedddda2dc5cdbf9d946d89ad6f5d43dd3d7d189d012cfdecdbfcc9bcb0dcbceca87cab3ca21cbafcb25cd83cf79d26bd60fdbd8df22e5dcea86f061f659fcd9014407000dc7120e194120d727e62fac387b41404a1a532d5b4862b168cc6da971ec7477777179337b7c7c797d6c7e037f317fd57e917d7c7b8c78c57474706d6bc665e15f7a59da52844c0946a53fae396f33322d75279421051c4f17c012c70ed00b0d09df0687052e042b03a902f40184019501a20126024d03b404d406b209e20c92106114c817d81a3c1dda1e0b209a208a2025202e1fc51d441c7c1a9418c416a4141712300f950b4107760221fd4cf742f110eba7e43aded6d73fd1aaca62c43cbe6ab845b374ae06aa6fa66ba323a119a0da9f28a046a1aaa21aa413a660a8e2aa29ae26b29fb608bc69c26dc950d111da27e385ec2bf678ff4f08ec10dc181d203527c52db933ab393d3f40445a49264e4d525456cf59525c515e835f995f0c5fbb5d6b5b7858dc547850984b5e46e040523be635af309c2bcb264422b41d3a19f5147410d80b5f078b02a4fd2ff9def422f190eeafeca1ebb3eb3eec45ed11ef19f163f329f6e3f88ffb68fe1f01ce03b7069a09750c640f3812e7148017ef19361c601e6d20592213248725972621272327a1268925df239a21a41e051bed168612080eb3099d05be012efeeffae3f72af5c7f279f03fee0ceca1e922e7b5e449e228e086de49dd9edc94dcf4dcd4dd3bdf01e130e3bfe584e877eb81ee97f1bcf4dcf707fb38fe3e012c04ea063409340bee0c380e630f7f1057112a12ec124d138a139f133a1386127311aa0f5b0da50a6407eb037700e8fc69f921f6e2f2b1efa4ec85e944e605e3b8df66dc52d979d6e0d3c5d120d0e8ce46ce0cce08ce4cceafce23cfd6cfbad0c6d10ad35fd4ced577d74ad969dbcfdd3be0b2e214e529e723e902eba0ec3feec5effcf024f21df3b4f336f485f47af460f41cf48ef307f372f2b7f120f1a0f01bf0c1ef73effdee73eec4ede4ec0eec5debc7ea6cea56ea6eeacbea84eb73ec8fedcaeed6efb2f082f12af2d9f2baf38ff46ef575f65cf74ff868f947fa06fbb1fbf1fb15fc4dfc52fc6ffcacfca4fc9afc8efc19fc78fb99fa26f97cf7b8f5bdf3f6f162f0c2ee4cedeeeb83ea47e92ee808e7eae5b8e463e31de2f4e0ebdf1edf89de0ade98dd3eddf4dcc5dccfdcfcdc47ddcddd65de10dff4dfd5e0b5e1c1e2b1e39be4afe585e63ae7fee767e8c7e868e9cae92feaa9ea88ea2deadde921e991e855e8bce72ee7b2e6bfe5f6e47be4c6e340e3bee2ade17be01edf50dd82dba4d992d7aed5ecd351d212d1f5cf05cf51cea0cd2acdd3cc38cc90cbabca5ac948c877c7b5c695c6d4c617c7f3c72ac96bca44cc57ce3fd098d252d54bd830dceae005e6cbeb0cf23af888fedb04a20a091052154c1a711f5225a82b8a32353a0742ca499b51bc58d45e15640c68d96a2a6df36e6770e6711973f1739074a87446746973d371ad6fea6c8869ec65e961815d16593954f74ec3490244ca3da9371431772abb24621fca1a8817ad144b12d710660f230e770d710c330b270ab2084807880611064b0686074d09ce0b140f9e126e16541ae21d2521f2231e26d027d9282d29fd282128b126ec24b4222b20921dd51a091857158912730f0b0c22088f037afe06f922f308edfee6dbe0d6da56d522d05acb63c7cdc38cc00fbee6bb17ba3fb903b952b9b2baa5bce1bed3c109c541c8ffcb13d054d44ed9eedee9e48debbaf2fdf97e014409da104818941f32260c2c6b311136293a473e3542e745b4493a4d49503553ae557857cd585859ea58c557ca55fb52974f9f4b35478f42c83d0e395b34ad2f312bc5268e22ea1e991b9d182816ac131c11c50e2e0c6e09f4065204c601e6ff68fe89fdb8fd71febbffdc015b044307b90a290e6b11811404171319ed1a761cdf1d401f6d207d216b2212238623b52386231123442206216c1f601de11a2b1861159712fc0f7e0dde0a0b08f1046a01a3fdd0f9ebf528f2c1ee99ebcfe892e6a8e415e3f8e110e15de006e0d3dfcbdf27e0cbe0dde198e3e0e5abe8e6eb3eef7cf276f50ef84efa46fc21fe0900f8010c0450069208ea0a5b0d910f93114e135b14de14f6146d148f1386120a114f0f750d350bc00830063603f6ff9afc0ef9a5f5a7f2ffefbdeddaeb0dea43e87de69de4a7e2b4e0c7def6dc6edb47da8dd954d998d952da86db23dd08df07e1e1e272e4b5e5b8e6b9e7e6e841eaddeba4ed66ef37f112f3d2f496f649f8aff9f1fa07fcc1fc56fdb3fda0fd5efdf5fc4dfcbafb36fb85fad5f916f926f85af7c1f63af6edf5b6f54ef5d0f42df44af35cf26ff172f099eff2ee68ee1fee1cee44eeb7ee8cefa3f008f2abf336f591f6baf781f814f9b8f954fa12fb0ffcf8fcccfd96fe02ff30ff59ff45ff2dff41ff23ffe6fe99fed9fdcffca7fb13fa3ff841f6c6f309f148ee6eebdde8cee60ae5a4e388e255e10ee0b6de23dd8cdb1edad3d8dbd750d708d70cd75dd7d0d770d850d944da52db8adcbaddfade67e0cde138e3b4e4eee5fee613e8f8e8ebe920eb36ec50ed80ee4eeff5ef9ef0d2f0ddf0e0f05cf0aeef04efededdcecf6ebbeea9ae99be844e707e6fbe4c7e3e5e261e2dce198e15ce1b3e0c5df6fde98dcaadab8d8e4d674d548d474d30ad3d9d211d3a9d349d419d5e2d541d693d6c4d69fd6b8d602d740d70ed847d98fda61dc74de4fe075e2cee413e7e7e94dede9f038f52ffa57fff804ed0a8210c715b81af01edf220527402beb2f6235423b99419948ab4f8356045d76629f66c269ca6b036def6d896ee66e296f206fc56e0d6ec96c006b936882650662f85d6d59a6544f4f9749e843e83dca37e2318d2bf924a91e381834124d0df80874050e03f40051ff71fe95fde9fca7fc2bfcc1fbc8fbe5fb80fcddfd9bfff801fb043508b70b470f7a126715ec17fb19e11b801dca1ede1f6c206220eb1fcb1e161d051b6a1863153012b60e0c0b600788036aff06fb31f6c2f0d7ea9be421debdd7d3d15ecc7ec77bc316c041bd41bbb7b970b8b3b721b797b690b6e0b66db7beb8abba06bd4ec068c400c963ce56d45edab2e048e7c8ed7df487fb83029009c810aa17281e6324df298d2ebc322136ca38343b423d063f04411443124533470c49374abc4a464aa7482146c342c63e8f3a5b366132bd2e6f2b7b28b7251923b1203a1ea51b111937164013a3103e0e4f0c2e0b680af009f509f209f0093b0a6b0aac0a6b0b600cbc0dc20fee1127146e164518b819ed1a9c1bef1b151ced1bc81bdf1b111c791cf61c2c1d1f1dae1ca61b231a07182a15ce11180e300a84062b03050021fd53fa6cf790f4b7f1c6eee1eb0ee94de6e9e30ce2b6e0fcdfc2dfcbdf03e049e06fe06be02fe0c1df66df6cdf2ee0ede19ce40fe8ecebbaef44f35df6cdf8adfa0bfcd2fc51fdbafd07fe7bfe1fffaaff3b00cc001301320125019800b1ff8efe0ffd7efb03fa64f8b3f6eaf4c5f267f0f2ed4eebade842e60ee44be22be19ae092e0f8e085e122e2c2e240e395e3afe368e3cde20ae255e111e188e1cae2eae4bee7ecea48ee83f13af461f6e6f7b3f81af948f93ff948f972f99ff915fae0fac9fbebfc11fecdfe27ff12ff75feaafddefcf9fb23fb46fa15f9a3f7fdf517f442f2b7f070ef86eeeced63ede1ec6cecf5eb9eeb86eb8ceba8ebd2ebdcebcdebcdebd9eb11eca2ec6aed6beeb1eff9f046f2b1f304f55cf6ddf73cf97dfaa5fb56fcacfcdbfcb3fc78fc58fcf0fb53fb89fa36f9a1f714f666f4e8f2b0f154f0e3ee54ed54eb25e9eae679e409e2a6df1cdda3da56d830d675d43ad360d200d2fed129d282d2f1d255d3c5d34bd4e8d4c6d5f0d655d808da05dc2dde91e027e3ade51ee865ea45ece6ed6fefbdf00af270f39df4bff5eaf6bef76bf8fbf8f0f885f8daf797f633f5f0f375f22cf12cf0faeee0eddaec68ebdbe942e851e683e4f7e26de136e047df5edecedd9addabdd2bdedade70dfe1dff2dfc7dfa2df89dfc2df4ce0e0e0a7e188e24be350e475e567e673e758e8c7e835e980e970e99de9f1e940ea1feb5bec82ede4ee3af03cf195f279f4d1f61dfa2afe5d02cf06540b830faf13f217f81b032045248128042d11325c37033d24435a49944fc5555b5b1f600764cb669868b969336a396ae8692d693268fa668465f7631d62e45f645d455a81564152194d2f47f7403b3a7233332d12273f210b1cd216d611960d8c0906066303f100e3fe90fd5dfc81fb49fb19fb1ffb9ffb25fceafc1efe53ffbe009302a7045107af0a720e7e127516e119b41cc81e1a20ed203a210a218d20a01f3f1e8b1c601ac617f414e911b90e910b5408e104440178fd6af941f511f1a9ec02e836e322def1d815d48fcf81cb57c8dfc50bc439c327c39bc3ecc4d2c604c9e9cb4bcfccd2b6d6c9daa0deade207e782eba1f074f689fc13030b0afb100b18451f2426a22cba32f637693c4c406943e8451448c449174b4c4c3f4dec4d644e6d4eee4de54c314be14800469842d33eb13a4136b431fe2c4f2803240f20981cd91974175615b0132912c710d60ff30e160e890df10c660c4d0c5b0ca80c9f0d0e0f1c1113148417261bd61e0922b0240427e028612a962b2c2c312cca2bfc2a1b2a4a295d28632737269b24b5227720af1d901a0d170613bf0e2f0a2905e5ff67fab3f449ef71ea37e6dfe252e03ade97dc51db35da5bd9bfd82ed8b2d74fd7f9d6dbd620d7d3d70bd9ccda08ddb2dfb8e212e6a6e94fed01f19bf4f0f708fbd0fd1900f2014c03fd033e042704a303f702360235012e0036ff1efe0bfdfafb98fafdf838f723f5f9f2dbf08fee26ec9fe9d1e6f5e34de1e7de01ddafdbc1da34dafdd905da75da63dbbadc79de6be045e2fce381e5cbe611e85be99eea03ec8bed2cef14f13af36ef5c6f72efa80fcd8fe1401db0215049b04480481039c02a201bc00cdff6dfeadfcc0fab8f800f7d6f5fcf46bf40af485f3e0f221f202f189efcdedb0eb75e962e766e5aae352e244e1c3e00ce100e2a5e3c9e5e0e7c8e977ebc4ecfeed56ef96f0d6f10ff3f3f3b0f465f5d9f53ff6a7f6d1f6f9f64df790f7e8f74ef859f81ff8baf7f8f613f61ff5c8f316f219f0abed18eba9e84ae61ce41ee215e011de20dc2fda64d8ccd658d536d47dd32bd35cd3f4d3c2d4cbd5ffd65fd81fda23dc2cde20e0b1e1bbe293e377e498e559e7abe94aec44ef71f290f5d1f812fceafe65015d037704f404f00437042c030902a90078ff9bfea6fdb3fca8fb0ffa37f86af686f4f1f2c7f197f06def35ee8becaceab3e86de622e4f8e1d9df29de20ddbfdc3edd79de1be0fee1cce34de58be672e70de877e89ee8b0e8d2e802e984e952ea29eb1dec01ed92ed19ee87eeb2eef3ee29ef1eef35ef47ef11eff1eebeee3beee6edb0ed60ed5bed79ed7aedebedfceeabf08df391f729fc4c019e068d0b4810e4142419501d872186258829cd2d2c32e8363e3cef41f5474a4e6e540c5afa5ed762956569676968c2689b68ed67ae66e364a66221605b5d745a6157c5539d4ff64a9745d63f063aeb33c72dcc278521341b2a15000f1909d703c5fe36fa87f63af39cf0fbeec5ed26ed41ed72edd9ed98ee2aefcfefc0f0b2f106f3f2f439f718fa7afd0601d1049f08190c480fda118e139814e31491140e1444132712d310ec0e5e0c6909fc053b026ffe83fa75f666f247ee11ead9e599e137ddb3d826d48ccff4cab3c6dac27cbf09bd8cbbe4ba5abbb1bc6fbebfc06ac30ec616c986cc0bd016d4a5d855dd91e26ae875eefcf4f1fbc40299097810fa16541da0237029c72eb233d837503b573ec0409b421344fb445c456d4527459744e7430043d3416140873e2c3c4839d335f231cc2d95299a25e021631e441b59189f1562138511ff0f060f460e970d4e0d400d7a0d680ec00f4a1134130d15ab166718001a711b1b1dc11e6d208122b92404277a29972b362d712ef72eec2e812e712de42b092ab8274b25ea225120a71dd41a8a171914a2100a0da5096b061303d8ffb4fc7ef97df6a1f3b1f0e4ed3debb9e8b5e64ee571e43be487e421e510e63ce78fe81cead6ebaceda8efb5f1bbf3aff573f701f96afab8fb0efd8bfe15009c0109032304e3045d057e055705f3042104e4025b0175ff5ffd4bfb15f9bef658f4b9f1feee5fecc9e95ce759e58fe3e2e162e0d2de3eddbddb2bdac3d8bdd716d704d785d751d870d9ccda31dcd5ddc3dfc7e1fde34ae669e878ea70ec29eed4ef6df1c9f21bf465f585f6b3f7eaf8f0f9ddfa99fbe1fbdbfb8bfbcafad0f9a5f814f745f54af305f1c1eeadecb7ea23e9f8e7f3e632e695e5c6e4f3e320e31be244e1b5e033e0f9dffddff8df39e0c9e077e192e2fee360e5fde6c4e871ea5aec68ee2ef0d4f12ff3edf368f4baf4caf404f57df507f6d9f6d6f7a0f848f9acf995f948f9ddf83ef8a2f7fdf603f6c7f44df375f177ef80ed95ebf1e9b3e8cce752e729e710e707e7ede685e6f5e546e557e474e3cfe256e243e2ace247e310e4f6e4d0e5b8e69be79ce8bce903eb83ec31ee23f006f2e1f38cf5a5f674f70cf825f830f850f820f801f81cf803f802f836f81ff8f1f7c6f72af757f66af5fdf34bf27af042eefbebe6e9d0e7fee597e462e38ce21ce2c3e187e14ee1cae01fe06cdfb5de4ade46de82de14dfe6dfc4e0d5e116e350e494e5cee6cae7bae8c7e9edea5dec0eeeb5ef35f16af218f33df3daf2e9f181f0daee3dedceeba9eaf6e978e9f2e88de806e81fe71de6c2e4e2e216e160dfc2dd0fdd1edd78dd9ade13e040e1c9e2a1e477e626e9bfeccff0f6f515fc8002970931118c18da1f0d27852d84334f39ad3e0444d749fc4f8c56ae5dd064776b807158769e79987b417c8b7be4796a770b7424700b6cc66789635f5feb5af9555a50fa49d5421f3b3d332f2b1623651bed13ab0c1106b9ff95f93cf45bef10eb10e8eae5a1e4c2e4aae558e73cea91ed32f14bf504f95efcacff98029f052a09fb0c72117b16a51b2921a426ab2b723066343c374b39203ac939d138d7360a34de30dd2c39285623d31d06185c12920cec06a0015ffc21f7caf11dec13e6abdf21d9a5d25dccd1c61fc245bed2bba3ba75baafbbd0bd50c08cc313c79dcad7ce77d347d8e0dddee3efe994f084f770feaf05f80cf413d91a9221f1271c2e2234c639f13ea84393476a4a424cd44c094c6d4a1e485645d14278401f3e153ce3393f3778344131832d8a2922256a20a21bcc1672129b0e680b4e09e7070e07e90605073207f30702095c0a920c250fed11431585189d1bd91eab213d24e7263929812bf02df92fe931ce33353580369b3706380a386337ba359133cc30592dd1290e26f621f11dbc193e15c510ff0bea06e201d4fceff786f37fefe0ebbde8f7e596e39fe104e0bddeabddc3dc07dc6cdb13db1fdb9cdbbcdc90de04e11ce4ade76ceb2cefb6f2eaf5c1f838fb6dfd6aff2901b802070415050b06e406b8079f084f09a809a809ff08b5070a06ec03880112ff63fc9bf9ddf608f448f1b3ee33ecf5e9fee72fe6b9e49ae3b3e224e2dee1cae1fde164e2f2e2b3e389e480e5b7e62ae8ece90eec67eed4f048f3a8f5ecf722fa56fc6efe71005d021504a505df0686077707b10645057a03ae012000f4fe2dfe9ffd19fd75fc88fb37fa76f835f687f3a4f0baed09ebc9e80de7eee57fe5a6e549e640e73ae8fce876e9afe9f4e99beac4eb76ed8eefb8f1ccf3bdf583f74ef93efb31fd26ff0a01ab0219047105a606dd072109310af80a510beb0ad9094a08440628045402b6005aff39fef8fc8afbfaf913f8f1f5b6f331f17feee3eb5ee934e7abe59be4f4e3a2e346e3cae238e271e1a2e008e09bdf84dfdddf72e03fe136e216e3ede3c4e474e51ee6d3e677e737e826e91cea2ceb3aece8ec32ed0eed56ec5deb69ea7ae9dfe8aee89ae8aee8e0e8dce8c6e8b1e84ee8bbe705e7dee58de45de343e2a4e1c9e15de268e3bde4b4e542e66de6f3e54ae5d4e47ce4a9e47ae588e6f8e7b1e930eb8eeca8ed0dee06eeb1edf1ec54ec0aece8eb42ecf7ec9aed47eebaee93ee0bee1fedd0eb9deaa7e9efe8a9e89ce88ae86de804e840e73ce6dfe459e3d1e13de0dcdeb8dda6dce5db68dbfedafada42db90db33dc05ddb9ddb8deebdf07e17ee239e4e6e5f7e766eadcecceef49f3fff664fb8f0018063c0cec129c195f203027932d923343394c3ecd421c47274b2d4f8b532258dd5cb5613d660c6aeb6c916ed56ecf6db06ba768eb64c9606d5cd8573f53b04ede49d5448e3f9c392d338d2c8225751edd176611510bf605cf0005fcfef740f401f1b5eedfeca2eb69ebbeebcdecfeeedcf165f5b2f917fe6e02be069b0a270e9811c314e3170e1b101e0c21e9237126cf28d82a5b2c782dd42d262d922bda2807259820961b1b1683109f0a4f04d9fd34f76af0e0e9a8e3acdd0cd8bcd288cd8ac8fcc3e3bf6bbce1b91cb8e2b64cb615b614b6c4b647b89bba3abefcc25bc86fcee7d43edbaee131e887ee03f599fbd701fb07090ea8131819621e23236e27442b582ed430ea328134bc35b1361c37e236f53521346931fb2df02984250e21c21cd7188115bf128310b40e1b0d970b120a7908e3066c052c0465033e03c2030b05f2063009aa0b2f0ea3103b130116f2182d1c811fc322062623290e2cd32e2231cb32c333cc330933c431f52fdb2d9e2b032927261a23931fc21bbe174f13c60e4c0aa70512018cfcbff7ecf23bee94e960e5c7e191deeadbd7d921d800d784d682d611d723d883d93edb4cdd92df16e2cee4afe7bdeaf7ed61f1f7f49ff859fc1100a8031e07540a150d570ff910db112412e8112f113510160fc30d590cdc0a2509380716059502beffaafc4af9c1f548f2e8eec8eb16e9b7e6abe404e39de177e0acdf16dfb4dea1dec2de2edf11e05ce11be34ee5bce751eafdec87eff5f148f462f667f865fa3ffc0dfec2ff2b015d025403f40362048e04450493036902ba00ccfec0fc9dfa8ef882f655f41cf2d7ef7eed3deb19e90be73ce5b0e35ee263e1bfe05be04be094e024e108e236e380e4e1e54be7a5e813eab3eb7ced9fef28f2e9f4f2f72bfb34fe0001740341058b067207db07140849084b084b084f0802087f07c3067e05eb033802380038fe68fc84fab9f819f759f59cf3f3f112f014ee13ecdce9aae7bae5f7e38ee299e1dbe05ce027e00be022e088e014e1c0e182e21fe384e3b7e3aae384e375e38ce3e6e392e46ee562e649e7f5e764e893e87ce84ae808e8aae74ce7e7e665e6f0e588e51ae5d5e4b5e499e4b3e4f6e436e59ee517e672e6eee683e706e8c4e8b5e9a5eae4eb75ed1bef15f14bf35cf57df7a8f990fb79fd5fffea0052028d034c04db04470542051505d5043f04ad034203b3023102b601dc00c3ff70fea0fc8afa49f8b4f511f37cf0d2ed42ebe8e8aae6bae43be32be29de17fe1a0e1dfe11de256e28de2c1e20ae359e395e3e5e33ee497e43ce518e606e74be8bce912eb97ec24ee77eff3f080f2d1f340f5a6f6a6f7a2f88bf919facafaa4fb53fc46fd83fea6ff1501ed02e9047d07e10ac00e47136a18971dbb22c327432c54301a346a37753a793d68407443c8463f4ad84d8d512a558c58885be65d7a5f0b60935f245eaa5b4e584454794f354ad4444b3fde39d134c62fce2a1a263a214a1c93179a12750d89088503b3fe99fae3f6b3f35df168efeeed59ed5aed1beef3ef79f2b0f5c4f938fef5020608f00c9c111416051a7d1d8c20ff220025a726e1270229232a1d2b0a2cbb2cce2c3e2cd62a5428e5248e20461b7215500ff008af02a8fcb5f6f8f07deb1be6fce054dc07d835d411d16ece5acc1ccb91caadcaafcb62cd8ecf65d2b6d549d967ddfae1d9e65bec6ef2c4f884ff7306210daf13fd19bf1f2b25362a8d2e5a329c351a380c3a873b5f3cbf3cae3cf43bab3ae03873369d338b30422df029962616237b1fa71ba417c6131c10b30ccb094607150577036102de0131022b03b604f4069d098c0ce40f5513bd16531ad41d2521782487273a2ade2c5c2fd03188344337d839443c1a3e363fad3f403fff3d0e3c31398d356531a22c902776223a1d1c184513760ed70981052d0110fd54f9c2f591f2e1ef56edfbeae2e8cbe6f3e4a7e3cae295e239e372e448e6e1e8f0eb64ef50f35bf74efb25ff930275050008330a1e0c040ed90f7a11ee121714da1452157e155115e914451450131a12b210130f550d950bd709150854068704920279004ffe24fc20fa7af846f7a3f6a7f633f731f89ef955fb3ffd4cff410102039004d205ce06ae0782085b09510a540b590c5c0d3f0eef0e6a0f980f6b0fef0e270e0e0da50be709d1076705bc02e8ff0cfd3bfa80f7e9f47cf241f04aee95ec11ebbbe985e86de78ce6f3e5ace5c2e51de6afe67ee774e896e9fdea93ec5dee64f083f2c7f43af79af9defb08fecfff400179023f03ac03e303aa031b038202b101d000190024fffcfdaafcc9fa88f814f62df31ef024ed02ea06e761e4c5e16cdf7cdda2db12dae6d8c0d7c5d60ed64ad5b2d478d465d4a7d454d515d6e7d6c5d761d8d7d859d9d3d971da4adb17dccadc5add9cddafddb0dd8fdd67dd34ddcddc51dcbedbf5da1cda36d92ad833d755d672d5c2d439d4b1d373d37ed3a8d32ed4efd49dd577d674d767d8bbd978db53dd85dff8e151e4d6e680e9f8eb79eef5f016f31ff51bf7cff88efa63fc01fea1ff330152022503a903960335039e0291015200edfe19fd25fb32f905f7eff406f3edf0ceeeb5ec4ceadfe7abe570e374e1dddf37de9bdc33dbaed949d85bd7a5d64ad67ed6e0d673d779d8b3d932db29dd53df80e1bae3b9e54be79ee8ace962ea02eb9eeb09ec57ec99ec9bec63ec28ecd5eb5eebfaea8eeae9e93fe98fe8b0e7eae64be681e5c3e428e45ae3b1e280e282e208e36ae44fe6e7e890eceaf004f620fca90269097a104b17ab1de923b629012f29340139793dee4151468c4ad24efc52ba56ec59525c945d935d565cd7593156b8518d4ca64646408d395032e42a8f231e1ccd14cc0db606b5ff1cf9a9f2adec99e71ce353df83dc33da6ed891d744d79ad7f8d80fdbdadda9e132e661eb6cf1fef7e0fe0b061b0dcc130e1a9e1f62246d28b82b572e6830ec31f13275336b33d932ab31d52f562dfb29ae259420ab1a1314240de50557fecef644efd2e7e9e09fdafed42bd020cca6c8c5c597c307c22dc14ac14bc219c4e4c67fcaabce93d317d9e9de3ae5eeeba5f28ff98f003d07d80d67148e1a88204426342b6a2fce32e934003646368535183426326e2f3d2cc428e424f320151d1619171501118f0cea0722033efe9df966f5a8f1aeee82ec1febafea1beb51ec67ee3ff1cbf40df9cffdee025208cc0d5313f018891e1a248129892e27334737d33ae03d5240fb41e142ec4213428f406a3e9b3b4c386234bc2f862ac124581e901781101d09c1019ffaabf32bed35e78ee15ddcc0d78fd302d03ccdfcca6ac9bdc8c5c8aec9a8cb63ced2d1efd54edadadea7e371e835ed13f2cff659fbcdff11041008f00b980feb12e1155218151a1f1b731b101b081a9318cb16b9148c123a109c0dce0acd079204680172fe9dfb1ef9f6f6fef465f33af261f102f11ff17df11ff205f318f478f539f74df9bafb74fe5a0153044607190ab00cf20ed21043124713eb132114d9131913dd113310440e240cdd097c07f9045b02adfffdfc65fae5f771f514f3bbf065ee31ec1dea35e89ce64ce55fe404e434e4f3e44de608e806ea4beca3ee0cf19cf32bf6b2f840fbaefd090067029e04af069108040a0e0bb30bc20b530b710af9081f070405a4024300edfd77fb05f999f606f483f125efc7ec8bea73e860e682e4efe28ae17ce0cadf4bdf19df45dfb1df6fe07fe1b7e220e4bbe564e71ce9e6ea9dec3feecfef37f18ef2e1f321f55af686f77df832f993f979f9f2f806f8b0f620f56ef390f1b5efebed24ec92ea37e9f6e7f3e626e66ee5f3e4b3e48ce4aee416e5aae598e6d1e725e9aaea43eccfed7fef50f129f336f567f7a0f904fc84fe08019d031a064b08350ab90bbd0c5b0d8c0d470db20ce20be90af3090e09240837073406fa04970315026500a6fef6fc4ffbd1f99bf890f7b6f60ef671f5eff49bf458f43cf455f479f4b9f428f5a6f556f644f743f858f96bfa39fbc4fb02fcdbfb7dfb06fb79fa07fabcf98cf98af9a3f9baf9c0f98bf902f916f8bef61cf545f34bf16fefb7ed1cecd5eab9e99fe8bbe7dce6e1e52de59de40be4dfe3f1e311e4bbe4d1e50de7dae800eb18ed7fef15f275f4f9f688f9b3fbd6fd0e002402a104d5078c0b16109115871bf221be28602fb735b93b024189456849774cd44ec6505e52cf534755b5560b582259bf59c9590c5979572e551752514e264a7f4581408a3b6e364c317a2c9d27a822dc1dcd188a13950eb1091605560119fe6dfbc1f9a6f826f8a3f8a2f91ffb67fdf9ffd5024706e009b10d08127b16131bf01f8824c528b52ce92f7b329634f435bb361237bd36f435e8346d33af31b52f2c2d1d2a81262122331de7173712680cac06ea0052fb13f61ff1aeecf6e8d9e562e3aae177e0c3dfb7df26e009e18ce27ee4cde6afe9f6ec8af09ff404f996fd83029207860c6c11fd15fc19911daa2033236925352777285629be299b29142912287c267024e221d61e831bf51737147b10c50c2509d105c8020500a1fd79fb77f9bef747f620f58bf48bf421f57af67ff80ffb44fef301ed05470adb0e7c134718181dbe214d269c2a792efa31fc3455371939263a653a033a0a399737ee3510340032c72f362d462a052754234a1ffa1a3b162911e50b5a06d10089fb75f6d6f1d8ed4aea5ce72be57fe37fe248e294e276e3fbe4c9e6e1e851ebceed62f02ef3f0f5a5f865fbf9fd6100d10233058f07060a6c0c9c0e9510351267133f14be14d7148b14dc13be123911750f8d0d910bad09f5075306e304af039002a001f1005800edffccffc2ffddff36009100f4007b01ef015202c10207032703470344032c032a0323031d03320336031f03ee027302a0017e00eefe00fdcdfa4bf898f5d2f2f4ef1bed66eacae765e553e380e1ffdfdbdeebdd36ddcddc8fdc92dcf1dc7cdd35de23df08e0f1e001e211e33fe4abe517e78de81bea76ebaeecddedc1ee7def38f0acf001f154f14ff11df1daf032f05aef69ee01ed5deb9ce979e752e55de355e18ddf18de99dc56db62da66d9b1d84ad8d2d78fd788d76cd791d705d876d82dd927da0cdb1fdc64dd88decedf31e154e26ce372e414e595e506e629e642e65fe633e6eee598e5e7e416e43ae318e2e8e0b9df4bded2dc65dbcdd94dd8fcd69fd570d472d361d279d1c4d011d0b6cfc3cf02d0bed0ead138d3ebd4ead6e6d825db85ddaedfe9e119e4fae5ece7e0e996eb66ed36efbef04df2c7f3dff4dcf5a0f6e3f6f5f6caf62ff67bf5b1f49ff398f29df173f060ef5eee2fed17ec25eb1bea3ee994e8cce71be78de6dae54be502e5b3e49ee4d5e4f5e438e5c2e53ee6f1e6f8e7e8e8ece90aebd5eb81ec25ed68ed8aeda1ed50edd5ec3aec2aebeee995e8e0e62ae585e3bbe120e0b7de44dd15dc25db3dda9cd929d9a9d846d8e9d76dd70bd7b9d672d667d692d6f4d6aad799d8c1d920db8cdc14deb1df39e1c9e251e496e5c3e6d1e791e854e92deaebead9ebfbecf9ed0def46f050f172f2dbf334f5b2f680f83dfa11fc46fe95002d036606f609e50d73124217351c7d21c426e62b0d31ef35623a823e1c421d45af47c5495d4b8c4c3c4d654d034d124ca84abd485746954358409f3c95380d340b2fd0293124421e5c185712500ca606310112fca9f7c8f385f031ee8beca4ebc1eb9aec31eeaaf09ef3fbf6d9fae2fe1a03a5072f0cb9105215a419b51d9b2117253428072b532d1d2f7130123108316330002ff92c6a2a3d278823671fd31aef15ec10ce0bb106ac01b2fcd4f737f3ddeee4ea6ce763e4c6e1acdf00decddc43dc59dc1eddb6defce0dde36be763eba1ef36f4e5f884fd3002af06db0ade0e9c1204164e19551ce51e1321a7227323b0235a236d222a21901f831d391bae18d815f2120210fb0c060a1a071f043b016cfeb3fb51f958f7cdf5e4f48bf4a2f448f56af6faf72bfae5fcffff89034b07180b180f36135c17bb1b28206a249f28982c273075336136bd38a03ae53b5d3c2e3c4b3bb539b0375035a932f82f372d612a9527b524b921ba1e911b3918cf1430117d0df80992067d030001eefe62fd95fc46fc81fc7dfddcfe9200cb0213055a07e409550cab0e3911a513d91524182a1ad51b721db21e791f0e202d20c91f3f1f721e691d7b1c8d1b921ab219b9188c173d16b114fe125711c70f750e790dbc0c4e0c230c1c0c4b0c9a0cdd0c240d5c0d6d0d8c0dcc0d2c0ee10edf0ff51028124c131b149514ac14371457131c127210820e6f0c340af307ce05a70378013fffcffc2dfa75f79ff4cdf12cefb4ec86eacae86ee787e62de63ae6b5e6a2e7cbe82ceac7eb67ed13efd5f08bf242f4fef5a2f73cf9dafa76fc27fee9ffa10140039a04a0055406a506aa067806fb0556059804a903b902d201c400baffadfe5cfdfafb94faf2f85ff705f6b7f4c0f33df3e9f2f1f25df3ddf38cf46df537f6faf6bdf74df8c6f844f9aaf90afa76facafa01fb1ffb08fbb8fa3dfa90f9aff8b0f797f665f52ff4f7f2acf14df0d5ee31ed63eb73e963e743e525e324e15edfebddf2dc87dca2dc51dd83de07e0d2e1c3e39be560e704e969eac6eb3aedc8eeb9f015f3adf59af8b0fba3fe820125044e06250896097f0a1c0b680b440bec0a570a67094b08f7064b0573036e012fffeffcbafa8ff8a2f6f0f465f319f2fcf0edef04ef46ee98ed17edd5ecb2ecbbec08ed81ed3aee55efb6f05ef250f446f620f8e1f956fb8dfcacfd93fe56ff0a007700a000960027006cff81fe4cfdf2fb76fa9bf887f649f4caf163ef3aed2ceb6de9f8e794e676e5a6e4fbe39ae378e363e370e39ce3d8e351e419e52be699e759e94feb57ed4def1ef199f2abf372f4d7f4d7f4bbf470f4e7f370f3f6f257f2e8f18df105f193f01ef060efa6eef8ed24ed87ec4eec4cecd0ec01ee9befb5f166f460f7b5fa9afee902b7073a0d38138d194f203c27202e0135953b8641c446204b7b4ef4509f528353b753475337527650004ed44acd46ea41643c4136ac2ff82819221e1b4e14980d1f073e01d4fbddf680f268ee8bea35e748e4f7e1abe039e0c1e08be246e5f6e8c7ed4bf36cf931000f07d90d9214be1a54208325022ae42d4a31da339035893683369d351534c631cc2e562b4827bc22ec1de418d213e20e140a6705cb0026fc75f7c1f229eee1e909e6bfe229e051de4add3ddd3bde3ae032e3ffe661eb33f053f58bfac5fff904f6099b0ee712a816c2194a1c2a1e611f2c2095209f207a200120061f9b1d991bea18cb154c12740e830a7c0653023afe3ffa6af6f8f2f8ef68ed5debc0e986e8d8e7b4e72ae86fe96deb0fee59f109f5e1f8e2fcd900a8047c084e0c0810ce138b17151b7f1eba219c2435277429252b542c012d052d6f2c5d2bc429bf2788253823db208a1e331cb5191d178a140b12c20fd10d100c550a9908b506ad04d5024b01170073ff4bff51ff85ffc5ffc2ff94ff4bffb9fe13fe7ffdc6fc09fc7afbecfa7cfa5afa45fa1dfae6f954f94bf8f5f64cf565f383f1b7ef0bee9fec6beb70eac3e971e985e912ea17eb75ecfded9fef4df1f6f2c5f4d6f60df971fbf2fd430063026a043906ef07aa09300b7d0c880d0e0e200ee20d410d720c940b750a150967072f05870291ff40fcc1f82bf567f1aeed3bea31e7eae488e3d6e2b4e2d7e2cce281e20ae269e1e8e0d6e046e156e206e421e681e8ffea62eda0efb9f186f30df56af697f7b4f8eef93ffba1fc00fe0effa2ff9bffc4fe3efd2ffb90f8aff5c3f2c0efeeec75ea2de85fe627e545e4ebe311e439e46de495e437e49ee30de366e22ee2c3e2e3e3c1e54ae8d7ea59edbdef90f102f339f4f0f460f5a9f58df54cf508f588f4f5f355f355f200f142efc5ecabe914e60ce20fde6eda27d773d44ad260d0d7ceb5cdc7cc3fcc25cc2bcc6ccce2cc55cd0dce35cfa8d0a1d21ed5b9d77bda4cdde1df79e233e5e2e7bbeaa5ed2bf05bf21bf42bf5ebf57af6b9f6fbf622f7dbf666f6a9f55ef4d4f2f5f080eee0eb36e985e65fe4e8e2eee19ae199e16ce120e1a2e0dddf45df0bdf24dfc8dfe5e03fe2ede3dbe5c8e7b5e975ebc1ecbeed9aee78efbef0a2f2fef4abf751fa71fce6fd98fe72fec4fdc6fc71fb13fad0f882f765f690f5caf43ef4f4f38ff31cf38bf287f142f0e8ee66ed1dec3aeb91ea4bea55ea5cea8aeadfea2cebb2eb6dec18edcded78eeecee56efcfef60f037f147f276f3bef4f1f5f7f6d5f77df8f8f841f940f906f994f8e9f742f7a3f6f4f54af56af41cf396f1d1efd7ed19eca2ea61e9b3e88fe8cfe8b9e92debc2ec75ee0cf036f138f247f368f4fef545f80ffb67fe49025806880aee0e6113f717ec1c2522a7278a2d91337e392b3f25440848a44ad04ba24b754a9f487a464c4428420b40d33d5a3b8d382b351031492cb9268e20441a0b14350e3b0901056d0183fec8fb0cf97df6e7f37ef1bfef90ee26eeddee58f08ff2bcf562f95bfdd0014306980a110f5a137217971b691fc822c9250b287e295e2a832a0c2a46291d289426c9248a22ce1fb71c4b19b0152512ce0ec90b2809df06d404df02d900b6fe73fc32fa3ff8c9f6e1f5a2f503f6d3f612f8c4f9bdfbeefd4b008502850469061b08b709960ba00db40fd911af13e914a415b8152c155e143e13b511fd0fe40d540bbe084106ff036a026a01b6004400b8ffdefe11fe8bfd99fda9fe9100f10280059c07f608cc093e0aab0aa60b210dec0e12114d1394154018371b3c1e3a21ae232825d325dd259f25b3252c26c0262c27e1267c254423af20571ef81cce1c971dd81ed61f11208f1f861e6e1dc21c841c981cdd1c031d191d631dd51d7c1e461fb01f881fdd1e8f1df21b711ae51860170a167b14b8121d11830f040ee60cc70b740af708f2067b041102cafff0fdecfc7afc71fccefc1bfd2bfd1efdbbfc1afc9afb4ffb8cfbcafc11ff5c028306e10ada0e0012ee13c31403153015d015291709190c1baf1c891d8a1ddd1cd51bce1ae319fb18eb176e166b140f12880f140ddb0ab5088b0667044902680017ff47febdfd36fd3afc7bfa28f8a5f573f31af2bbf10af2acf23af372f399f328f467f57df729fab2fc84fe68ff44ff59fe23fde5fbb7fa9cf97af851f752f6aff58ef5f3f5a3f643f782f738f76cf65ff584f425f44df4f2f4d0f587f60af76df7bff75df87ef9e5fa66fcbafd76fea6fe8ffe64fea3fe97ff1f012d036d0540076608b208ee0769069804c20250016600caff59ffc7feaefd09fcd3f9fdf6c6f36ff020ed43ea2fe8fee6c0e653e749e845e9efe9ffe976e995e8a6e703e7f2e686e7a1e80cea86ebe4ec1dee3bef5ef099f1e5f229f443f51cf6c4f65df71df83af99efa06fc2afd95fdf5fc78fb5cf901f707f5b4f30bf324f3c6f39ef4aef5c9f6b7f785f804f904f9c4f86af825f876f898f97bfb0bfed70049030c0511064d062806fa05b8059b057c053405e104870435040604db03950319033c02040183ffb1fda2fb6df91ef7e1f4fef2b8f13af18ef1a0f215f48cf5d5f6aff712f83df83df826f82af824f810f832f87ef810f92bfa8cfbfcfc6afe68ffd2ffc3ff0affc5fd30fc35fa0ef8f2f5c6f3bff1fbef4beedcecc5ebdbea3feaf6e9d8e9fee95eead3ea5febdeeb22ec33ec0aecabeb46eb10eb30ebaeeb8decb3edc9eeadef67f0c9f0faf057f1c6f142f2eaf24df31df37bf235f13cef08edc6ea87e8d8e604e6f4e5e6e6dde842ebe3edc5f084f34af6aef9a4fd3e02d107e70d1d148f1ad220a926642cda31fb36173c02419745d649654dff4f7b519a5179504c4e2e4b8b478043f93e173a9334592ecd27ff203f1a1114490ee308f20305ff36fad4f5baf145eebaebcae9b9e8a6e850e919eb07ee9af1e8f5adfa56ff2b043609390e9e135419ce1e0f24d828ac2caf2ff0313633a3333233a6311f2fcf2bca275023981ea21974141e0fa309310404ff39faf7f53ff2e1eee0eb3ee900e778e5c7e4d9e4c5e528e76ee89ee9a1ea6bebaaecb8ee88f15ef5eef986fef002c5069409860bb30c2e0d6b0dad0dff0d6c0ea90e550e230dcc0a5407ee02e7fdc0f8daf379efe5eb13e9dce623e5a3e33ee204e10fe098dfc5dfaee055e263e4b1e655e900ecb1eec2f1e5f400f861fba9feb801e504d5075a0aa30c5f0e800f4010d710721149127213851439153a155114ae12d6104e0f5e0e2c0e760ea80e940e3b0ea30d5c0ddc0dfb0ea810b1127614d6150517f217c618bb19851adf1ad01a571a8a19c9184518b917da1666150113c10f340ca6085d059802eeffe4fc5ff931f58cf023ec5ce880e5d8e323e300e33ae37ce3ade307e4bae404e619e8edea57ee1ff208f6ebf9b4fd690105056d08a70ba80e5611d9132f162b18e519451b121c8b1ccd1cb81c8f1c391c3e1ba0194217de13db0f9f0b3f073803c4ff8cfc82f991f658f3f9efd1ecf4e9aae73ee684e55be5dae5cde616e8c4e988ebf7eceded41eefaed9feda1ed2fee61efe8f02ef2d7f2c8f21bf23cf19ef071f09ef0f9f01af189f021ef07ed6feaa1e709e5e4e249e17be07ae000e1fee12ae30ee4b0e429e577e514e651e7ffe823eb7fed79ef02f12ef2fdf2eff35df51ff733f947fbc4fca0fde2fd86fdf7fc54fc61fb28fa7ff82df692f3f4f06aee5eecdbea9de9bde823e884e7fee687e6e0e529e576e4ade303e3a1e26fe28de211e3d4e3c2e4c6e597e614e747e753e795e769e8e1e9dcebe9ed70ef1bf0c2ef87eef8ec81eb5eead7e9c0e9b8e9bce9a0e939e9eae8d4e8d6e838e9e6e979ea1aebc1eb1cec6cecb8ecb3eca6ecc5ec0eedfeedd6ef56f261f58cf82bfb0cfd24fe7efe8afe8ffe8efe8ffe54fe94fd48fc5efae0f712f512f20bef5bec2deaa1e8dde7aae7abe7b0e77fe709e79ee681e6c9e68ce79ae88ae931ea87ea86ea7feac8ea77ebb4ec94eee6f09bf3adf6ddf91cfd5f005d03fd0517084c098709c208f1068304e70157ff40fda8fb29faa1f8bff627f421f1e8ed97eaafe74ee53be39fe163e058dfd1dee5de69df74e0c6e1fae21ce438e567e604e81bea76ecd2eecdf036f229f3def3b0f4c2f5eaf60af8dff841f984f9d8f944faf2fa87fb80fbe9fabaf90ef891f67cf59ef40df46cf342f2daf078ef4eee11eefceebbf035f3fff579f8bcfa06fd7fffc9023c079a0cbe124919971f92254b2bbd303236be3b0541cd45bf497b4c234ef24e114fd94e494e134d1d4b33484844d73f363bac36a032e32e1e2b4527ff22381e5d198014d40fca0b2e08f6046f02660001ffc0fe63ffda0047030506e3082c0c850f04130217e41a651ea7212424f825bd274229a22a312c742d4c2e002f342fd62e162e922c3a2a6a272c24ce20bc1dd61af717fe148d11a80d9809a1054f020700c9fe91fe12ffcbffa0009301a2022d045b06db08600b920dfe0ebc0f2d1075100011111239133014e7140b15d314d414121589152b1638162315f3129e0f910bb7076e04e801530038ff2ffe35fd19fcfafa48fa11fa6afa74fbd8fc65fe1c00c9018803ad052808fe0a2d0e3e11f1134e163418d419891b421de51e6b207a21de21b321eb20831fab1d661bb418d9150c1378106a0eff0c1e0cb20b850b520b060ba70a5c0a6d0a0c0b4d0c1c0e29103e1241141616e417d919c31b8e1d291f4020f22090210e2291222f236a230b231d225e20f81d4b1b3318bd141611010d97082b04b3ff60fb7bf7e4f3c0f048ee60ec26ebaaeaa3ea0bebe7eb08ed98eeaef012f3c0f5a8f88cfb95fef601a505b509030e02126015f5179c198f1a321bbb1b441cc21cf11c8d1c851bfb1927185016bb1463131312b110140f140de50aac0856060404c80177ff42fd72fbf6f9e0f845f8ccf756f725f742f7e0f75ef98cfbfbfd66004c024c0393035203a602de010301d3ff3bfe38fcc8f931f7d4f4dff26ff17ff0d4ef1fef35eeffec7debd7e947e8dee69de593e4b1e303e3dfe297e358e543e805ece6ef50f3cbf52bf7f3f7d4f84cfab3fcd3ffee027105ec063507c2061d0694057b05b405cb059105cc0441032f01bdfedafbd5f8d4f5d0f233f047eef4ec61ec66ec70ec58ec0bec5aeb9dea2beaf8e922eaafea50eb07ecececd0edb4ee94ef29f05cf046f0e4ef5befdcee61eee4ed5fedafeccdebc6ea9de975e869e779e6b2e508e55be4c0e34be3fbe206e36ae3dee349e482e455e40ee404e459e45de50de7f0e8ccea57ec42edd7ed6aee21ef5af010f2d3f381f5d8f69cf72cf8c0f852f918fac9fae3fa69fa48f98cf7d7f57ef48af338f33df31bf3c7f20ff2d6f08fef6fee87ed2aed48eda0ed43ee13efe1efd0f0d8f1c3f295f338f483f496f496f498f4cef44cf5e9f585f6edf6e6f679f6d1f50ff576f420f4daf38df318f34cf25af17bf0a7ef06ef92eefced59edc9ec49ec3becd2eccfed32efb2f0c2f160f281f2f9f13df18df0d4ef77ef82efa4ef0cf0abf02af1bdf165f2daf243f391f36af3e0f2fbf1b3f063ef58eea2ed4ced1eedbbeceaeb94eae0e814e76ce523e428e344e26ae173e042df1ade0edd05dc26db56da4fd946d86dd7ced6e4d6f5d7c1d93cdc4cdf7ae2c8e571e94fed65f1d3f544fa99fe1d03cf07ca0c54122518e11d6f237b28e12ce4308234b037983a073dd03e02406140bf3f233e663b913707330f2e02294024cc1f8b1b5417e212290e38092b044effd0fae0f6d3f3c4f1d4f035f197f29df40af74df939fb1ffd0aff4d015704d407840b520fa012421588174419a01a121c6c1daa1e0a203621fd2179226322ac219b20401fcc1d831c601b4b1a1e199c17b4156213c710390ee90bfa09a708dd0775076c0783077a075107f3066b0621065f0649070c096b0bce0dc10fdb10d410e90f8a0ef90c7d0b260a92087d06e903d6009afdcdfaa9f837f769f6c6f5d5f476f392f164ef7eed43ecffebd0ec52ee0ef0acf1d0f28ef34bf42cf55bf6ddf742f94cfa22fbdcfbdafc9dfe0501a003fe057807b80721074606b80507062d07800855091c097b07d6040602bdff84fe93fe74ff9300a4017602380380049e0695093e0d08114414a61632182e192b1aac1bd01d5220b6226b24fb24662405232221111f0f1de11a58188f158312680fa60c2b0abc072905fc010efebaf95af584f1ceee37ed99ecb4ecf7ec35ed97ed13eeddee2cf0b8f175f381f5bcf752fa85fd1c01db049f080f0c090fbc114214a716ff181b1ba51c701d6b1d801cd01aae184316bd138311bb0f640ebb0da50dba0de10dd60d2f0d170ccd0a5a0921086e070f07fb063c078607c7072c089608e60831094c09f4082e0804076b05a9030f02a20073ff7bfe5dfde6fb1ffa03f8c7f5c1f3e9f121f049ee19ec90e90be7ebe4aee3ade3c2e477e633e85be9b2e96be90ee946e983eadaec0af088f3e4f6ecf993fc13ff990106043d0609082209a309c2099c09820985096a093409c508db07aa063f0575039801c2ffccfd00fc75fae6f86ef70af669f4aef2f8f029ef7ded2eec2deba9eac5ea54eb3bec4aed21ee91ee93ee39eecbed9cedcded5bee15efa9efd6ef8aefdeee0dee4beda6ec0cec44eb19ea8ee8d0e62be50ce4aae3fae3e6e420e641e73ce80be995e91ceac8ea7eeb6eecb0ed10efacf08af25df428f6d8f722f91dfadafa44fba4fb1dfc8efc19fda3fde3fdfcfdeefdadfd95fdaefdb8fdb4fd47fd01fc05fa7cf7a0f417f22bf0c6eeeced4feda2ec19ecf1eb57ec88ed5cef54f111f34cf4f1f458f5ddf5aaf6c4f7f5f8def949fa37facff94cf9e1f894f84ef8e7f749f788f6c7f526f5c6f491f450f4f3f36ff3c1f225f2b2f132f192f09eef17ee41ec88ea39e9e0e8c1e98feb09eeacf0c2f20df476f406f442f385f2e0f184f149f1e4f082f041f033f0a6f06ff116f261f2fff1def085ef6beef3ed65ee81efccf0e2f15af23ef2eef1c1f114f2f0f2e4f38cf47ef47ff3fef175f033efa5eea7eebdeedaeeceee77ee41ee3fee3bee71eed8ee49ef45f0fcf13bf42af78bfacafdec00f203b5068f09ad0cd70f191353162a19b81b191e41207822db243827a4291f2c8d2e2831f833bb365239623b7a3ca23cef3b843ad838133720351233a830ac2d642aef269923fe202a1ff41d421d581cb91a9b180d16951332120512f612f91432171419cd1a221c401db01e0820fd20a4217a219d20e01f681f871fa6201b22582345246324d5234923cb228922b122b6225622b1219520421f1b1ef51cd51bb61a2f194d174315ff12dc102a0fcb0de60c8f0c7b0cb50c470dde0d7b0e240f8b0fcc0f20106b10dc109411351292129912e2116c108d0e4b0cf7092208d3061106fb051006dc0550051f044f027100bafe58fdaefc89fcaffc39fde0fd72fe1bffacff0f008b001601b401aa02c103cd04f4050e071c0882093a0b270d480f36119212601394134b13ef129e124f121d12e911a01179119411fc11bd12a5136114c914d514a4148814ce149315bf160a181c19b219b7195c19f318c3180a19c619a31a551b921b091bcc191e181a1604141d124210790ede0c3d0b9309fe07440658045f023a000afe17fc5efa04f945f8f2f7f5f740f85ff814f867f752f631f59af4cbf4f7f519f8b0fa4efda8ff7701c302c303940459052106d8067607ef074908a20808098e09370abf0af20aa00a8b09de07f8052004c8022d02040213021702a601da00070045ffd3fecbfeccfe9dfe37fe79fd96fce4fb5ffbf3fa7ffaacf962f8cff624f5b6f3d8f28af2b8f245f3f4f39cf427f570f560f5edf402f4bbf252f1f7eff4ee86eeabee4fef40f021f1c5f11df223f20ff209f2f5f1c5f156f175f05fef7fee1feeaaee33f032f22bf493f5d5f507f594f3cdf160f0c2efd9efacf01ff2bdf37df556f7e4f819fad8fac5fa13fa2af93ef8d6f733f8e2f885f995f976f84ef6a3f3e9f0e4ee00eeefed6cee0fef51ef4bef43ef48efa5ef4cf0aff098f0f2efa1ee29ed17ec7ceb6beba5eb79eba4ea25e9f9e6a6e4aae214e111e0a2df79dfaadf55e05de1e5e2d7e4ade623e8e2e88de86de7f2e56be47fe36ce3dae3a1e45fe59ae593e598e5c7e595e6f3e746e94aea9aeadae989e824e7f0e581e5d0e545e6b3e6c8e637e681e516e512e5c5e5fce619e8f4e86be96ee990e939ea67eb2fed3feff6f01ff2a0f274f20ff2c2f1a1f1cff11cf232f209f29cf1f6f071f032f01df02cf019f098efc5eebdeda7ecddeb64eb03ebb1ea47eab3e95ee9a6e9afeaacec58ef0ff267f4fff5a4f6c4f6dff648f761f814fae8fb91fdbdfe36ff46ff20ffc7fe65fedbfdebfcc7fb98fa7bf9ccf87cf82ef8bff7e2f65df58df3c4f129f01bef9fee6aee74eeaceef6ee92efacf02df20ff415f6d2f715f9cef9fef9e7f9c9f9bbf9bef9b3f96af9caf8d3f7b4f6b6f510f5ecf456f519f6f8f6bcf729f82cf8d6f728f73bf62af5f2f3a0f25df13ff076ef3cefa5efc2f08ef2cdf445f7b8f9e2fbb3fd3fff9f000f02ae0361051707a708cf09990a290b8e0b030cab0c620d150e9f0ec00e870e220eb70d9e0d090ed40ecf0fa910f7109810980f140e530c7d0a9d08c706f80453033202d1015e02f30331069e08d00a490cef0c130df00ce90c5e0d240ef70eb00fee0fa30f320fd00ec60e660f7910a511bb125a135e13041365129911cd10db0fab0e660d2b0c3f0b030b870bb00c4c0ef80f7811bb12b51385144b15f31584160817561777177f174417da166816dd155e151915e114ac148b143d14c4135713cd122f12b8114111ca10811027108a0fac0e400d430b1b09ef060a05db03460322036c03d2033304c2047b0583062908530ae70ccf0f80129414e9154816ec156e1516153215f81508170c18ee187a19bd19ff19291a111aa1199918fe1628154f13a0112a10ae0e050d430b99096b08f9072208a6082d096d098f09e309870a910bc50c9b0ddb0d820d9d0c7f0b570a030996073406fc045f04b104bd0533079b084a090509e5070f06f2030302700067fff1febffe8afe1cfe49fd53fcaafb9ffb5cfc91fd80fe82fe3bfdd2fa21f826f68ef599f6cff84ffb70fde1febeff86008b01bd02c3031a0482033a02d900150062009e014703ab0426058204e902b50066fe58fcbbfaacf914f9c7f8c4f80af9a6f9cbfa7cfc71fe4b0099010f02d2014101be00870081005100c5fffefe68fe8cfeb2ffa501b803240574059a04fa023701b9ff8dfe98fda4fc97fbaefa48fa9dfabbfb5afdf4fe1b00a200970052002e003d005300210044ffa2fd91fba3f976f89df839fae3fcfcffc5028a041605ae04cc031103ef024903be03e30361035d026c011601a101ed026204510556056f04f3024901a3fff9fd17fcd7f95ef713f567f3b5f20cf31cf466f56ef6cff66ff675f528f4e0f2e7f15cf14df1c3f1bef247f45ff6d9f85bfb7afdd7fe44ffdefef9fdf4fc0bfc4efbacfaf9f922f93cf866f7bdf665f651f64ef634f6d9f524f544f475f3e4f2c7f20df375f3f1f384f43df56ef639f84ffa46fc87fd8afd4bfc1efa93f76cf526f4def387f4caf53ef7b5f810fa4ffb9cfce9fd0bffe0ff2000b2ffe0feeafd13fdaafc9dfcaefcccfce4fcf6fc2dfd88fddcfdf7fd99fdb0fc61fbe2f97af864f7aef64df633f63ff659f679f6a1f6d8f62ff7b7f765f81ef9bff923fa27facaf927f970f8e5f7cbf752f876f9ecfa50fc31fd45fdb0fce3fb57fb7afb4efc58fd14fe22fe69fd68fcdbfb43fcd9fd5100ed02f204d6056d0505040f02e7ffd2fdbcfb61f9bbf6ebf34ef190ef39ef68f0dbf2ddf593f85bfa0bfb0efb29fb19fc45fe6d01b1041007bf078806050437010aff04feeefd10febcfd8efcb1fad9f8a6f763f7faf7e1f88ff9daf9e1f913faf3fa9dfce7fe880108041c06df076909d00a380c840d790e0f0f3b0f010f960e080e4a0d740c8b0b8b0aa409f1085f080a08060860085909150b750d4e103c13d215ec1773196c1a0b1b491b0c1b661a371970174215ac12d30f3e0d3e0b360a950a140c1b0e271067117811bd10900f6b0eea0df60d400eb30e190f900f96104f12ba149917191a9b1be51bce1abe18711645149a12c1118e11e111a81279132114a514f8145b15261640176d184b1945191f1811166d13af10380e040cff09130825065c04f202fc01a001f901f7028c0484066408c5094e0ac6097908e70666055804d5037a03090360023f01d1ff7efe63fdcdfc19fd2efef7ff5602bd04b306f20719082f07a605cd031c0209018600640076005f0004008afffdfe8afe5afe5afea2fe6effd80013033106d809900ddd1035135f147e14ca13a012691154106b0f9a0ea10d3f0c4f0aca07d404c201f3fec8fc98fb8ffba9fcb9fe62013704e9064a09420bd60c020e9a0e740e8a0dfe0b1d0a3d088506d904f2029800cefde6fa6af8d1f643f6adf6caf73cf9ccfa6dfc0bfe9dff2001920203047d05e70602086c08cd071c06ab030901c5fe22fdfafbe9fa83f9a5f78bf59df352f2e0f131f22ff3bbf4b4f627f9f4fbacfe0501ca02de0398044105aa058c058204390221ff15fcccf9bdf892f853f877f7fff57ff430f4bbf598f8b8fbc8fdd5fd53fc80fa61f99df9d2fab9fb72fbdef972f74af54cf478f455f52df646f67bf5fbf3d9f132ef0aec60e8a1e477e165dfdadec7df97e1d4e326e638e807ea7feb47ec4aecb3ebe5eab3eaa9eb99edfbefd3f122f2eff0d4ee91ec22ebdcea3febfaebc7ec68ed31ee3eef1ff09df07cf097ef89eed7ed83ed99edc3ed84ed2ded28ed9cedbdee21f0e8f0cff0e1ef56eee5ecccebaaea46e975e74de599e3fce26fe392e47ee541e5c8e396e179df6bdebcde05e0cde17de3b5e4ace59fe695e7a6e8afe96cead4eac2eaffe998e89de667e4d4e284e28ce3abe5e3e7fbe8a0e833e78de5f4e4fae524e8aceaaaeca8ed41ee51ef57f17df412f802fbe2fcb6fddcfd1bfeb1fe3cff68ffcbfe37fd2cfb23f95cf734f6aef5a8f543f65af782f86bf99ef9d5f879f714f61af5f6f479f50cf667f675f64cf65ef6cff632f713f711f60ef4a1f1afefcfee34ef80f0e3f1ccf218f310f375f3e6f473f7e3fa94fe9f0188032b04920327025e0065fe6afc68fa31f8ccf538f37ff0f8ede9eb89ea3cea0feba9ecb7eea7f0dcf146f20cf25af185f08fef3bee8aecb5ea42e9fbe84beafcec5cf05df33bf5f5f50ef66cf6ccf71dfab6fcb4fe3eff18fec2fbfff89af618f583f4b6f486f5cff697f8bbfad2fc77fe4eff2fff7efed1fd8efdf6fdecfe0d002d013a021d03e103620464041904f3036704d7050a081f0a470b130bd709c5080509100ba80eb212f215f817e01824197319d519ef19ca19a619231a341cf71f9024c428072b652a36275322da1cf8171a14601120105610e511af14db17871a811cd31d171f30211124f426e228b92842267f22951e9d1b281aa4195c192319f3186019131ba81d3e2005221f2295205f1e451ce31a711a6f1a811aa71aca1a101b6f1b3f1b2f1a76185916aa1424146314b2146e140113dd10360fc50ec00fab1132137b13a8125b11b21071112913ee14cc1508150413c610ef0eec0db10d860d280df20c210d1a0ef70ff011321358134b12b910a80f910f87100012d2124e125f10340dbf0919079e05650538063d07dc07ee0756078a065a064707b109890ddf119315a81764172115fe11ef0ea30c110b36094b0673028cfe4cfc4efdb8016108510f4e143916841576138611a910ae10af10bf0f540dcf094306d7037d0371050109110d6a10fa118211880fc80c2a0a64087c0736075507a207480892096a0b770dff0edf0e7c0c1a089d029dfdbafa8afa8efc6cff61016401acff54fde4fb5ffc8dfe5d017a03f6030203a201ed0094016a037f05d906d00671058303f7016e011302670370044c049f02d6fffefc4afb96fbc9fdcc004d035404b30350027001c4012f03bc0409055403e3ffc1fb58f8a8f6d4f65af865fa40fcc7fd37ffce00af02b40467064d0702074c053a020bfe27f93ef411f033ed03ec6cecd5ed8cef12f138f26af35cf571f891fc1701df04f206e906fe040e0229ff1dfd77fc53fd45ffb201ce03c30431042a022bff0efc4df9c2f614f4c8f0c8ecf2e86be60be625e80cec82f0aff435f82dfb04feaa0089021f032202d9ff49fd3bfbcef9b4f841f7f4f424f2a8ef47ee52ee55ef6cf0eaf0b2f03ff052f046f1e4f2a7f412f61ef746f8f3f900fcb2fdf4fd06fc35f8c2f336f09feeedeefaef6ef082ef66ed31eb04ea62ea2cecc5ee96f185f48ef765fa8ffc66fda6fc07fbcff914fa22fc03ff120139017cff11fdc2fb6ffc8dfeb60060010b00d9fd7efc1bfda9ff9302b003ef01c2fdd7f874f5fef436f7d4fa41fe560007010401ea00f200d000e7fff5fd34fb1bf84ff542f308f2aef134f25ff3c8f4d3f5c8f57ef484f2d9f092f004f25df443f68af6fcf4d5f2f5f1a6f3fdf780fdca0125033f0125fddcf80ef614f55ef5cef56ff559f452f312f30ff409f623f8b9f99dfafdfa64fb32fc45fd4dfee5fed0fe3cfe6afd80fc9dfb96fa28f955f71cf56af25fef11eca8e8b0e5d0e377e3cfe479e7aceac4ed6ff0d8f280f5a8f811fc09ff9f00510089fe48fcccfaeafa50fcdcfd4ffee2fceff9def61ff56cf578f7fef9b3fb29fce9fb22fcd2fdf00089045f078d0824080207080695055f05c6047903c2015300ccff10004f009dff64fdcff9f6f504f390f1b0f1ebf28ff46ff6d1f8fdfb1100b004ef08e60b010d3e0c450afe073b06a30553060008540ace0ce10e5b1033118411ba112a12de12ad131f14b01348121f10ab0d860bdd0990088507af0667065507b609340dfe10d713f2148614601384128b12e9125a12b90fa00a11040efe6bfa2cfaf0fcec004304f205ec05430575053907620a1f0e4b11471336148614b214d4145b14ba12e30f3c0ccb08b9066b067b0717093f0a730a110ae2099a0a7a0c130f9f117613411415143513a7114c0f0e0c12080304df005fffdaff0b0209050408890a510c5e0db00dec0cd00a790752033fff2cfc66fabbf997f94ff9dbf8c5f889f971fb2efea100bf01340164ff5ffd69fc23fd5aff3802b8044506f00649071e08ef098d0c460f1e1128111f0f950ba70797045503fd03e5051908e9093b0b830c550edb108d13381596140111bd0a0503bafba9f6dcf447f6b8f954fd61fffcfe86fc84f9bcf73df8c4fad0fd6fff63fee8fa96f66ff3cbf2acf4c9f78afa26fcedfce7fd170092034c07cb09250a90082e065304b903080423040f03a30084fdb7fa02f97ef8c1f864f96ffa3efc09ff7c02b0058f07a407790623058d04d004f304a703520081fbb6f681f356f256f213f289f001ee3aec42ed15f212fa3d032e0b4f106f124f12e610c30efd0b9708ed04bf01c2ff14ff2eff57ff2dfff8fe8dff5f01db039005db04e6007cfa9ef36dee2eec8ceceaedcceebcee66ee5fefe3f2bdf871fff6049a07060751041f01d1fecbfd4bfd0ffc26f973f4edee2eeab8e774e84cec33f28ef8a6fd3b00020088fdfef9e4f60ff53df495f3eff180eee8e9e0e522e4cae57fea3df0aef45ef65ff582f333f3e1f55ffbbd0121069c060603defce0f668f311f3d0f470f6a2f59bf15deb1ee56ee1aee144e544ea38ee5befcced1aeb3ce9bbe9a8ec81f06bf3eff39cf16eedfee89ee51fe46ce4a4e5eee6bae7d8e7c7e74de8f8e9f8eccbf062f4c2f65ef768f6e9f4e0f3c3f380f454f56ff5e3f464f4c2f49cf69af95dfc70fdeafbe4f7b1f200ee0aeb5eea86eb80edaceff1f18ff413f895fc6d01990518086908ea066804a401f0fee4fbe7f7f1f2abed73e9e4e7b6e960ee73f40ffad6fd92ffdeffafffcaff30005300b9ff3efe33fc64fa9ef945fa5dfca0ff90039f073d0bc90dc20e000ecf0be2080706c30314029e0011ff92fdc3fc55fd75ff6d02c604fe04660299fd3ff83ef4e4f269f4edf718fcbcff1a02fb028f0235017bff25feecfd2cffb101ab04f406af07ca060d059b035a036704fc05fb06aa0619052803f501fc01cb024b0358028dffc1fb8af857f7a2f89dfb87fe9fff1afe8ffa8bf6def3cdf364f697fae9fee20193020c0130fe40fb86f9ccf9e7fbf0feb1012d035903150371030c058707430962081b0413fd68f5fdefbaee8bf1baf69afbd0fdd3fc03fab2f712f8fbfb6002f2083f0de70d4f0b2d07ae0367027f03ed055808cd09730a650bb20dc71122172a1c231f1b1ff41b89166d10ff0a1207d304ab03b802580148ff15fddafb53fcbffeab02a7065509510aee0926094809c00ae90cb10e090fb30d950bfd09110a2d0c480fdc11dd12d611690f120dcb0bca0bd20c2e0e8b0f7f11b9149019a61f72252429be292c278022631dc918d5142c113e0d3a091d06ce04d505dd087e0c810f7f11871242134e14481568153314b511ef0e4d0d8b0d8d0f55125d14e314121453124810400eba0b6908c4049401e4ff85002303b106300a140dad0fbd128116701a421d6c1d611aea147f0ece08d5045a02ab005cff6cfe76fef8ff7602d604f3053e0577034702f902d605d109f80cd40d210cc608640537037c02dc02c203b404d4055007b30838092a083805070110fdc9faeffa32fd7900a2030906bf075409180bbf0c9c0d070ddd0ad6072605c403fd035e05ea06bf078e078f0643051c043403630274014900edfe92fd65fc81fbedfaabfabcfa0ffb8cfb3cfc26fd49feb2ff3e018d02450328032a02a20014ffd8fd08fd7ffce8fb1bfb56fa2bfa39fbbafd29014d04bf057f04a30095fb76f70ef615f8d3fc58028f065408bd07d205f503f902db0227037603c1036a04c1058107cf089b0843062a029dfd40fa5df943fb0dff1403b105c405110354fedcf80af4e2f0bdef5bf025f268f4a9f6bef887fad0fb70fc49fc7afb75fab6f971f95ef9d6f852f7cef4eef1deefa1ef7bf103f55df98dfd0b01bb039b05a4069f065405f9020b0027fd01fbf8f9e5f994fad0fb45fda6fe91ff87ff4cfe0dfc54f9e4f624f5edf3e0f29ef13af09cefc2f0e9f376f8d9fc15ff1afe38fabdf477efb2eb8ae978e8fbe7f0e7fbe8feeb0ef152f746fd5b01ee02920293013801d1018b023a02fcffe0fb43f7cef37ff27df3e9f561f812fae4fa12fbdefa0afa02f89af444f041ec59ea7aeb3bef6cf46af9ebfce7fe00009900910025ff7dfbc6f559ef32eafde7eee899ebeeed4eee88ec29ea55e983ebd7f0f1f7abfe5d033f0586043f0272ffe0fc3efbd0fa45fb13fc6bfc80fb48f986f66af40af476f5b1f771f9acf957f8bdf64af693f73efaf7fc3cfeb3fd3dfc47fb03fc6ffe39018c020701a6fcd6f67df138eed4ede7ef5df348f7e4faa9fd52ff9fff7afe47fcc6f9cdf7f4f61ff7aef7faf7c9f7a2f782f81afb4fff0f0498077a084c06b20131fc6af715f4f9f152f028ee31eb4ee8e0e627e8c2ec0af43afc4c03b007ea08c507b3052a04040400053606d1068906020687061b09cb0d78132918281ae21815156710420ce4087905c4001efa57f272eb80e795e712eb03f052f4c5f694f721f8aff984fcd5ff1102e7015bffb7fbdbf861f897fa56fed201860301034401fcff82002e030907660af50b5a0b5d09a2079e07e309030eaa124016be17e3164b144611130f530eed0ef70f2710a90e780b800734049302b302bc0338042503b100eafd4ffcfdfcd1ffbe0391074d0acf0bb70c830d650e500fe60f0c100210c60f220fc20d1e0b47074b037b00f3ff160211066b0ae60dfe0f28115212fb13db15ed160316c7120d0e5f0977063306fe07720a160c070c9b0af8082308ad08650a5e0ccf0d6a0e110ef40c5f0b6f096607bd05d9040f05520602089609ce0a930b330cfb0cae0dea0d620df80b1b0a7c08590790069c05b803a200dbfc42f9ebf68af60bf8d2fa11fe1901b2030d069408a10b0b0f4012921420154d13450fc309e0030fff7afc87fce8fe9a023d06bf08b3096909c808ab086e09b80a850bb90ad30704031ffd55f77af2b0eec8eb89e9fde7bee79ce9feedaff4b5fc81049d0a2f0e110fd60d820b1a094007f405cb044a032601a0fea3fc20fc81fd7300e80383067407dc069e05cb0410055a06dc07aa087f08ba07f606dd068f074208da0793054401aafb3df68df29cf16df314f721fb2efe71ff17ffeffddffc83fccdfc0afd6efc94faaff797f470f219f2ccf315f707fbb0fe7f016f03d80413062707bb0742077805c7020f004afe3bfecafff801a5030d04f902ff0026ff2efe61fe97ff4c01fb023604ad0456044703ca017500b5ff7fff84ff1cff8bfdc3fa49f7c8f3d2f086ee76ec34eac5e7bfe50ee551e673e9b0edd3f1e2f4a6f67bf709f8ddf8ebf9abfa80fa01f95ef670f32ef15cf038f110f3bbf45ff59bf4ddf272f189f16ef3aaf6fbf9d7fb91fb81f9aff679f4d6f3d4f4e6f62ff9e5fad4fb29fc4bfcd4fc1afe00002102a2037303f10015fc8df5c7ee1fe94be554e398e258e279e287e346e632ebedf136f990ffea032a061c07aa07440892087907ee03ddfd52f642efd3ea52eaa6ed64f350f964fd99fe10fd03fa32f7e4f597f62af9ccfc8a00fa0300078209790ba00c5e0c520aaa061602b4fd9afa66f905faa6fb3afd0efebffd61fc87fab7f825f7f5f519f548f45ef34df21ff134f01ff066f161f4def804fecf027506b308f9091c0ba60c620e6d0faa0e540b780511feabf6abf0e7ecb0ebc9ec9aef7df3c5f7a8fb81fef3fff7ffe9fe41fd5efb8af9f6f7d8f6b1f6f9f7b2fa62fe100285041005d903ab0188ff0bfe0efde5fbcef995f6d8f285ef53ed9bec17ed47ee1bf0eef212f762fce9011f06c20785066e035400aafec5fed1ff3100acfe4ffb35f7baf3d2f17cf1f9f1a4f278f3f7f4a0f73dfbb0fe8900fcff86fdd2fac9f976fb4fff85032c06570681043a02100174019002f4026501aefdbef807f4b6f04defa7ef4df1baf384f64ef9a7fb3ffd58fea4ffe601af05bd0adf0fdb130916971676167c168f16be15c9120a0d5b05b5fd3af849f6aaf7befa9cfdedfe70fefefcc7fbbbfb51fd5600450496089b0cab0f65119b118010a70e730c0c0a6a074504b8008dfd9ffb89fb6bfd63001603b0040805a0046c04ea04d705b4063007a7072f09b70c38127818481dc01e651c4e17ca113c0ea20d670f0f12dc13fd13fe12dd117511161201131a13c611f80e5f0b2b0825068b050d06ba06b606b505e4033102e20192033007e80b08102612e711ac0f980c130abe087808cc08180927094709b709950abd0ba70cfc0cde0c890c750c1b0d720e3d103712e5130115ac1509166b165117b418251a071b7b1af817c813b20ec009f105a2039f026c0272026e025f0246025402b30254035504e105d707340af70cd60faa123d15fb168417b1168114ac11430fd20d860dfa0dee0d460cb4088803d3fd12f943f69ff5a7f653f8c0f9adfa88fb4efddf005106d70cfc123017ac18ad173715ae12f9102110c40f4d0f3f0ec90c710b830a280a3c0a0c0ad208040653010ffb4bf48aee56eb9deb47ef52f51efc1e0285061409cf09ec087f06a60221fe24faeef75ef84dfb97ffe4032d071709240af00a8e0b8d0b400a28076802d5fc9bf7bff3d3f110f251f412f8acfc4201d104a0068506d8046102d3ff6ffd2afbb9f8e7f52af354f1edf038f2eef4fcf74ffa74fb5afb62fa52f9a5f84df815f8baf707f721f682f5a3f5d7f644f9b7fc940003041f0613068603e2fe1cf961f3aeee37eb67e88fe55ae234df60dd26def2e105e8b0ee4bf452f878fb45ff1505a00cf2139f18d3187d14c60d9007cf03be02ae022201a2fc85f5b2edabe70ae5e1e534e98fedebf137f69cfaf6fef60222060a08e1082109bd082807bc032ffe51f72bf1e8ed8eee6af24af7a1fa1dfb6df996f784f7cff94cfdcbffb8ff2cfdb8f955f713f72ef8bef838f76cf3c1ee90eb8aebc6ee08f482f9fbfd580104044a061108ab089c076b051f039e013e013c014600e5fdd0fa8af8bef8dffb81006304b105ee0371007cfd9ffcf2fd2c00880116014fff8bfdfcfcc3fdc8fe94fe4ffc68f865f4bef1dff01df105f156ef16ec61e89be5e3e45be627e95eec81ef7af28ff5daf8fbfb89fe5900b80184036206240aef0d6e107510e30d7c0961048eff2efbaaf66cf158eb11e5f9df4edd88dd52e096e425e975ed94f1e2f5c1faf8ff970494072208ff05b20139fc98f6aef10ceef6eb76eb56ec23ee3ef007f243f339f46ef57bf7b5faa4fe5302ed04dc0526059c0317021201b0007b00b7ff1efed9fb79f9f2f7e5f73ef981fbd5fd64ff13006300f4003f022704dc056e066105fe02500094fe91fe3f00cb020305fe058105eb03df01f5ff5dfec2fca6fabcf7f9f3afef78ebe6e761e545e4c6e405e716ebbcf04af7d6fd5f031807c208a1082907d9040f02f4fec3fbf7f813f781f668f77bf93efc5effc0028306c90a330fe912f9149814ab11250d6d08c104df029302cc026c02f10093fe32fcd7faf9fa23fc4afd64fd09fcbef9b6f729f79ef88dfbaffebe00f4005effe4fca3fa2ff979f8f7f7d9f6b0f4e7f18eef04ef6af1ecf683fe4306f60bfc0d0f0c4a07a8013afd2bfb56fb93fc5ffdadfc89fa1bf805f7b8f89afdb2040e0c84118a130f126b0e930a3108d3079508dc086f072d04290008fd0efc5efde4ff30025a034203a20286026303ee0491069a07ae07080717063305a1047f04eb04020694071b09e609450922074604f8016d0113032e065509360b4b0b500aac095e0a680cbe0ec40f7e0e550bb007220582044e052606e10551046f02980172026904fa05a705230390ffb3fcfafb9dfd7a001f03e3042106fd075e0bd20fb3131315ac12da0c8405f1fecffa82f91dfa48fb10fc1afcbefb97fbeafbc7fc28feedff1e02de0409084f0b5a0eda10a612c5134d14451491130d12af0f770c7e081904b3ffbbfbbff836f741f79bf8b2fad8fc8afeb6ffc4004b0291046207120aaa0b780b8d0992066e0304019effbefeb0fdedfb40f92ef6b8f3b2f2a3f3a8f62ffb3c00c904d507a8081b07a30347ff40fb91f8cff7e4f81afbaafd0200c801fd02d5035b04870465041204c903db037d04a5050c0750081c093e09aa088307f7053204720202012b0033006301e2039107180ce2102015f617cd18791725144d0f96096f0305fd88f63bf08fea4be643e4eee44ae8c0ed3cf4c2fabc00fc05c70a6f0fc3130c1749189b16df11ca0abf025cfbb9f52ef2a4f0c3f035f2e1f495f8acfc37005e02cf02fd01e7008a002f0130029202b301bfffd0fd4cfdd6fef90157054c07d9062c044b006afc5bf939f7b1f576f490f364f357f46af61ff9b6fb75fd04fe8efd87fc7afbd6fad6fa99fb0efde8feb500f70131025501f3ffd5fe94fe45ff4000570092fed3fa0ff6ccf16fef9feff8f16af51af9bafc8800eb04c209210ed210c910b70d6e084a0291fc4bf804f6c6f576f7cefa27ff8c03ef0685081c0822066a03ba0075feb3fc74fbc1fac9fabafb66fd4dffd7008b0146012e0070fe1efc26f9a1f522f296efe0ee75f0e4f3dbf7dffa12fc9dfb91fa51fab5fb89fea201a303e103bd026b0150011403310656092a0b070b610970076206c40632088509a6091708f004e50002fd17fa82f85cf863f9fefa85fc95fd2efeb7fed1ffe5019c04fa06e607b306b0033200c0fd47fdabfed4005e027d02430169ffb7fd72fc50fbc8f987f7c3f41bf21ff01cef2cef50f09cf22cf6dbfa0b00af04c707ee088b088907c1066e061206e8049d02ccffbffdadfdf4ffbc034307cd08bc07df04e4016300fb00d90237049803be00ddfc02faecf9f7fcef01a9063b090109b406c4036801deff63fefefb56f81cf4c6f0c0efb3f130f6f1fb920131068209af0b110dd70d120eee0db80dc70d690ea90f25115b12f412c612df118610f20e070d7e0a1d07d70207fe7df93cf604f5f6f580f894fb1dfe88ff0c0071008b01ac037306fa083e0aa6095807f8034200c7fcbff92bf71af5bdf36ef379f4c7f6e8f952fd760007032105fd06b6083d0a3f0b5c0b6a0a88083606360429036603eb0439077309c50a960ab2088005df01b0fe9bfcecfb68fc8afd13ff0e019303bb065a0aa90db50ff90f8e0e220cc1093f08bb07ae076c07910620057b030302b40034ff2ffdabfa29f853f671f532f5e0f4cdf3f3f12df0b9ef67f10ff59af987fdd3ffa60020019f02e605960a570f911236134811c30dfe0907075b05cd04c404b9047304f2035803c5022102180160ffe2fcbcf974f6e8f3ccf27af3eff591f961fd84007002fe0274024101b1ffd2fd86fbcef800f6bdf3ddf20cf452f702fcfb001305aa07d7085109140ac10b2d0ea6103012ef11bb0f490cbc08380673054706c307ac080c08a40512026cfeabfb3ffae5f9e2f9c0f9b3f96afaaefcda003f065a0bb00e6b0fbc0de20a5308c506fb05f2047402fffd3cf892f292ee43eda4eecef18ef5cdf8e5fac9fbb3fbf4fa03fa5df958f927fab2fb6ffdaffe1affdafe7ffeb9fef2ffdb019b0370041504e202ad013701a201880247037b03550365032504a305540765084708fd061905530312025601c500d6ff65feb9fc1efbdcf923f9c1f86df80cf878f796f668f5fdf3a2f2edf177f2aff494f87bfd7f02f806900a510d6b0f9510f60fb30c84062bfe8df5f8eeebeb5becd5ee49f13af2aaf112f141f22cf640fc80028d060f075104e9fff6fbfdf920fa8dfb30fd2dfe63fe61feb1fe8fff0501ce026d04680542057d03e3ffdafa70f5fcf092ee90ee57f0b2f2a4f4d7f5c2f644f8d2fa12fe1501b8026802af00a7fe4ffd32fdf3fd89fe36fe0cfdd3fbbafb9dfd470175057a080709e8062a038aff9cfd0afe4c0013032005cc0538051904190353025e01a8ffd5fc05f9dff448f1f8ee4bee4fefb6f1e1f42cf80cfb11fd29feb4fe22ffabff43008e001d00e3fe6cfd99fc38fda1ff610360077c0af50ba40b090aef07ce05c3039f01edfe6afb62f769f31df016ee90ed58ee11f076f259f598f8fdfb2fffbe014e03de03e503f2035604200504067d065a06ef05ab05cf055006a40602060804f70090fdc7fa5cf979f9b2fa5efc01fe68ffa80000028703f804d3058d05d003a60091fc6df825f569f389f35ff550f8a0fbb6fe2b01fc027404df055d07c0087709ea08d10662036dff19fc49fa39fa64fbd0fc98fd5ffd78fcadfb9dfb5ffc95fda6fe1dff0bffebfe31fffeff1501fa013502a1018f0083ffedfe0dffe1ff0801f1012b0283012d00e2fe91fec8ff5c0264058807b507d705ec026a006afffaff18015601d8ff01fd35fa04f942fa7cfd2f01bd03620486035d0229027503ce0519084709e8082e07a904e9011eff35fc36f983f6d9f4fdf43df722fb84ff0203b60490043a03ab018100a3ff7dfe8bfce6f97ef7b2f684f800fd20034609f80d8b103c11ad104e0f210dcd092305a4ff70fabaf645f5dff577f7cbf816f968f888f76df7b0f841fb74fe8601f4038305480689066006c105bb046503c901060048feb2fc6dfbc8fa01fb05fc73fdbefe4bffd4feb4fd9efc32fcb2fcd0fdd4fe36fff9fea7fe02ff5b0031026803e40238001dfc22f8bcf597f535f72bf91afa94f934f83ff7e8f770fa0dfe6c0165039a039b0270010401bd015d034a05f00603088f08c308dd0816096d09b709cf095e09eb0746058101e8fc2ff839f4b2f1f9f018f2c7f489f8d2fc2501ff04d3073c090e096007be040302f3ff25ffcbff8901c803f70585071b08ae073c06ea03280184fe91fccdfb4afc91fdf2feceffe1ff6cff0dff49ff39007401530257026b01f2ff82fe82fdfffcd0fcd3fc28fd1afedaff3d029b040c060906aa0480026200ebfe02fe28fdfffb87fa41f9edf8fbf93ffc13ffbb01d2036805d2064e08ad096d0a0e0a52086e05eb0157fe2efbe9f8e9f78ef81afb4cff4f040c096a0cc90d500da10b630903077b047d01e0fdeaf94cf6ebf38bf36df536f90cfecf0268062d0802084b06cc0355015cffe3fd84fca7fadff742f47ff0adede7ecdaee66f37ef996ff3e04b5063907d206a9065b079e087409de088506010396ff72fd07fde8fd12ff98ff29ff24fe47fd33fd15feacff8601370383044c057705f204c00314024f00e0fe12fef0fd56fe16ff16005d01ed02a3042906fe069f06d304c90103fe42fa4cf7a2f563f561f62bf845fa5efc4efe1000bf016e031d05c90650086709ac09c70894065603d4ff12fdd5fb4dfc05fe030048015b01670003ffe3fd84fd07fe55ff3a017b03c205840733087d078105df027a00f7fe55fef8fd17fd32fb83f801f6cdf488f50df861fb21fe52ffd9fe5dfdfffbb8fbbcfc71feddff32005dff11fe5efd0efe2f0009039b053007ba07c107e4076108f80812093b087f0647040e0224009dfe6bfdaafcb2fcd9fd1500e2028a058307ac086109140ac00acc0a74093d06690117fcbcf76bf567f524f7a7f914fc03fe7cffbd00da01a502e0025c022c01b8ff73fea6fd70fdb7fd4dfe2aff6f004602c204b707bf0a580d090f970f1b0fce0d090c260a54089b06ea041403ee007cfef9fbf0f907f9aaf9defb20ff7202d0049a05cb04fc021401e0ffdbfff600b10287040106cc06ea068e06de05fd040d040703d4017200f8fe92fd8ffc44fcdcfc38feedff60010902c101da00f4ffacff2e000e018801f60046ff33fde6fb43fc7efeeb0148057e073808cd07f8065b06ff0563050f04e4014fff20fd01fc0ffce0fca9fdbffd09fde5fbf2fac3fa82fbe5fc56fe30ff0dffd3fdbefb60f969f75df68bf6e2f7e5f9f4fb9dfdaffe4bffb7ff200073006c00e6ff11ff5ffe52fe27ff8100a101d901e90031ff8afdabfcb9fc46fd8efd0bfdeafbdafaaafacffb00fe4c00c7010402490175007800b101ad036a05da056f046f01e0fd09fbc8f94bfa21fc6efe53005b017701c80097ff31fec9fc8afb8dfac4f913f968f8e4f7e8f7dff8f8faf8fd3301db037b05210648066a069e068606a005b503330100fff2fd4afe82ff89006400bdfe06fc38f951f7ebf61df893fad0fd5e01ca04920735095709ef0753052f0252ff3cfd02fc75fb38fbf7faacfa8efac0fa3cfbe8fb8dfc06fd76fd28fe3dff8f00b9012d02990131007cfe0bfd35fcd2fb6dfbc3fa02fabef9b4fa38fddd00ab049707f108b7087207b805d103af011cff10fceff869f61df553f5e3f655f91ffcd7fe3c011a033a047004c903980260019a006f0096008300bfff41fe80fc2ffbdefaa5fb03fd33feb8fe91fe40fe8dfee9ff11022a0429056104f401d1fe32fc06fb86fb2efd1effb200c20185024b031e049a04500424037501f7ff4cff84ff0500f7ffd3fec0fc96fa6df9ecf9f8fbd6fe97019203b7045f05e1055b06a10664067905f9032302420085fe06fdf4fb95fb1bfc84fd75ff400141023e028401c100a8008d012703b804940565054904c6026d016b0098ffadfe69fde6fba5fa30fad8fa8bfcbffeb300ce01d7010901f2ff2fff2dff0a008c013f039a04220594040103cb008dfee9fc43fc95fc75fd50feadfe66feabfdd3fc1dfc8efb11fb97fa40fa6afa74fb6cfd0800c002ec0428067a061a064b05420406038301c5ff06fe8afc8bfb26fb47fbadfb1cfc7cfcc3fc05fd75fd2afe13ff0900b600b000c0fff7fdb5fb9df941f8e1f75df837f9def90efaf1f908fae2fac5fc75ff3c023304b20488030601e9fd07fbf5f800f829f833f9d4fad7fc11ff5c0198038505d20637078b06e404b00293001dffa2fe0bffd9ff770091003400d5ff0f003c012f034a05b806c4063e058f0287ff0cfdcefb0efc89fdb7fff201a603790458046e032102eb002f002300a30035014c018d0000ff29fdc5fb72fb63fc42fe8000b102b104ae06e4082a0bd90c2e0dab0b6f0853048900e7fd90fcfbfb55fb12fa57f8d7f65ff667f7b4f97ffceefe7e002b016c01e001e0026c044c061e088a095f0a810ad509520815066303950008fe01fc9dfafaf958fafdfb09ff3703a507f90af60b170ad905a20026fc9df949f98dfa6bfc2bfeaeff48014f03b905fd0759095309f907c8056c036a01e7ffc8fee8fd39fdb7fc60fc2afc13fc3dfce5fc38fe1e000a022b03db02100164fedbfb5dfa17fa61fa34fac8f806f6c0f24af0c6ef91f12ef58ef98efd6f002b0233030e041a0558066207c1072707820511034e00abfd84fb0ffa4ef92af98cf95cfa86fb03fdbffe880020024403b50360036f022801d7ffbffef4fd58fdc6fc2afc8efb2afb56fb65fc83fe910113053e082f0a320a19085a04e7ffcffbdcf845f7c5f6e6f65df731f8a1f9d8fbbcfee301c3040c07c908300a680b610cbf0c060c0b0a0e079d035d00c4fde6fb8efa76f97cf8b4f745f755f7f4f710f97dfa1bfccafd4eff5c00bf006b009effe8feeafeeaff9a013203bb039502e8ffa1fce4f977f860f8e6f819f991f8c7f7d2f7b8f9b6fddc026f07cc093c094c067e0278ff29fe76fe88ff63008b0047005300570184036e063609fb0a4a0b290a0508940587034202d001eb010902a0017900dbfe65fdbefc42fdb0fe3100da004300b5fe1cfd94fcb5fd2b00eb02c4040405d3031c020e015b01db02ba04e6059505c3032c01cafe5dfd1afd92fd08feeffd3bfd6dfc49fc57fd84ff1802ff034d04c7020a0048fdbffb27fc57fe60010f048d05ba052605b304f704cd056f06fb050904070126febdfc7efd0d003903a2056b06b1056b04ac03f80313052b064f061705ce022a00e0fd63fccdfb00fce6fc8dfefe00110460075f0a880c890d580d190cf7091907b2031b00dbfc84fa8cf915fac1fbebfdf6ff76014b02aa02d002bf024d025301c9fff2fd61fca9fb0bfc5afd12ff92006f019b0159010601d600be008000d9ffa1fee4fcecfa26f9fcf7ccf7c8f8c8fa4ffdbcff6e01fd017601520023ff57fe1dfe55febcfe2bffb8ff9200d7017303090516062106ec049d0299ff5efc71f92cf7a3f5cef4b4f45bf5dbf66af90dfd6501d1058b09ce0b310ce30a6e0878058b02e5ff6efd09fbdcf858f71cf7a8f8fdfb7100e3041f086009a508a9067204dd023d02380217025701ebff3ffe09fddffcc3fd2aff6100dd00760093ffe1fedefea0ffd600f10169020502e90076ff08fed1fcd8fb05fb2dfa42f95ff8a4f727f706f74ff7edf7ccf8ddf9fffa18fc31fd59fe97ffec003d024603c503a103f302f9010d01700026000600e1ff95ff2fffeffe1ffff3ff750175038c0541072a08ee077806f903d10077fd75fa32f8d9f67ef622f7adf804fb03fe4b0146044306b0065a059f0262ffc0fc98fb2dfc1cfe9200ad02db030d048a03a502950175003ffff8fdbcfcaefbcdfa06fa53f9c7f895f806f947fa41fca7fe170130039c041d057f04a902ccff7ffca2f91ff891f8e6fa74fe400256052d07ba07460720067a045d02c0ffc6fcd4f976f73df67ef61cf888faf2fc92fe01ff69fe70fdeefc8afd62fff8017c042a06ac0644069c054f059a052f066606a805dc0388018cffaefe32ffac003f022e034a03f902f802e003b005bd071509f808380750041a015cfe7cfc75fb05fbf2fa39fbf5fb38fddffe8300a401f10172018200a0ff24ff0bff04ffabfeddfdddfc38fc6ffca7fd80ff3a012802120247016a00150074002b01aa018b01d400f1ff7bffccffc900f101b002a402c0014c00adfe30fd04fc46fb0ffb74fb79fcf0fd87ffea00ed019f023903d70347041a04e4028c0093fdecfa82f9c4f96ffba5fd70ff50006c005600a10072014f027c026c0125ff4efcdff9a2f8ddf845fa37fc22fec7ff3801a7023704c90507079a0755073d0677044402e8ffaafde4fbfefa3ffb91fc81fe51003f01e10069ff84fd06fc8cfb2efc7efdc4fe60ff18ff27fe11fd5cfc58fcf3fcc7fd6efeb6fea9fe8ffec4fe56ff00005900100020fff9fd47fd83fdb8fe76000202b60260023f01d6ff9ffec8fd2bfd87fcc3fb11fbebfae2fb3efecd01ef05c8098f0cdd0dcd0db60ce90a8b087c058c01e5fc32f863f456f267f223f476f64af80ff9f5f8d0f88ff99dfba1feae01c7036f04e003e4026602ed025404fd0537078707de06960515048c02040170ffccfd36fce7faf7f94ff9c4f84af812f881f8f1f95afc3bffc9015003a3032e03ac02a5021b038c033d03d201a4ff80fd35fc2ffc2afd5afe08fffcfe76fefdfd02fe84fe1fff7cff91ffa2ff1900220163022303bc02000163fed1fb26fabef957fa46fbe5fb00fce1fb20fc45fd79ff6f028a052508c509380a96092a0852067004da02c3012e01f100cc007900d1ffe5feecfd32fdf8fc54fd36fe6effbe00ef01e3027f03ac036603b4029d014600e0fe86fd49fc46fb95fa56fabdfaf0fbe1fd5700fe0273056c07cd089109b9094f095b08fb06740521044803f702f702d00200024b00d5fd1bfbcaf884f798f7ebf823fbbefd39004202b9039b04fb040205d904a1047704620451042604cc034303a9022302c8018b013c019d008dff14fe65fcc5fa74f98ef820f83af8edf84efa64fc0bfff201c0042007d708c809e9093509be07c205a403d901aa0006007bff79feb6fc74fa80f8d9f719f908fcadffc1024f0436043e038302c7021104ab058e0609062c049301f7febafcb7fa77f8bcf5ddf2c0f066f054f231f6e3fa12ffd4011d039d033c0484054307a708bc080407bb03c2ff32fcd8f9faf854f963faaffbfbfc32fe47ff2500a700a900250035fffdfda5fc64fb7efa48fa17fb08fdd1ffc0020205fd059d056a044403db0252033204a604ea03ca01b8fe8afb1bf9f2f704f8d9f8def9acfa30fbb0fb8efc05fe06002e02ed03d904e1045004ac036d03ad031c044404c903ae025f01780061000e010502a0025d02250157ff93fd6cfc34fce7fc35fe9fffb0001c01d100ffff0dff68fe57fed6fe9eff480082004700e6ffc8ff3a0042019002a80334042704b6033703df029102fb01d7001cff21fd84fbd2fa2dfb4afc8bfd56fe79fe44fe46fefafe77004a02b5031e045c03c601150008ff02fff3ff7501fa02060464042e04a6031703be02a702a2027302f6012c014d00a8ff6fff86ff97ff3bff41fedafc89fbdffa25fb27fc4ffd04fef8fd58fdbcfccdfce3fde7ff7102e704cc06e30720089a0787062d05d203b102e4015201cd003e00baff84ffe1ffd7000102bd027a020c01dbfebbfc77fb6dfb68fcc1fdbdfef8fe95fe15fe0cfee7feaa00f60241050207c4075807e305c6038b01c8ffddfec4fe25ff82ff78ff01ff7cfe6dfe31ffb10061028f03bd03df026801040028ffdffee3fed4fe7cfe03fec8fd13fee1feedffd100460145010501ba008300650066009900280127026d0391041d05ca04b20355024b01fa00620121029e026502500187ff76fda0fb6bfa0ffa97fad2fb6dfd1affa200e901f002b80328041a047e036c022d011a006eff2cff1fff11fff6fef4fe31ffa6ff0f00faff19ff86fdc5fb77fa01fa61fa29fbd2fb19fc26fc55fceefcf7fd28ff160089009f009f00c50026019c01e901ef01bd016f0111018d00b9ff8afe37fd28fcc4fb31fc29fd1efe90fe58fec7fd7cfd05fe79ff71013803340438049103ca02500232022b02e10123010a00e7fe04fe7cfd4afd63fdccfd9cfedeff6801df02e703550447040704d703c603a9034b03a102d2010c015d00a0ff8efe03fd3afbacf9caf8baf842f9f3f989fa33fb6ffca7fecf013e0500085a093e09510876072a072d07ad06d2046d0140fdacf9eaf760f865fa9dfcc6fd68fd02fcacfa5cfa53fb05fd7ffefdfe6afe55fd8efc99fc64fd59fec8fe62fe6cfd99fca2fcdafd1000b9023a053907ae08a7091a0ace097708f00576029bfe0afb3df85af63cf5b1f4b3f46df516f7aff9eafc41002a035105b1067007a8075b077a06fd0410030e0152ff05fe22fd81fc05fcc2fbf8fbd7fc4dfefaff4f01d8017b0187007effbcfe44feb6fd9cfccafa9af8d2f643f660f7eaf90dfddfffcb01ce0263031b041f0515065806640522030f00f6fc7dfae3f802f88ef764f7aff7daf840fbd6fe17032807210a5c0bbb0a9c089f057402a0ff5bfda3fb64fa94f93ff988f981fa10fcf3fdd7ff71019f026c03f7034f046d04380492037c022901e9ff0affc6fe2fff140027011e02c102020318035103d803a4046d05b50513057c034301f0fe0ffde6fb62fb3dfb50fbabfb8bfc2bfe86003a03ad055c071008e2071207d3052604ec0120ff06fc26f917f73cf695f6c1f73df9a8faecfb33fdadfe69003302a50364044d048b038202a6014b0183012302cf022d03fe0235020401d5ff12fff5fe6afffeffffffeafec3fc27fa1cf89ff70cf9e1fbfefe3d010802ae0125016401c102af041406f105fe03e400dcfd0cfceafb13fd94fe79ff48ff33fee4fc1afc45fc6afd2eff0c019902a603390470046e043a04b203ae02230126ff02fd2dfb10fad6f961fa54fb39fcbffcf0fc22fdc9fd33ff5001a7038c056b061506cc041b0385014b0055ff5bfe2bfde5fbf3fad7fadefbeafd660084029603590302021f0057fe17fd6afc16fcccfb5dfbdffaa1fafafa08fc99fd42ff91003e0158013e015701dc01c502c5036e047f0409045a03db02e4027b035004e804d104c903e6018eff40fd69fb49fae4f908fa73faeffa5efbc6fb54fc4afdd9fe0e01b4034f06430812098e08f706e6040903d0013f01fc007d005fffacfdcafb47fa96f9d2f9b5facffbcefca8fd8efebaff2f019b027303480316024c00a3fec1fddbfd8cfe21fffdfeeefd4efcddfa52faf8fa9cfcaffe8f00dc019202ec0227035b0366030b032302c40042ff11fe9efd16fe54ffee005f022f0321034b02fb0092ff60fe87fdf1fc76fc03fca7fb95fb09fc22fdbffe920038025e03e903fb03db03d3030d047e04eb040005780445039601cfff60fe99fd7bfdc8fd23fe40fe14fed9fde3fd69fe5dff6b0024014101d0003500f6ff7200ad014a03af045405fc04cd033202a9008fff03ffeafe08ff24ff1cffe6fe8ffe2dfed4fd89fd45fdf6fc8afc04fc8efb71fbf9fb48fd3aff65013c0355049e045e040304e203ff0300046d030002dcff86fdb7fbfefa78fbcbfc5afe8fff1c001500d4ffbcff00008b0015014d010601540086fff4feddfe42ffe4ff5f006100caffc1fea4fddbfca2fcf2fc83fd01fe3cfe51fea3fea5ff9101370404073109180a7e099907e804fa0132ffb9fc98fad9f899f704f735f71ef88cf942fb0dfddbfeb1008d024a04a70569066c06c505c104b103ca0212027301d3003400c5ffb7ff0d009000e100b300040038ffeafe8bff1401f7026004ac04ca034e021901cf0070015202900294018eff64fd38fcc4fcf7fef8019d040b061b064a055e04ef030f045d045f04d203d702e101650191013c02fa02560310033002f900cdff05ffd2fe2affd9ff8400d5009d00f7ff3dffe1fe36ff390083018002bd02260212012000d5ff50004501290287023f029301f000a100a200a600510079ff48fe2bfd94fcbffc9cfde8fe530099019c0243036b03ed02bf01020008fe42fc0afb7afa75fac4fa3dfbdefbc0fcf1fd53ffa0008801d9019c0109015e00bbff1aff64fe90fdc7fc54fc75fc36fd5dfe84ff4b008f0072003a0024002f001b008cff4efe70fc53fa85f88cf7b2f7fef836fbf3fdbc0016039c041105780411034a0188ff06feccfcbffbcdfa13fad5f94dfa7afb14fd9efeaeff2e006d00e500ec0174030005de058b050104b90176ffedfd71fdd7fda0fe3fff5afff3fe5dfe00fe22fec8feb0ff7d00f1000e010e014501e301cd02aa031104c603dd02b501c30056007900f6007e01dc010b0230027c020c03d10394040605e4041104ab0208019effd6fedafe87ff7e005401d6011f0280023e0352045305a305cb04c8022400b2fd28fcc2fb31fcd6fc34fd3dfd5bfd1bfecdff3502a0044406b0060606e404fa03a903d703180405048c03f902b402f2028903fc03cb03c102080108ff2afdb4fbbbfa4cfa87fa91fb68fdc4ff1602c70380046004df037f0378039d037e03c70291015c00caff36006a01b10235037a02a70070feb8fc10fc75fc5efd18fe36fed1fd6dfda5fdbefe74001202d1024202860047fe5dfc75fbc4fb01fd94feefffc20015013b0190013d022003d703ee031f03870197ffe4fddafc89fca1fcaffc6cfceefb9cfbe1fbdffc44fe6effcaff33ff0dfe13fdeafcc2fd41ffb9009201a0013201db001201ef01260330049904310411037e01c1ff0efe88fc4cfb79fa28fa5dfafafad1fbbafcacfdbefe07007f01e902e703240485033902a00012ffbcfd91fc6ffb50fa6df925f9c5f94ffb63fd65ffc700540147011c014a01f701df027b034b031d022300dffde6fb9ffa2dfa74fa35fb35fc48fd50fe2fffc9ff0800f0ffa7ff6dff76ffd7ff760010015e013801a700d8ff0aff66fefafdb6fd83fd57fd3dfd51fdaffd62fe5bff720075013d02bd020103280345034e031b037e026301f1ff87fe9dfd8dfd63fed1ff57017802f402d7026002d1014801b300effff3fee7fd23fd00fda9fdfdfe9b000702e1020f03b7022302a20164016f01af01060250026e024602cd010a0122004dffbcfe84fe9afedbfe2cff91ff2a001401460278033c0431043e03ad01150017ff12fff7ff570197023a0317035c026b019c001700c4ff65ffcdfe01fe43fdf3fc5bfd83fe2100b801d2023503f9026f02f501be01bf01c201900113016000aaff22ffdffee4fe2fffbeff9500a601c402a103e703600311023d0046fe80fc1bfb1bfa78f937f972f94efad1fbcafdd5ff77014f0240027401480025ff5bfe10fe44feddfeb2ff97006301f2012b0204028101a60076fff1fd24fc37fa7cf85af72af70cf8d0f9fbfbf8fd51ffdaffbbff49ffd9fe98fe7bfe5bfe13fea3fd2ffdeffc1afdcffd0cffb00080022b045605af050d0583035b0102ffddfc22fbd5f9e1f840f80af877f8abf998fbe8fd1b00bd019702bc027202fe018001f6005400aaff2eff22ffacffb200df01cc022e03fc0261029601bb00c8ffaafe68fd3cfc81fb7efb32fc47fd37fe9bfe6ffe17fe2cfe1affdc00ef029d045705fe04e1037a022101daff76feddfc4dfb60fac5fad7fc4f004e04b0078e099a092408e3058403680190ffcefd06fc60fa3af9fbf8d5f99bfbcdfdceff2501b001ae019801de01aa02cd03d5044d05f904fc03c502d5018001bf0136026802f801dc0067ff1efe78fda1fd69fe58ffeeffe2ff4aff90fe3afea2fecaff5301af0268035503ab02d7013e010c01270149013e010501de001701d901f702f303310448033d018cfef7fb2afa7bf9c9f9aafab2fbaffcb6fdfcfe95004e02b90362041404f7027c0124003dffd1feb4feb0feaffebefefcfe7dff37000801c40147027b025702d8010b010b0004ff1efe71fdf5fc8dfc25fcc6fb9ffbf3fbf2fc9afeaf00d202a504e6057a065b068b05110403029cff3bfd53fb3afa0afa97fa85fb81fc63fd3afe30ff56008d018102da0267024001bdff4dfe48fdcffcd6fc39fddefdbdfed2ff0e0146023403930337032a02ae002eff1dfecdfd47fe4bff61000f0110016e007cffa4fe25fef9fde0fd93fdfdfc56fc06fc69fc96fd50ff2201a002930303041804ec0372038602100132ff4efde2fb53fbbbfbe4fc60fec2ffc9006c01c601f201f401c0014901a4000900bcffedff980081014f02bd02b0024502b0012201a8002e0090ffb6fea4fd7dfc74fbbcfa77fab4fa6efb92fc04fea5ff5301eb024b045005e205fc05af051e056f04ba03fe02280228010700ecfe10fe9ffd9cfde1fd32fe65fe76fe8ffee4fe94ff89007d011a0223029001930080ffa6fe30fe20fe56feb0fe19ff91ff2200ca007101f30131022b020302ec01090251029102880211023e0153009eff4dff56ff80ff92ff76ff47ff38ff6fffdeff4f0081005900f1ff8bff61ff79ffa0ff82ffe8fee3fdcdfc1efc2efc05fd5afec3fff200db01a902900394047805d6055f050e0435025000cbfed0fd44fdf1fcb6fc98fcb7fc23fdbdfd3cfe56fef0fd33fd7efc2dfc73fc45fd71fec1ff1d018102ee0348055706d906a506c80581042203ed01f50023004bff4efe2cfd03fcfbfa30faa9f95ff957f9acf990fa27fc6efe1d01b603ae05a5069006c105b904f303a503b103bc0361036b02ec0034ffa8fd95fc15fc0efc4dfca2fcf8fc55fdccfd6afe29fff7ffba006301f1017102ef026f03e0032104090476036402f3006aff25fe75fd80fd36fe51ff74004d01aa018501f100110007fffcfd24fdb8fce9fcc4fd29ffd3006e02bc03a70436057a057b053405a304db03ff0233028201d4000000f4fecbfdcbfc3cfc35fc8bfcdffce5fc94fc3dfc5bfc4afd04ff1e01fc0227048504620431043f048c04c9049c04d50393022b01f5ff1dff91fe1ffea2fd1cfdbcfcbafc37fd22fe43ff4c00f7001b01ad00c4ff97fe77fdc2fcc5fc9afd15ffcc003802ef02d30213021b015000e9ffd3ffcbff89fff0fe20fe67fd12fd44fde4fda9fe41ff7fff6dff45ff49ff9dff2c00b300e6009f00faff4eff06ff69ff6f00ba01bd02f3021b02560013fee5fb47fa78f978f91ffa42fbc6fc9bfea900bc027b048905a805da046903cb017500a9ff61ff5bff3fffcefefdfdfcfc1bfc9ffba9fb23fcd8fc91fd33fec5fe6aff3a0030011b02b902d4025e0282018d00cdff6fff6fffa3ffd6ffe3ffc8ffa2ff9effdaff5600f4008301d201ca017301ed006400fbffc2ffafffadffa2ff80ff4cff19ff02ff1cff6effe9ff7000e60040018a01e2015b02ef026e0397033b03610250016d0009003200a800fe00e0003c0052ff8dfe45fe92fe43ff01008300ae009c007b0070008200a200c000df0012016c01ef017e02ef021b03fd02aa024a02fa01bc017601050158007cff97fed7fd55fd13fd03fd19fd59fdd7fd9ffea7ffc200b301440265023002dd019f019201ab01c901c50187010c016a00bfff2dffcefeaefec7fe02ff3fff64ff68ff53ff37ff1fff05ffd2fe75fef2fd6efd25fd4bfdf0fdf7fe1e002101da014a028c02bc02dc02d2027802b801a00061ff3afe5dfde4fccefc12fd9ffd65fe41ff010069005400c8fffafe39febefd97fd9ffda7fd9ffda5fdfbfdcffe120071017802d6028402c301f70063000e00caff63ffcbfe25feb0fd97fdd6fd3cfe87fe8efe53fefcfdb6fd9cfdb5fdf9fd5efedffe75ff13009e0002013b015e018b01d4012d02620237028801610002ffbefddbfc75fc7dfcd0fc52fdfdfdd3fed0ffd600b30131023502cb011a015600a6ff1bffbbfe84fe76fe8ffebffef1fe10ff17ff1cff41ffa4ff47000a01bc01320257023002ce0143019900dcff24ff9bfe71fec1fe83ff7f006101dc01c90139017100cbff91ffd7ff790027018f01840114017700f1ffa0ff72ff34ffbefe1cfe93fd7efd11fe2dff59000201c600b7ff59fe68fd7bfdb7febc00dd0273042a051c05a8042e04d003630398023e016fff98fd4cfcf5fba5fc0dfea0ffd60062014701c5003000c9ffa7ffbaffd6ffd5ffa1ff4cff02ff00ff6fff4f0068016002e002c60233027b01f500cb00e400fd00d5005e00c4ff52ff42ff9aff2900ab00ed00e800b60079004000ffffa6ff33ffc0fe79fe83fee4fe84ff3700d7004d01900198015701c500eefffefe3cfee7fd13fe9bfe2dff82ff80ff53ff4affa3ff62004201e5010d02c1014601ee00df00fa00f2008800bdffdbfe4bfe51fee5feb0ff42004b00c5ffebfe0ffe6ffd1cfd09fd24fd6afde9fdabfea8ffc000c40190020f033a0311038f02b101860039ff07fe2efdcdfcdbfc34fdb4fd54fe2cff5600d0015b038904e70439049b027b006bfedffc05fcc2fbd7fb11fc69fc01fd01fe6fff1c01ad02bd030d049803960265015d00b2ff62ff41ff18ffc6fe57fe05fe14fea7fe9dff98002201ed000100c2fec0fd76fd05fe2dff70005c01c001c201b801e7015502bd02ba020502a700fefe91fdd0fcdbfc7dfd4dfeecfe35ff4dff80ff13000f013e024303c503a203f40207023301b3009500bc00f4000d01ec009300130084fff4fe63fec7fd1ffd78fcf6fbc7fb14fcecfc37febfff3f017d025c03e003250452047f04ad04c0048b04e203af020b0139ff9bfd88fc32fc89fc4afd19feacfee6fedcfebbfeacfec0fee8fe06ff0bfffafef2fe18ff84ff36001101e8018f02ea02fb02e002bc02ab02a8029102350271014e0002ffe3fd39fd1efd71fde3fd2afe26feeefdc6fdecfd77fe41ff00006f0072002500c7ff92ff99ffc4ffe4ffd7ffa4ff77ff82ffe2ff8000220187018d013e01ce00710047004d006600730068004a002a0013000b00110027004e008100ad00b4007b00050076ff04ffd9fef5fe28ff33ffeffe76fe14fe1bfeacfe98ff7000c7007100a0ffc8fe61fe9dfe58ff3000c800fa00ea00dc0009017201e7012202fa017301b200e6ff25ff72fec7fd2efdc7fcb7fc0efdb7fd84fe4afffaffad008301870291035904a0045a04bf032803da02ce02b5022302d800f1fee3fc40fb72fa86fa37fb1ffcf9fcb5fd6ffe47ff3a001f01c1010102e7019e0154012601150112010b01f100b7005100b8ff00ff57fe00fe2ffeeafef7fff5008a0194013601bf006d0046000f0079ff61fefffcdafb8ffb7bfc82fe1c018f034a051e06450625060706e80581057804a4022e0085fd29fb74f982f83bf870f800f9e2f91afba3fc6bfe4b001902a903cf0465054e058b044203bd01530045ffa7fe5ffe42fe33fe34fe61fed1fe79ff2b00aa00ce0099003800e4ffc4ffd4fff3fffaffdeffb4ffaaffe5ff670006018501b10182011f01c800ae00d80021014c013001d0005f001a0026007100b700ab00210028ff0cfe30fde0fc32fdfefdf7fec9ff3b003c00eaff7aff22ff08ff2eff7cffc5ffe6ffd5ffa5ff7fff83ffbaff0b0047004a001400d2ffc8ff32001c014f0269030604f4034c036602a8014c0145014a010c01690089ffc6fe74feaafe31ffa2ffa6ff2dff71fed5fda4fde2fd51fe99fe85fe29fed7fdf4fdbafe1600ab01fd02ab038f03ca02a901800086ffcefe48fedafd77fd26fd02fd2afdb1fd93feaaffbe009101f601e2017001d90054000300e0ffcbff9dff51ff0bff0cff8dff9700f3013e0310043204af03cc02dd011c0195002c00b9ff24ff73fec5fd3dfdf6fcf2fc28fd84fdf3fd66fed3fe32ff7fffb8ffd8ffd9ffb7ff71ff13ffb7fe80fe90fef1fe8dff3100a100af005c00d5ff5dff2eff54ffa8ffe9ffe6ffa0ff51ff49ffbeffaa00c601b7023d035803390321032e0347033003b502d201bd00caff3aff18ff31ff37ffe8fe33fe43fd62fcdafbd3fb47fc0bfdebfdbafe63ffe9ff5b00c9003a01ad0113025a026a023102a601d300d6ffdafe0afe82fd47fd4ffd8bfdf3fd81fe2effe0ff7000bc00b80080004a004c009a001d01a301000226022e023f027402c5020e032b030b03bf0266021a02da018c010b0140002affe8fdaefcb2fb28fb2dfbbefbb7fcd8fddcfe8bffd6ffd4ffb6ffadffceff0f004c0065005200290012002800630098008b0018004dff6dfecffdb1fd17fec3fe5effa4ff90ff59ff54ffc1ffa700d601fd02d903490457042504d5037e032503c6025802d30133017c00c0ff1bffa6fe69fe56fe4bfe2bfeedfda8fd82fd9ffd06fe9bfe31ff99ffbeffa3ff65ff24fff9fee9fee7fed9fea5fe3efeb5fd36fdfefc3ffd04fe2bff68006701f001fd01b90162012d012601370136010a01bb0076007400db00a10190025603af038603fb024f02c301750153013001e3006400cfff54ff19ff1cff3cff44ff0eff98fe02fe7efd38fd41fd88fdecfd49fe8cfebcfeeffe38ff99fffcff3b003900f0ff77fffcfea5fe84fe8bfe9bfe97fe76fe4bfe35fe55febdfe6cff4d00440134020303a9032a049804000560059c058705fa04ef0392023101150061fffdfea8fe25fe66fd9cfc21fc43fc17fd66fec6ffce0045013501d70071002f000f00f0ffabff2bff74fea6fde5fc54fc0bfc13fc67fcf0fc89fd10fe6ffeaffef1fe5cff0600df00b8015c02ab02b002930283028c02970274020402510195001e002300a60071013202a402ae026702ff019f0155011301bf005000d5ff74ff55ff88fff9ff7100af008000d8ffd7febafdc7fc2cfceffbf3fb04fcf8fbc4fb84fb6ffbbefb8bfcc4fd30ff880093013a028e02b102c202cb02bc027702e9011b0133006dff05ff20ffb7ff96006801db01bf0127016200d8ffdbff780072015e02de02d1026002e101a001b80101023002060271019700bcff1cffcdfeb2fe95fe3bfe8cfd99fc9cfbe1faa8fa0bfbedfb05fdf7fd7dfe82fe2bfec3fd98fdd3fd6dfe34ffefff7a00dc003b01bf0176024103e3031e04d90330036602c10167014d0146012401d9007f0046004e009400ef002e0136011301ed00f00029018801e40118020e02c60148019f00d5fff6fe19fe57fdc6fc6dfc3efc22fc09fceefbe1fbf7fb40fcbbfc57fdf8fd8cfe0dff85ff08009c003701b701f601dc017701f900a400a60006019b0126026f0268022c02ed01d501f30132026c027d025402f6017c010801bd00b100ec005a01d60133024a020f028d01e100240061ff91fea7fda3fc9afbbafa35fa32fabafab5fbeffc2efe42ff12009e00f30020012c011601db0081001700b0ff58ff14ffddfeb0fe91fe88fe9ffed4fe23ff84ffffffa300790176026c03210465043304ba0342030e0333039503f4031404d2033403540253014b004dff64fea0fd0ffdb6fc8dfc7bfc68fc46fc1afcfcfb06fc4dfccdfc71fd19feacfe20ff7bffccff15004c005a003100dcff82ff56ff7cfff1ff8700f9001301c9003f00b6ff69ff70ffbcff23007d00b600d300ee0020017801f1017602ec0239034e032c03e502930254023a02470268027b025c02ef013201360020ff12fe22fd55fca1fb03fb86fa49fa6dfa02fbf6fb17fd2bfe06ffa3ff1d0098002501ab01f701d0011e01f8ffa2fe72fdaffc81fce5fcbcfddcfe1d005e01850279031e0462044004cd033103a002470239026502a702ce02bd026f02fa017c010f01bb0074002600c5ff4fffcefe51fee3fd87fd3efd08fde8fce7fc0afd4efda7fd00fe44fe65fe64fe4efe3dfe49fe88fefcfe98ff3900b300db009e000b0051ffb7fe7afeb5fe59ff31000201a1010502400269029002b102bd02ac0282024f022002f601c5017b011901ae005c003e005a009a00d400df00a40029008affe9fe64fe06fecffdb8fdbbfdd8fd0efe5afeadfeeefe06ffe8fea0fe50fe27fe4afec4fe77ff2900990096001a004dff76fee2fdc2fd1afebffe6dffe7ff12000200ecff05006b000f01c6016102cb020e034c039e03ff0349044a04de030a03fa01ec0012007eff1fffd2fe79fe0ffea6fd5dfd4cfd7cfde1fd69fe03ffa1ff3b00bf0012011701bc000d002fff5dfeccfd94fda7fddffd0ffe20fe16fe09fe15fe44fe8cfedcfe29ff78ffdfff720033010902cc025003800361031103b7026d023a020e02d4017f010f0192001b00b9ff73ff4cff47ff6dffc0ff3a00be002401460111019300f5ff6aff13fff8fe0aff2eff54ff7affa3ffcffff1fff4ffc4ff5cffccfe2afe90fd09fd99fc3ffcfefbe7fb0cfc7dfc3dfd42fe73ffb000d201bc0257039c03940357030403b6028102670263026802670256022e02ef019b013901d20070001c00dbffaeff8eff6dff3dfff1fe8cfe22fed9fdd5fd29fec5fe7aff0e00550047000400bcff96ff95ffa0ff8fff48ffcffe41fec1fd63fd2cfd13fd12fd2efd73fdeafd8efe4cff1200d0007f011b029c02f6022103270324033603660397038d030c030102960030ff3cfe00fe74fe46ff040056002600a3ff20ffe5fe0cff78fff2ff44005b0042001600f0ffd4ffb3ff7dff2bffc7fe6cfe36fe37fe72fedafe52ffb8ffe9ffd3ff78fff9fe8cfe66fea7fe45ff0d00b9000e01fb0098002100d0ffc7ff05006a00cf001a01440159016a0180019a01ac01a9018d0158011301c4006d000d00a4ff3dffeffed7fe0eff97ff5d003001de01420256022c02df017a01f500390037ff03fed1fce9fb7dfb97fb0bfc91fceafcfefce4fcd5fc04fd8dfd63fe62ff61004301fd0193020e037803d6032c0471048e046104cd03cb027a011d0002ff5afe1efe19fe0efedafd92fd7dfde3fde6fe5c00e20104037b034803ad02010281013301f1008c00eeff2eff7bfe06fee1fdf7fd1afe1afedbfd62fdd4fc68fc54fcbcfc9dfdd2fe1c003e010f028702b802b50284021b026e018a009cffe2fe8ffeabfe0aff66ff88ff69ff38ff40ffbaffad00e5010c03d1030b04c40326036602a801f30041008cffe0fe5efe2efe68fe06ffd9ff9f001a012901d2003a0092ff04ffa4fe6efe4ffe2efef4fd94fd13fd90fc3ffc57fcfbfc21fe8cffe100ce012f021c02d801ac01bc01fb0137023e020202a4015b0157019601e301ed0172016a000effc4fdeefcc0fc2efd00fef1fed7ffa90070013102d70239033803d10221026001b400240097fff4fe3dfe97fd2ffd1cfd4dfd8efdaffda3fd8afd93fde2fd6dfe07ff7effbcffd3fff7ff5200f200bd018202120356034d0303038902ec0137017400b1fff9fe57fed6fd8cfd8bfde0fd7bfe2fffc0ff0400fbffdaffedff66003a011d02ab02a1020802350198007e00e5008501fb01ff018901c900070071ff0affb2fe3dfe98fdd2fc17fc9ffb95fb0bfceefc0efe27fff6ff4e002b00bdff53ff3effacff8a008d015702ae0298025f025f02cf0294034a047d04e903a9022601ddff16ffbefe80fe03fe2dfd3efcaafbd7fbe0fc7ffe35008a0141026c024d0227021202f801a601f300e5ffaefea2fd09fd05fd81fd3bfee2fe3bff40ff11ffe4feeefe49ffedffaf005a01c201d601a1014201de008d00540029000000d5ffbbffcbff13008a00060150013c01ca00250095ff52ff69ffacffd6ffb1ff3fffbbfe78feaafe4eff2800ed007301c50114028d022f03c303f50385036d02e40045ffe2fde4fc44fce3fba8fb9bfbdafb81fc89fdbafec0ff5b007e005600270019001c000000acff45ff27ff9fff9c009c01f0013801c5ff8bfe9dfe79009d03b10643088f07eb048b01cefe83fd9dfd6afe23ff5cff2ffffcfe13ff77ffe3fff7ff7dff8afe7ffde9fc46fdc2fe060137033b043503070093fb7bf777f58df684faf3ffda0483073a078004b80072fdbefbe3fb74fdcaff6a023e052e08bd0a0e0c0d0b1207860019f951f375f166f406fb8d02ca079a08e10486fe73f82df5cdf5bef94eff9c045808070ac909fb07ed04ee0083fc90f84af6cff69cfa15017008260ed40f340ccc03eef8f8ee26e961e99deff4f96005c00eba134013b10dab04a6fa5bf219ee16ef07f52bfedc07700f0213f611ee0c6f055ffd8df660f29bf13bf470f9ccff94053e09d809460741022dfcd1f6e7f3aaf457f9e5002e09930f0012c80ff009b40271fc9ff858f7a4f75df8f4f8adf92efbbefdc100e802f602a100f9fcfef989f939fcf900830597074206670249fe40fc6efd20014705b8076c0705054b02fc00ad0179039c049a03300085fb7af79df562f6daf873fbdefcb4fc8ffb9bfaeffa01fd7d007904de07e309510a8a0944081e074a0677051204b60187fe3efbd3f8f5f7acf856fa0cfc1bfd61fd41fd53fdfafd32ff9f00cb016902700205025c019400bbffdcfe12fe8bfd7afdfdfd06ff5d00b201b9024a0363032303ac0216026801a300dcff38ffe0fee2fe27ff77ffa1ffa3ffaeff130004016902d903c704c104ad03ce01aaffc2fd64fc97fb32fb00fbe9fafffa6dfb55fcaffd37ff790004019d0075ff21fe67fde2fdadff4702c8044a065306100533038f01b500b5003301a901bd016201cf004f000f000300f0ff8bffa2fe3cfda6fb69fa17fa0ffb40fd11009902f803c2033502140044fe52fd60fd42fe89ffd500ed01bd0234033503a6028c012000c6fee2fdaefd25fe0bff14000501c00133024b02ee010f01caff6ffe6dfd23fdadfdcdfe0300cb00df004c006cffa7fe42fe44fe85fedafe31ff96ff1800a80016012a01cf003600c7fff0ffe5007a0234047d05ec05670523047502a600e0fe2ffda1fb56fa85f961f9fff948fbfcfcc7fe5f0095015c02c102e302da02b3026702e401210128001fff41fec2fdbefd2dfee3fea8ff4d00b700e200de00ca00cb0003017f012802bb02dd024202d600dcfedcfc73fb0efbc0fb3efd04ff9800b2014f029302a1027e0210023501f0ff7cfe44fdbcfc27fd6dfe1d0092013d02e701cc007aff94fe85fe55ffb1001a0224039b0386030c03510261013b00dffe6afd17fc2bfbd7fa25fbeffbf4fcf8fddafea0ff5f002601e0015d026f020b026601db00be002501d1014a022a0256011d0013ffbbfe49ff7d00d001b402da0247024301270034ff83fe09feaffd64fd27fd09fd26fd9efd78fe9affba007a018e01ec00dfffecfe8ffefafef4fff20067010e011300fafe57fe7dfe5bff8b00900118022202ee01cc01ee014a02a302b30252028c019d00d2ff67ff6bffb7fffdffedff50ff29feb7fc64fb99fa98fa5ffbadfc20fe65ff5c001601c00177023003ba03d90372039b029901c1004c0044008600d400f800d7007500ebff57ffcbfe53fef9fdcdfde7fd5cfe2aff2e002501c501dc016a01a000caff20ffb7fe7afe49fe1efe14fe58fefefeeaffd00059015901e7005400fcff13008c002901a201cb01a8015a01ff009e0028008cffd2fe24fec4fde9fda4fed1ff1f013902df02fd02a302f4010b01f4ffb5fe61fd2afc52fb16fb89fb8efce1fd3cff6d0068012e02be020403ec027802d0013a01f3000c015c0196017701f30036008bff29ff18ff2fff33ff01ffa2fe40fe0cfe20fe72fee3fe4dff96ffb5ffacff81ff41ff00ffddfef5fe57fff7ffb2005d01de0136027a02bd02fa020a03c0020202e700b7ffcdfe66fe89fefefe74ffa9ff89ff2fffccfe89fe77fe93fedcfe58ff0e00ee00c50145022a025c0108008dfe51fd91fc55fc7afce0fc7ffd6bfeb0ff3701b602d0034004030457039a021802e601e501df01ab013e01a500f3ff34ff71fec0fd48fd35fd99fd54fe1aff91ff80fff2fe2dfe95fd77fde6fdbffebcffa0004d01c301160257028502940275022202a6011d01a40052002f002c002f001c00e4ff8fff39ff08ff19ff6cffdeff34003200b4ffcafeb3fdcffc70fcbcfc99fdbefed6ffab0036019301df0118021b02bf01ff000d0047ff02ff5aff1b00de003e0113018300e6ff96ffbaff3a00d6004d0182017b01580134011b010401e200af006d002700e2ff9aff43ffd5fe50fec0fd42fdf0fce3fc21fda3fd53fe15ffc9ff53009b0097004f00dcff66ff1cff20ff7dff29000301e501af0248039f03b0037f031a039b021a02a5013501b6000c002aff18fef3fce2fb09fb85fa6ffadcfadcfb68fd56ff5a01100325047404180458038d02f5019e01630112018200b7ffdefe36feeffd14fe81fe01ff66ffaaffe6ff4100c4004c018f0145015000d9fe48fd13fc92fbdafbc5fc05fe51ff7900660111027c02ab02a8028902630245022902ff01b2013f01b1001d008fff06ff7dfef4fd88fd63fdadfd74fea0fff60032021e03970394031b033f022101f2ffe6fe1cfe98fd3ffde9fc88fc35fc29fc95fc7dfdacfec4ff7800b000950077009600fe008401e501f101a9013a01e600de002f01c5017202040352033f03c202ee01e700defffafe4afeb8fd20fd68fc99fbe7faa2fa0bfb36fcf7fdecffa701dc0276039703810367035a0347030f03a202130288011f01d5008600020031ff30fe40fda5fc81fcc3fc35fda4fdfefd58fed1fe76ff2b00bb00fb00e30090003400f6ffddffd7ffd2ffc7ffc2ffd7ff0c005700a900f6003e018a01d7010f021002c2012a017200dbff97ffb2ff0c0068008b0064001300cfffd2ff2e00c300510194016701d300090043ffa3fe2bfec2fd47fdb2fc18fca5fb89fbddfb9efca3fdbdfebcff7f00010154019301da013e02bb024003b8030c0432042b04f5038903d802d701880007ff8dfd5efcb5fbaefb3afc22fd1bfee1fe4eff69ff5eff63ff9cff0b008d00f2002201270123013e018201cf01f701d5016c01e5007a00480042003700f6ff6fffc2fe2dfee3fdf3fd3dfe87fea1fe80fe41fe19fe3bfec1fe9dffa6009d013e025802db01e300bbffc0fe40fe56fee7fea7ff4800a000ba00c100e3002e018401bb01c401b301ba0100027702d702c9021802df0085ff8cfe40fe97fe3cffc3ffecffc2ff7aff41ff15ffc6fe26fe3ffd69fc15fc8dfcb8fd13fffeff110058ff4cfe92fd9dfd78fed6ff4401670222038803b403b003770301035d02b4013501f600e800e100ab002a0066ff83feb4fd2ffd1afd7dfd4afe55ff59001d0186019d018e018c01ab01d201d2017c01c400d6fff5fe5dfe20fe26fe35fe23feecfdb2fdabfd01feb6fe9dff780013015a01630160017701b401ff012602fc017801ab00c2ffe8fe3bfec3fd83fd85fdcffd5efe1effdcff6600a400a00085008400b60007015001710165014a014c018001d0010d0200028b01c800f3ff54ff23ff6aff00009e000001fa009000f2ff5bfff0feb5fe86fe3afec7fd54fd1efd5bfd0cfeeafe92ffb8ff55ffb0fe3bfe4ffef8fef7ffe300630161010d01b4009600c80028017c019a017b013401ef00cb00cb00dd00eb00e300c100940067003b000e00d8ff97ff5dff4bff78ffefff9d004b01bc01c6016001a700d3ff15ff83fe1efed8fdabfda3fdd4fd39feadfef7fee8fe85fe19fe0efeb2fe0400a7010303a1035f037a0261017200c6ff3bffa5fe00fe79fd5afdcdfdaffea9ff5b00930069002c002b0084002001c3013202570241020b02d601b301a3019b018f01640101015b007fff99feeffdc0fd1ffef4fef9ffd80051014e01dd00210049ff77fec3fd3ffdf6fce2fcfcfc39fd8ffd00fe96fe4cff06009900d700ac003900c5ff98ffd6ff6d0016018701a50188016e019201fa016d029d0255029b01bd002d0041000d01510290033904ed0390025d00d6fd95fb1bfab0f953fabefb87fd46ff9d004f0148019f0094ff93fe0ffe4efe49ffa300c8013c02dd01e700dcff39ff35ffadff5800f70079010002a7025503bd0385038402e7002fffe7fd57fd66fda8fd9dfd05fd04fc05fb87fae0fa0ffcd3fdd0ffb2013c035404e704ea0469049203ab020102c801f401430261021002410128001cff71fe66fe16ff6a001e02c703d704cc046c03e400c9fdeffa0cf95ff8adf865f9f1f90ffaf1f900fa99fad4fb74fd13ff74009e01c8022904b8051607c1076207fd0505042302e3006f009500ec001401ee009d005500380048006a0084009b00be00e600ef009c00b5ff45fea0fc42fb99fad3fac0fbf4fc03fea8fed5feb6fe87fe7ffec8fe7fff9e00fe0159034b048a0409040103d701f30080005e004600fdff77ffddfe6cfe37fe22fefbfda4fd3afd12fd83fd9dfe1d008701620284022402a001440121010101a500ffff43ffbcfea4fef2fe60ffa1ff9fff80ff90ff1200090134023c03db03f403a20319038002f2017501f80062009effa2fe7dfd65fc96fb33fb35fb66fb7efb5ffb27fb1dfb80fb60fc85fd9dfe7fff3f001b014b02c30329050c063106b105ee04580419040104b803f502b90154002fff86fe54fe62fe6efe59fe38fe2afe3ffe6efe96fe9efe8cfe82fe99fedbfe36ff87ffb3ffb8ff9fff70ff34fff5fec6fed2fe4aff37007301a80270038c030e03410284011801fb00f000b7002d005bff6afe86fdc0fc13fc83fb25fb1efb99fba6fc25fedaff8201db02c4033a044a041104ba035f0304039502ef01f200b2ff75fe97fd67fdfbfd14ff450028018a01790141012d016201d5014f028c025d02bc01bf0091ff64fe57fd73fcbefb3bfbedfae2fa23fb9ffb33fcb8fc0dfd35fd63fdd5fdbbfe2400ec01c9037105a80643072d076a06100554038e011c003fff0fff65ffefff5f0086005e000400a9ff6dff64ff91ffe5ff3f0075005600bbffaafe55fd0efc33fb03fb7ffb79fcacfdd8fedcffb900770112028102b502a8026b021d02d10183012801ad00180093ff4dff61ffc4ff44009c00a3006000f9ff9dff6eff6bff7fff98ffaaffa8ff84ff26ff7afe8ffda7fc16fc24fce4fc1ffe74ff96006401f4017b021c03c5034e048f0476041d04b0033e03be02190243014b0060ffb0fe4dfe2bfe2efe3ffe56fe7bfeadfed0fec3fe71fee2fd49fde5fcd6fc10fd5bfd6dfd14fd5bfc89fb08fb44fb77fc8afe17018803500528062b06c0055e054f058405a905660598046c0344026e01f1009800120036ff28fe42fdd3fcf5fc71fde3fdfefdbbfd4ffd0cfd2ffdbafd74fe12ff5aff31ffa8fef5fd53fdf9fc15fdb5fdbffe01003a012402a102c002b002ad02ea02750337040805bc0526061d067f0531042d029effe4fc7bfad8f833f870f835f918fad1fa5efbf2fbc4fcecfd54ffc8001a024303490420059f058705b00433037701fcff25ff0fff80ff12008700d00005015801e90193022003680336037a025201dbff41fec5fc8cfba1fa08fab9f9acf9f2f99efaabfbe8fc0cfed9fe48ff88ffeeffb700e10127032a04a8049e043b04b7033b03ca025a02f201a30180018901a201a0016c010d01a700680065008e00bb00bf007a00e1fff7fecefd88fc5afb86fa3efa8cfa43fb13fcb9fc22fd85fd43fe9bff79016b03d0042e0578042203da0131014f01ed018802b2025502b3012401e200e100de009900f6ff10ff2cfe81fd24fd0bfd11fd14fd06fdeffce0fcf5fc4cfd06fe28ff8f000502450303041f04b60302035402ed01d901f3010202d1015201a9001400d0ffefff48008a007000efff39ff9efe60fe84fed0fef3feb3fe1bfe6dfdfbfcf5fc4cfdb9fdfbfdeefd9bfd3afd0afd38fde7fd22ffce00b90295040a06dd060507a006ea05180538043603f5017700eafe95fdb8fc5ffc6bfcbffc43fde8fdb3fe97ff71001d017501680111018800d4fff5fedafd85fc36fb45fa00fa8efad2fb76fd21ff9c00e9012d038204df051107ce07f0077d0797066b0510047e02a80094fe75fc9afa4df9aef8aff820f9d3f9abfa9efbb3fcf1fd4dffa900ef010e03eb0365046504e103eb02b8017c0062ff8ffe12fefafd6bfe6fffd30046026003cd03a0033503e202d402fe0208039102820114009ffe67fd88fce2fb42fb9efa1dfafdf961fa37fb4efc5ffd2bfeb3fe23ff94ff2200e800ce01b0027f0321046c045204dd0325034a027601c10019007eff08ffcbfee9fe84ff770071013302900282023d02ef01a2014401a900bbff9cfe93fde7fcaefcbdfcc8fc72fc91fb56fa23f96df8a4f8e5f9f0fb60feb6008c02c5037604cd0408053d057105ab05e305140638062b06b905b004fc02c20066fe5dfc0dfba0faedfa9dfb49fc9bfc7dfc1bfcb4fb86fbbcfb4dfc0ffdd5fd72fecffe01ff1fff42ff93ff2300ec00e201dd02a403220455044d0442045c049804db04ed04a80415045703a20212028001a90058ff78fd43fb2ef99ff7d8f6d2f63ff7d1f755f8d1f894f9edfaf9fc95ff5202ab044806fd06d60625062c051104fe0208022f017f000300b6ff90ff9cfff0ff8b006b018d02ad037404c2048104a80372022601e1ffbdfed2fd13fd68fccdfb3afb9afadef915f961f8ebf7e8f785f8c4f97afb72fd7dff6601f9022804fa046e05a805ed0569062307f00769082708090733050b0303016dff5efeb6fd3efdd8fc86fc51fc3dfc3bfc2efc00fca8fb42fb04fb19fb81fb14fca4fc09fd35fd4afd7dfdf9fde3fe3e00d70183030d052f06c606db068606fb0578051f05ee04d0049f042f045a0318027a0094fe9ffce5fa8af9abf848f830f848f895f805f999f952fa08fbb6fb7bfc66fd93fe300027022704d505de061f07be0601061d05300457039702e8015a01f600a7007500660060006800850087004400a5ff98fe49fd22fc7efb85fb2afc16fdd6fd18fec1fde8fcd1fbdafa49fa45fadcfa05fc9efd77ff4a01d7020904f504b9056606f2063707ff063606000591031b02c70080ff12fe7cfcf0fac0f944f998f990fadbfb07fdcafd36fe85feedfe9eff80003c018b014d01880080ff92fef8fdc1fddbfd2cfea4fe49ff1e000c01f401b2021e033a033b0346036b03b60303040d04ae03d8028701d9ff09fe46fcb5fa73f985f8e0f78ff79bf703f8caf8e6f937fbaafc40fefefff7012b046006370852096c098008c4069a0464026a00dcfec1fd0dfdcdfc0afdb8fdc9fe030000018d01aa016301f0008a003200c0fff7febefd3ffcb4fa6ff9c6f8b5f818f9edf90dfb5afcfcfddcffa601350368041d058305df054106a606eb06cf062d0606058203e5015a00ebfe9bfd68fc53fb79fa05fa1afabdfacffb11fd3efe37ff0600bb0077014402f1023d03f702f601520079fee1fcdbfb95fbf9fbc6fcc0fdcafee7ff27018202d103e4048b05ba059b0560053305340556055d0507052a04a4027f0000fe7cfb3ef9a1f7e1f6f5f6c4f730f9eafaadfc62fedbffe7009001f0011e025402bf024e03d503250403044e033102ff00f9ff5bff53ffd2ffb400e80146039404ba059806fe06d9063106060559034501fcfeb9fccffa8ef908f920f999f911fa40fa38fa2ffa77fa6dfb2efd82ff01021f046e05df059a05f1044104b20356033903380349038a03e8032d042c04b103ab024f01e4ffc3fe44fe8efe8effee002c02dd02bc02c7015e0001ff0cfeb0fdddfd26fe18fe83fd71fc1efb08faabf92cfa73fb33fde8fe2f00fe00880129023d03cf04b806aa083a0a3e0bbd0bac0b050bbb0994078604ee0054fd56fa7ff8eff758f837f915fab4fa19fb76fb06fcdcfcf3fd3cff75006601f60106029d01f20024005effdbfea0fe9dfeedfeb3ff0d01150398051508fe09e10a890a2c094c07740509041c037202b701bb0078ff17fed6fccefbe2fadff9a8f866f785f66cf655f732f9abfb4cfeb700b9023a043605b105bb055905b6041e04bf039703920385034303dd0284025b0289020b039e03080437041d04be034903d60246028401920066ff11fec8fcb2fbdafa43faeaf9c9f9dcf924faabfa6cfb5cfc70fd9afec5fff2002a027903d6042c06680772082b099a09ca09b1095609b5089e0701060004c301a1ffeefdbffcfefb7afbedfa43faa0f93cf94cf9ecf904fb5dfcb4fddbfec9ff83002501c2014b02b102fd02290342037903e0036004e3043d053105ac04d503f7027302a602ac034605f30624086e08a207d8056d03b900f6fd58fbf1f8c7f60df502f4b8f335f467f526f76cf934fc65ffdc023006dd08aa0a950bb60b610bcb0adc098008b806910455026100f0fe16fec8fde2fd58fe41ff9e004102d303ec042d05840434039a0103008dfe28fdb9fb39fac8f8baf75bf7c4f7e8f893fa7bfc70fe51001702e203b7057c071709730a750b0d0c2f0cd40bed0a70097107ff0431025cffcdfcaefa4af9bbf8cbf84af901faa9fa33fbc5fb93fcc5fd4cff0701b402e60370046204ca03e9020b0238017500d0ff3bffc3fe91febefe58ff48006d01c00220048205f506500860090e0a1a0a5a09e407cd053d038800f1fdb4fbe6f97cf869f788f6d9f59af5e8f5e5f6b1f80bfb90fdecffc4010f030904d104a205850635079507710798066705300408034302eb01ba01b901ec015b0229031d04f1045905e304a103da01adffc7fd6bfc35fb5bfa8ef92af8fef6f4f59df4b1f511fa99fd9bfe41ffcdffbeffd6fff8ffdefff0ff0400faff0d000e000500190015000d0017000800ffff0300f0ffe6ffe9ffdfffe9fff9fffbff07000e000a0011000e00020004000100fdff0400050002000300fcfff9fffbfffaffffff020003000c00130014000f000000f7fff4ffebffeffffafff5fff4fff9fff3fff3fff7fff4fff7fffbfffcff0300030004001100160015001f00210019001800110008000600fffffafff8ffeeffe6ffe3ffe1ffe5ffe6ffe4ffeaffeefff5ff06000e000e00130014001000120011000e000c000600faffeeffe5ffe9fff6fffeff01000100ffff020009000f000f0011000f000300f7fff7fffbfffeff05000a000b000b0008000100fcfffafffefffefff8fff7fffcffffff0300050006000c000a00fdfff7fff6fff2fff3fff6fff6fff6fff3fff3fff6fff4fff6fff9fff4fff2fff9ff000006000c000c000d0014001c0020001f001e001d0011000300fefff9fff4fff1ffebffe5ffe4ffe6ffeaffedfff4ff02000b000c00140016000e00;
end
endmodule

//// global definitions 
//`define EOF        -1
//
//// file names 
//`define IN_FILE    "../../../scilab/test_in.bin"
//`define ENC_FILE  "../../../scilab/test_enc.bin"
//`define DEC_FILE  "../../../scilab/test_dec.bin"
//
////---------------------------------------------------------------------------------------
//// test bench implementation 
//// global signals generation  
//initial
//begin
//  clock = 0;
//  rst = 1;
//  #40 rst = 0;
//end 
//
//// clock generator - 50MHz clock 
//always 
//begin 
//  #10 clock = 0;
//  #10 clock = 1;
//end 
//
//// test bench dump variables 
//initial 
//begin 
//  $display("");
//  $display("IMA ADPCM encoder & decoder simulation");
//  $display("--------------------------------------");
//  $dumpfile("test.vcd");
//  $dumpvars(0, test);
//end 
//
////------------------------------------------------------------------
//// encoder input samples read process 
//initial 
//begin 
//  // clear encoder input signal 
//  inSamp = 16'b0;
//  inValid = 1'b0;
//  // clear samples counter 
//  sampCount = 0;
//  
//  // binary input file 
//  infid = $fopen(`IN_FILE, "rb");
//  
//  // wait for reset release
//  while (rst) @(posedge clock);
//  repeat (50) @(posedge clock);
//
//  // read input samples file 
//  intmp = $fgetc(infid);
//  while (intmp != `EOF)
//  begin 
//    // read the next character to form the new input sample 
//    // Note that first byte is used as the low byte of the sample 
//    inSamp[7:0] <= intmp;
//    inSamp[15:8] <= $fgetc(infid);
//    // sign input sample is valid 
//    inValid <= 1'b1;
//    @(posedge clock);
//    
//    // update the sample counter 
//    sampCount = sampCount + 1;
//    
//    // wait for encoder input ready assertion to confirm the new sample was read
//    // by the encoder.
//    while (!inReady)
//      @(posedge clock);
//    
//    // read next character from the input file 
//    intmp = $fgetc(infid);
//  end 
//  // sign input is not valid 
//  inValid <= 1'b0;
//  @(posedge clock);
//  
//  // close input file 
//  $fclose(infid);
//end 
//
//// encoder output checker - the encoder output is compared to the value read from 
//// the ADPCM coded samples file. 
//initial 
//begin 
//  // clear encoded sample value 
//  encCount = 0;
//  // open input file 
//  encfid = $fopen(`ENC_FILE, "rb");
//
//  // wait for reset release
//  while (rst) @(posedge clock);
//    
//  // encoder output compare loop 
//  enctmp = $fgetc(encfid);
//  while (enctmp != `EOF)
//  begin 
//    // assign the expected value to a register with the same width 
//    encExpVal = enctmp;
//    
//    // wait for encoder output valid 
//    while (!encValid)
//      @(posedge clock);
//    
//    // compare the encoded value with the value read from the input file 
//    if (encPcm != encExpVal)
//    begin 
//      // announce error detection and exit simulation 
//      $display(" Error!");
//      $display("Error found in encoder output index %0d.", encCount+1);
//      $display("   (expected value 'h%x, got value 'h%x)", encExpVal, encPcm);
//      // wait for a few clock cycles before ending simulation 
//      repeat (20) @(posedge clock);
//      $finish;
//    end 
//    
//    // update the encoded sample counter 
//    encCount = encCount + 1;
//    // delay for a clock cycle after comparison 
//    @(posedge clock);
//    
//    // read next char from input file 
//    enctmp = $fgetc(encfid);
//  end 
//  
//  // close input file 
//  $fclose(encfid);
//end 
//
//// decoder output checker - the decoder output is compared to the value read from 
//// the ADPCM decoded samples file. 
//initial 
//begin 
//  // clear decoded sample value 
//  decCount = 0;
//  dispCount = 0;
//  // open input file 
//  decfid = $fopen(`DEC_FILE, "rb");
//
//  // wait for reset release
//  while (rst) @(posedge clock);
//
//  // display simulation progress bar title 
//  $write("Simulation progress: ");
//    
//  // decoder output compare loop 
//  dectmp = $fgetc(decfid);
//  while (dectmp != `EOF)
//  begin 
//    // read the next char to form the expected 16 bit sample value 
//    decExpVal[7:0] = dectmp;
//    decExpVal[15:8] = $fgetc(decfid);
//    
//    // wait for decoder output valid 
//    while (!decValid)
//      @(posedge clock);
//    
//    // compare the decoded value with the value read from the input file 
//    if (decSamp != decExpVal)
//    begin 
//      // announce error detection and exit simulation 
//      $display(" Error!");
//      $display("Error found in decoder output index %0d.", decCount+1);
//      $display("   (expected value 'h%x, got value 'h%x)", decExpVal, decSamp);
//      // wait for a few clock cycles before ending simulation 
//      repeat (20) @(posedge clock);
//      $finish;
//    end 
//    // delay for a clock cycle after comparison 
//    @(posedge clock);
//    
//    // update the decoded sample counter 
//    decCount = decCount + 1;
//    
//    // check if simulation progress should be displayed
//    if (dispCount[31:13] != (decCount >> 13))
//      $write(".");
//    // update the display counter 
//    dispCount = decCount;
//    
//    // read next char from input file 
//    dectmp = $fgetc(decfid);
//  end 
//  
//  // close input file 
//  $fclose(decfid);
//  
//  // when decoder output is done announce simulation was successful 
//  $display(" Done");
//  $display("Simulation ended successfully after %0d samples", decCount);
//  $finish;
//end 
//
////------------------------------------------------------------------
//// device under test 
//// Encoder instance 
//ima_adpcm_enc enc
//(
//  .clock(clock), 
//  .reset(rst), 
//  .inSamp(inSamp), 
//  .inValid(inValid),
//  .inReady(inReady),
//  .outPCM(encPcm), 
//  .outValid(encValid), 
//  .outPredictSamp(/* not used */), 
//  .outStepIndex(/* not used */) 
//);
//
//// Decoder instance 
//ima_adpcm_dec dec 
//(
//  .clock(clock), 
//  .reset(rst), 
//  .inPCM(encPcm), 
//  .inValid(encValid),
//  .inReady(decReady),
//  .inPredictSamp(16'b0), 
//  .inStepIndex(7'b0), 
//  .inStateLoad(1'b0), 
//  .outSamp(decSamp), 
//  .outValid(decValid) 
//);
//
//endmodule
////---------------------------------------------------------------------------------------
////            Th.. Th.. Th.. Thats all folks !!!
////---------------------------------------------------------------------------------------
