module read_info_driver #(
  parameter integer NUM_PU = 1,
  parameter integer D_TYPE_W = 2,
  parameter integer RD_SIZE_W = 20
)
(
  input  wire clk,
  input  wire reset,
  input  wire inbuf_pop,
  input  wire read_info_full,
  output reg  inbuf_empty,
  output reg  rd_req,
  output reg  [RD_SIZE_W-1:0]rd_req_size,
  output reg  [PU_ID_W-1:0]rd_req_pu_id,
  output reg  [D_TYPE_W-1:0]rd_req_d_type,
  input  wire [PU_ID_W-1:0] pu_id,
  input  wire               stream_push,
  input  wire               buffer_push,
  output reg                stream_full,
  output reg                buffer_full,
  input  wire [D_TYPE_W-1:0] d_type
);

localparam integer TESTCASES = 500;

localparam integer RANDS = 1000;
localparam integer NEGEDGE_RANDS = RANDS;//1000;  // Number of times the test executes
localparam integer POSEDGE_RANDS = RANDS;//NEGEDGE_RANDS + 1;
localparam integer PU_ID_W = `C_LOG_2(NUM_PU) + 1;
//localparam integer RD_REQ_SIZE_W = `C_LOG_2(10) + 1;
localparam integer RD_REQ_D_TYPE_W = 1;

  integer ctr;
  reg[2:0] state;
  reg counts_equal;
  integer counts_equal_ctr;

  parameter idle = 3'd0;
  parameter start = 3'd1;
  parameter send_reqs_init = 3'd2;
  parameter send_reqs_complete = 3'd3;
  parameter finish = 3'd4;

  integer d_0_count;
  integer d_1_count;

  integer reqs_sent;

  reg pass;
  reg fail;

  test_status #(
    .PREFIX                   ( "RD_INFO"                     ),
    .TIMEOUT                  ( 1000000                  )
  ) status (
    .clk                      ( clk                      ),
    .reset                    ( reset                    ),
    .pass                     ( pass                     ),
    .fail                     ( fail                     )
  );

  integer read_count;
  integer read_info_pop_count;
  integer d0_pop_count;
  integer d1_pop_count;
  integer rd_pointer;
  integer wr_pointer;


  // Arrays of random numbers to replace $urandom and $random system tasks
  reg[RD_SIZE_W - 1:0] rd_req_size_urands[NEGEDGE_RANDS - 1:0];
  reg[31:0] rd_req_pu_id_urands[NEGEDGE_RANDS - 1:0];  // NUM_PU is 1, so can maybe just use 0 always
  reg rd_req_d_type_urands[NEGEDGE_RANDS - 1:0];
  reg inbuf_empty_rands[POSEDGE_RANDS - 1:0];
  reg buffer_full_rands[POSEDGE_RANDS - 1:0];
  reg stream_full_rands[POSEDGE_RANDS - 1:0];

  // Indices into each array
  reg[NEGEDGE_RANDS - 1:0] size_idx;
  reg[NEGEDGE_RANDS - 1:0] pu_id_idx;
  reg[NEGEDGE_RANDS - 1:0] d_type_idx;
  reg[POSEDGE_RANDS - 1:0]  inbuf_empty_idx;
  reg[POSEDGE_RANDS - 1:0]  buffer_full_idx;
  reg[POSEDGE_RANDS - 1:0]  stream_full_idx;

  
  initial begin
    ctr = 0;
    state = start;
    counts_equal = 0;
    counts_equal_ctr = 0;

    pass = 0;
    fail = 0;

    rd_req_size_urands[0]    = 20'd6;
    rd_req_size_urands[1]    = 20'd1;
    rd_req_size_urands[2]    = 20'd9;
    rd_req_size_urands[3]    = 20'd6;
    rd_req_size_urands[4]    = 20'd4;
    rd_req_size_urands[5]    = 20'd8;
    rd_req_size_urands[6]    = 20'd3;
    rd_req_size_urands[7]    = 20'd7;
    rd_req_size_urands[8]    = 20'd3;
    rd_req_size_urands[9]    = 20'd9;
    rd_req_size_urands[10]   = 20'd4;
    rd_req_size_urands[11]   = 20'd2;
    rd_req_size_urands[12]   = 20'd2;
    rd_req_size_urands[13]   = 20'd1;
    rd_req_size_urands[14]   = 20'd9;
    rd_req_size_urands[15]   = 20'd3;
    rd_req_size_urands[16]   = 20'd3;
    rd_req_size_urands[17]   = 20'd5;
    rd_req_size_urands[18]   = 20'd3;
    rd_req_size_urands[19]   = 20'd8;
    rd_req_size_urands[20]   = 20'd1;
    rd_req_size_urands[21]   = 20'd9;
    rd_req_size_urands[22]   = 20'd9;
    rd_req_size_urands[23]   = 20'd10;
    rd_req_size_urands[24]   = 20'd8;
    rd_req_size_urands[25]   = 20'd2;
    rd_req_size_urands[26]   = 20'd10;
    rd_req_size_urands[27]   = 20'd6;
    rd_req_size_urands[28]   = 20'd5;
    rd_req_size_urands[29]   = 20'd10;
    rd_req_size_urands[30]   = 20'd10;
    rd_req_size_urands[31]   = 20'd4;
    rd_req_size_urands[32]   = 20'd1;
    rd_req_size_urands[33]   = 20'd9;
    rd_req_size_urands[34]   = 20'd8;
    rd_req_size_urands[35]   = 20'd2;
    rd_req_size_urands[36]   = 20'd10;
    rd_req_size_urands[37]   = 20'd8;
    rd_req_size_urands[38]   = 20'd8;
    rd_req_size_urands[39]   = 20'd7;
    rd_req_size_urands[40]   = 20'd2;
    rd_req_size_urands[41]   = 20'd4;
    rd_req_size_urands[42]   = 20'd7;
    rd_req_size_urands[43]   = 20'd3;
    rd_req_size_urands[44]   = 20'd7;
    rd_req_size_urands[45]   = 20'd8;
    rd_req_size_urands[46]   = 20'd4;
    rd_req_size_urands[47]   = 20'd6;
    rd_req_size_urands[48]   = 20'd1;
    rd_req_size_urands[49]   = 20'd2;
    rd_req_size_urands[50]   = 20'd7;
    rd_req_size_urands[51]   = 20'd3;
    rd_req_size_urands[52]   = 20'd2;
    rd_req_size_urands[53]   = 20'd2;
    rd_req_size_urands[54]   = 20'd8;
    rd_req_size_urands[55]   = 20'd7;
    rd_req_size_urands[56]   = 20'd9;
    rd_req_size_urands[57]   = 20'd4;
    rd_req_size_urands[58]   = 20'd1;
    rd_req_size_urands[59]   = 20'd1;
    rd_req_size_urands[60]   = 20'd5;
    rd_req_size_urands[61]   = 20'd10;
    rd_req_size_urands[62]   = 20'd5;
    rd_req_size_urands[63]   = 20'd2;
    rd_req_size_urands[64]   = 20'd3;
    rd_req_size_urands[65]   = 20'd5;
    rd_req_size_urands[66]   = 20'd7;
    rd_req_size_urands[67]   = 20'd4;
    rd_req_size_urands[68]   = 20'd10;
    rd_req_size_urands[69]   = 20'd4;
    rd_req_size_urands[70]   = 20'd1;
    rd_req_size_urands[71]   = 20'd1;
    rd_req_size_urands[72]   = 20'd3;
    rd_req_size_urands[73]   = 20'd10;
    rd_req_size_urands[74]   = 20'd4;
    rd_req_size_urands[75]   = 20'd4;
    rd_req_size_urands[76]   = 20'd8;
    rd_req_size_urands[77]   = 20'd2;
    rd_req_size_urands[78]   = 20'd2;
    rd_req_size_urands[79]   = 20'd10;
    rd_req_size_urands[80]   = 20'd5;
    rd_req_size_urands[81]   = 20'd6;
    rd_req_size_urands[82]   = 20'd2;
    rd_req_size_urands[83]   = 20'd5;
    rd_req_size_urands[84]   = 20'd1;
    rd_req_size_urands[85]   = 20'd5;
    rd_req_size_urands[86]   = 20'd9;
    rd_req_size_urands[87]   = 20'd5;
    rd_req_size_urands[88]   = 20'd7;
    rd_req_size_urands[89]   = 20'd10;
    rd_req_size_urands[90]   = 20'd8;
    rd_req_size_urands[91]   = 20'd2;
    rd_req_size_urands[92]   = 20'd5;
    rd_req_size_urands[93]   = 20'd5;
    rd_req_size_urands[94]   = 20'd7;
    rd_req_size_urands[95]   = 20'd10;
    rd_req_size_urands[96]   = 20'd2;
    rd_req_size_urands[97]   = 20'd7;
    rd_req_size_urands[98]   = 20'd1;
    rd_req_size_urands[99]   = 20'd6;
    rd_req_size_urands[100]  = 20'd9;
    rd_req_size_urands[101]  = 20'd7;
    rd_req_size_urands[102]  = 20'd3;
    rd_req_size_urands[103]  = 20'd7;
    rd_req_size_urands[104]  = 20'd6;
    rd_req_size_urands[105]  = 20'd8;
    rd_req_size_urands[106]  = 20'd5;
    rd_req_size_urands[107]  = 20'd5;
    rd_req_size_urands[108]  = 20'd1;
    rd_req_size_urands[109]  = 20'd6;
    rd_req_size_urands[110]  = 20'd4;
    rd_req_size_urands[111]  = 20'd9;
    rd_req_size_urands[112]  = 20'd2;
    rd_req_size_urands[113]  = 20'd8;
    rd_req_size_urands[114]  = 20'd6;
    rd_req_size_urands[115]  = 20'd9;
    rd_req_size_urands[116]  = 20'd7;
    rd_req_size_urands[117]  = 20'd3;
    rd_req_size_urands[118]  = 20'd2;
    rd_req_size_urands[119]  = 20'd10;
    rd_req_size_urands[120]  = 20'd6;
    rd_req_size_urands[121]  = 20'd1;
    rd_req_size_urands[122]  = 20'd5;
    rd_req_size_urands[123]  = 20'd1;
    rd_req_size_urands[124]  = 20'd6;
    rd_req_size_urands[125]  = 20'd6;
    rd_req_size_urands[126]  = 20'd10;
    rd_req_size_urands[127]  = 20'd2;
    rd_req_size_urands[128]  = 20'd4;
    rd_req_size_urands[129]  = 20'd8;
    rd_req_size_urands[130]  = 20'd10;
    rd_req_size_urands[131]  = 20'd1;
    rd_req_size_urands[132]  = 20'd1;
    rd_req_size_urands[133]  = 20'd4;
    rd_req_size_urands[134]  = 20'd4;
    rd_req_size_urands[135]  = 20'd3;
    rd_req_size_urands[136]  = 20'd2;
    rd_req_size_urands[137]  = 20'd6;
    rd_req_size_urands[138]  = 20'd9;
    rd_req_size_urands[139]  = 20'd10;
    rd_req_size_urands[140]  = 20'd7;
    rd_req_size_urands[141]  = 20'd9;
    rd_req_size_urands[142]  = 20'd8;
    rd_req_size_urands[143]  = 20'd10;
    rd_req_size_urands[144]  = 20'd2;
    rd_req_size_urands[145]  = 20'd8;
    rd_req_size_urands[146]  = 20'd9;
    rd_req_size_urands[147]  = 20'd5;
    rd_req_size_urands[148]  = 20'd10;
    rd_req_size_urands[149]  = 20'd9;
    rd_req_size_urands[150]  = 20'd3;
    rd_req_size_urands[151]  = 20'd5;
    rd_req_size_urands[152]  = 20'd10;
    rd_req_size_urands[153]  = 20'd6;
    rd_req_size_urands[154]  = 20'd1;
    rd_req_size_urands[155]  = 20'd9;
    rd_req_size_urands[156]  = 20'd1;
    rd_req_size_urands[157]  = 20'd10;
    rd_req_size_urands[158]  = 20'd7;
    rd_req_size_urands[159]  = 20'd5;
    rd_req_size_urands[160]  = 20'd9;
    rd_req_size_urands[161]  = 20'd2;
    rd_req_size_urands[162]  = 20'd5;
    rd_req_size_urands[163]  = 20'd3;
    rd_req_size_urands[164]  = 20'd1;
    rd_req_size_urands[165]  = 20'd2;
    rd_req_size_urands[166]  = 20'd4;
    rd_req_size_urands[167]  = 20'd5;
    rd_req_size_urands[168]  = 20'd3;
    rd_req_size_urands[169]  = 20'd5;
    rd_req_size_urands[170]  = 20'd2;
    rd_req_size_urands[171]  = 20'd6;
    rd_req_size_urands[172]  = 20'd3;
    rd_req_size_urands[173]  = 20'd2;
    rd_req_size_urands[174]  = 20'd3;
    rd_req_size_urands[175]  = 20'd5;
    rd_req_size_urands[176]  = 20'd10;
    rd_req_size_urands[177]  = 20'd3;
    rd_req_size_urands[178]  = 20'd2;
    rd_req_size_urands[179]  = 20'd10;
    rd_req_size_urands[180]  = 20'd8;
    rd_req_size_urands[181]  = 20'd4;
    rd_req_size_urands[182]  = 20'd10;
    rd_req_size_urands[183]  = 20'd8;
    rd_req_size_urands[184]  = 20'd9;
    rd_req_size_urands[185]  = 20'd6;
    rd_req_size_urands[186]  = 20'd6;
    rd_req_size_urands[187]  = 20'd6;
    rd_req_size_urands[188]  = 20'd9;
    rd_req_size_urands[189]  = 20'd7;
    rd_req_size_urands[190]  = 20'd7;
    rd_req_size_urands[191]  = 20'd4;
    rd_req_size_urands[192]  = 20'd6;
    rd_req_size_urands[193]  = 20'd9;
    rd_req_size_urands[194]  = 20'd5;
    rd_req_size_urands[195]  = 20'd5;
    rd_req_size_urands[196]  = 20'd9;
    rd_req_size_urands[197]  = 20'd6;
    rd_req_size_urands[198]  = 20'd4;
    rd_req_size_urands[199]  = 20'd3;
    rd_req_size_urands[200]  = 20'd9;
    rd_req_size_urands[201]  = 20'd10;
    rd_req_size_urands[202]  = 20'd7;
    rd_req_size_urands[203]  = 20'd5;
    rd_req_size_urands[204]  = 20'd8;
    rd_req_size_urands[205]  = 20'd5;
    rd_req_size_urands[206]  = 20'd1;
    rd_req_size_urands[207]  = 20'd4;
    rd_req_size_urands[208]  = 20'd10;
    rd_req_size_urands[209]  = 20'd5;
    rd_req_size_urands[210]  = 20'd6;
    rd_req_size_urands[211]  = 20'd4;
    rd_req_size_urands[212]  = 20'd7;
    rd_req_size_urands[213]  = 20'd8;
    rd_req_size_urands[214]  = 20'd5;
    rd_req_size_urands[215]  = 20'd1;
    rd_req_size_urands[216]  = 20'd5;
    rd_req_size_urands[217]  = 20'd9;
    rd_req_size_urands[218]  = 20'd5;
    rd_req_size_urands[219]  = 20'd1;
    rd_req_size_urands[220]  = 20'd1;
    rd_req_size_urands[221]  = 20'd2;
    rd_req_size_urands[222]  = 20'd6;
    rd_req_size_urands[223]  = 20'd6;
    rd_req_size_urands[224]  = 20'd10;
    rd_req_size_urands[225]  = 20'd1;
    rd_req_size_urands[226]  = 20'd9;
    rd_req_size_urands[227]  = 20'd9;
    rd_req_size_urands[228]  = 20'd5;
    rd_req_size_urands[229]  = 20'd5;
    rd_req_size_urands[230]  = 20'd3;
    rd_req_size_urands[231]  = 20'd3;
    rd_req_size_urands[232]  = 20'd4;
    rd_req_size_urands[233]  = 20'd9;
    rd_req_size_urands[234]  = 20'd7;
    rd_req_size_urands[235]  = 20'd3;
    rd_req_size_urands[236]  = 20'd1;
    rd_req_size_urands[237]  = 20'd10;
    rd_req_size_urands[238]  = 20'd2;
    rd_req_size_urands[239]  = 20'd2;
    rd_req_size_urands[240]  = 20'd3;
    rd_req_size_urands[241]  = 20'd2;
    rd_req_size_urands[242]  = 20'd5;
    rd_req_size_urands[243]  = 20'd4;
    rd_req_size_urands[244]  = 20'd5;
    rd_req_size_urands[245]  = 20'd10;
    rd_req_size_urands[246]  = 20'd3;
    rd_req_size_urands[247]  = 20'd6;
    rd_req_size_urands[248]  = 20'd4;
    rd_req_size_urands[249]  = 20'd4;
    rd_req_size_urands[250]  = 20'd3;
    rd_req_size_urands[251]  = 20'd10;
    rd_req_size_urands[252]  = 20'd10;
    rd_req_size_urands[253]  = 20'd3;
    rd_req_size_urands[254]  = 20'd3;
    rd_req_size_urands[255]  = 20'd1;
    rd_req_size_urands[256]  = 20'd7;
    rd_req_size_urands[257]  = 20'd10;
    rd_req_size_urands[258]  = 20'd6;
    rd_req_size_urands[259]  = 20'd4;
    rd_req_size_urands[260]  = 20'd3;
    rd_req_size_urands[261]  = 20'd9;
    rd_req_size_urands[262]  = 20'd2;
    rd_req_size_urands[263]  = 20'd4;
    rd_req_size_urands[264]  = 20'd3;
    rd_req_size_urands[265]  = 20'd1;
    rd_req_size_urands[266]  = 20'd8;
    rd_req_size_urands[267]  = 20'd10;
    rd_req_size_urands[268]  = 20'd2;
    rd_req_size_urands[269]  = 20'd4;
    rd_req_size_urands[270]  = 20'd7;
    rd_req_size_urands[271]  = 20'd9;
    rd_req_size_urands[272]  = 20'd1;
    rd_req_size_urands[273]  = 20'd4;
    rd_req_size_urands[274]  = 20'd1;
    rd_req_size_urands[275]  = 20'd7;
    rd_req_size_urands[276]  = 20'd8;
    rd_req_size_urands[277]  = 20'd6;
    rd_req_size_urands[278]  = 20'd2;
    rd_req_size_urands[279]  = 20'd1;
    rd_req_size_urands[280]  = 20'd2;
    rd_req_size_urands[281]  = 20'd1;
    rd_req_size_urands[282]  = 20'd7;
    rd_req_size_urands[283]  = 20'd2;
    rd_req_size_urands[284]  = 20'd3;
    rd_req_size_urands[285]  = 20'd8;
    rd_req_size_urands[286]  = 20'd10;
    rd_req_size_urands[287]  = 20'd5;
    rd_req_size_urands[288]  = 20'd5;
    rd_req_size_urands[289]  = 20'd7;
    rd_req_size_urands[290]  = 20'd3;
    rd_req_size_urands[291]  = 20'd3;
    rd_req_size_urands[292]  = 20'd7;
    rd_req_size_urands[293]  = 20'd6;
    rd_req_size_urands[294]  = 20'd9;
    rd_req_size_urands[295]  = 20'd9;
    rd_req_size_urands[296]  = 20'd10;
    rd_req_size_urands[297]  = 20'd8;
    rd_req_size_urands[298]  = 20'd10;
    rd_req_size_urands[299]  = 20'd7;
    rd_req_size_urands[300]  = 20'd4;
    rd_req_size_urands[301]  = 20'd1;
    rd_req_size_urands[302]  = 20'd10;
    rd_req_size_urands[303]  = 20'd5;
    rd_req_size_urands[304]  = 20'd1;
    rd_req_size_urands[305]  = 20'd1;
    rd_req_size_urands[306]  = 20'd2;
    rd_req_size_urands[307]  = 20'd6;
    rd_req_size_urands[308]  = 20'd2;
    rd_req_size_urands[309]  = 20'd4;
    rd_req_size_urands[310]  = 20'd4;
    rd_req_size_urands[311]  = 20'd10;
    rd_req_size_urands[312]  = 20'd8;
    rd_req_size_urands[313]  = 20'd4;
    rd_req_size_urands[314]  = 20'd10;
    rd_req_size_urands[315]  = 20'd6;
    rd_req_size_urands[316]  = 20'd7;
    rd_req_size_urands[317]  = 20'd5;
    rd_req_size_urands[318]  = 20'd4;
    rd_req_size_urands[319]  = 20'd3;
    rd_req_size_urands[320]  = 20'd3;
    rd_req_size_urands[321]  = 20'd2;
    rd_req_size_urands[322]  = 20'd1;
    rd_req_size_urands[323]  = 20'd2;
    rd_req_size_urands[324]  = 20'd5;
    rd_req_size_urands[325]  = 20'd1;
    rd_req_size_urands[326]  = 20'd7;
    rd_req_size_urands[327]  = 20'd6;
    rd_req_size_urands[328]  = 20'd8;
    rd_req_size_urands[329]  = 20'd9;
    rd_req_size_urands[330]  = 20'd9;
    rd_req_size_urands[331]  = 20'd6;
    rd_req_size_urands[332]  = 20'd2;
    rd_req_size_urands[333]  = 20'd8;
    rd_req_size_urands[334]  = 20'd2;
    rd_req_size_urands[335]  = 20'd5;
    rd_req_size_urands[336]  = 20'd2;
    rd_req_size_urands[337]  = 20'd9;
    rd_req_size_urands[338]  = 20'd3;
    rd_req_size_urands[339]  = 20'd1;
    rd_req_size_urands[340]  = 20'd2;
    rd_req_size_urands[341]  = 20'd5;
    rd_req_size_urands[342]  = 20'd8;
    rd_req_size_urands[343]  = 20'd8;
    rd_req_size_urands[344]  = 20'd3;
    rd_req_size_urands[345]  = 20'd3;
    rd_req_size_urands[346]  = 20'd3;
    rd_req_size_urands[347]  = 20'd1;
    rd_req_size_urands[348]  = 20'd7;
    rd_req_size_urands[349]  = 20'd8;
    rd_req_size_urands[350]  = 20'd8;
    rd_req_size_urands[351]  = 20'd6;
    rd_req_size_urands[352]  = 20'd6;
    rd_req_size_urands[353]  = 20'd1;
    rd_req_size_urands[354]  = 20'd4;
    rd_req_size_urands[355]  = 20'd10;
    rd_req_size_urands[356]  = 20'd4;
    rd_req_size_urands[357]  = 20'd9;
    rd_req_size_urands[358]  = 20'd9;
    rd_req_size_urands[359]  = 20'd1;
    rd_req_size_urands[360]  = 20'd10;
    rd_req_size_urands[361]  = 20'd3;
    rd_req_size_urands[362]  = 20'd4;
    rd_req_size_urands[363]  = 20'd2;
    rd_req_size_urands[364]  = 20'd1;
    rd_req_size_urands[365]  = 20'd10;
    rd_req_size_urands[366]  = 20'd10;
    rd_req_size_urands[367]  = 20'd6;
    rd_req_size_urands[368]  = 20'd3;
    rd_req_size_urands[369]  = 20'd9;
    rd_req_size_urands[370]  = 20'd9;
    rd_req_size_urands[371]  = 20'd9;
    rd_req_size_urands[372]  = 20'd3;
    rd_req_size_urands[373]  = 20'd8;
    rd_req_size_urands[374]  = 20'd5;
    rd_req_size_urands[375]  = 20'd1;
    rd_req_size_urands[376]  = 20'd8;
    rd_req_size_urands[377]  = 20'd3;
    rd_req_size_urands[378]  = 20'd8;
    rd_req_size_urands[379]  = 20'd1;
    rd_req_size_urands[380]  = 20'd1;
    rd_req_size_urands[381]  = 20'd5;
    rd_req_size_urands[382]  = 20'd7;
    rd_req_size_urands[383]  = 20'd5;
    rd_req_size_urands[384]  = 20'd7;
    rd_req_size_urands[385]  = 20'd10;
    rd_req_size_urands[386]  = 20'd3;
    rd_req_size_urands[387]  = 20'd6;
    rd_req_size_urands[388]  = 20'd7;
    rd_req_size_urands[389]  = 20'd5;
    rd_req_size_urands[390]  = 20'd9;
    rd_req_size_urands[391]  = 20'd2;
    rd_req_size_urands[392]  = 20'd2;
    rd_req_size_urands[393]  = 20'd9;
    rd_req_size_urands[394]  = 20'd8;
    rd_req_size_urands[395]  = 20'd1;
    rd_req_size_urands[396]  = 20'd10;
    rd_req_size_urands[397]  = 20'd10;
    rd_req_size_urands[398]  = 20'd7;
    rd_req_size_urands[399]  = 20'd6;
    rd_req_size_urands[400]  = 20'd1;
    rd_req_size_urands[401]  = 20'd5;
    rd_req_size_urands[402]  = 20'd10;
    rd_req_size_urands[403]  = 20'd5;
    rd_req_size_urands[404]  = 20'd6;
    rd_req_size_urands[405]  = 20'd6;
    rd_req_size_urands[406]  = 20'd4;
    rd_req_size_urands[407]  = 20'd3;
    rd_req_size_urands[408]  = 20'd8;
    rd_req_size_urands[409]  = 20'd8;
    rd_req_size_urands[410]  = 20'd10;
    rd_req_size_urands[411]  = 20'd5;
    rd_req_size_urands[412]  = 20'd5;
    rd_req_size_urands[413]  = 20'd3;
    rd_req_size_urands[414]  = 20'd4;
    rd_req_size_urands[415]  = 20'd9;
    rd_req_size_urands[416]  = 20'd7;
    rd_req_size_urands[417]  = 20'd2;
    rd_req_size_urands[418]  = 20'd10;
    rd_req_size_urands[419]  = 20'd5;
    rd_req_size_urands[420]  = 20'd7;
    rd_req_size_urands[421]  = 20'd2;
    rd_req_size_urands[422]  = 20'd8;
    rd_req_size_urands[423]  = 20'd2;
    rd_req_size_urands[424]  = 20'd1;
    rd_req_size_urands[425]  = 20'd2;
    rd_req_size_urands[426]  = 20'd5;
    rd_req_size_urands[427]  = 20'd8;
    rd_req_size_urands[428]  = 20'd5;
    rd_req_size_urands[429]  = 20'd6;
    rd_req_size_urands[430]  = 20'd9;
    rd_req_size_urands[431]  = 20'd9;
    rd_req_size_urands[432]  = 20'd3;
    rd_req_size_urands[433]  = 20'd6;
    rd_req_size_urands[434]  = 20'd3;
    rd_req_size_urands[435]  = 20'd5;
    rd_req_size_urands[436]  = 20'd1;
    rd_req_size_urands[437]  = 20'd10;
    rd_req_size_urands[438]  = 20'd4;
    rd_req_size_urands[439]  = 20'd1;
    rd_req_size_urands[440]  = 20'd9;
    rd_req_size_urands[441]  = 20'd10;
    rd_req_size_urands[442]  = 20'd4;
    rd_req_size_urands[443]  = 20'd8;
    rd_req_size_urands[444]  = 20'd1;
    rd_req_size_urands[445]  = 20'd9;
    rd_req_size_urands[446]  = 20'd9;
    rd_req_size_urands[447]  = 20'd9;
    rd_req_size_urands[448]  = 20'd6;
    rd_req_size_urands[449]  = 20'd1;
    rd_req_size_urands[450]  = 20'd6;
    rd_req_size_urands[451]  = 20'd9;
    rd_req_size_urands[452]  = 20'd7;
    rd_req_size_urands[453]  = 20'd9;
    rd_req_size_urands[454]  = 20'd2;
    rd_req_size_urands[455]  = 20'd7;
    rd_req_size_urands[456]  = 20'd6;
    rd_req_size_urands[457]  = 20'd7;
    rd_req_size_urands[458]  = 20'd1;
    rd_req_size_urands[459]  = 20'd2;
    rd_req_size_urands[460]  = 20'd6;
    rd_req_size_urands[461]  = 20'd4;
    rd_req_size_urands[462]  = 20'd6;
    rd_req_size_urands[463]  = 20'd8;
    rd_req_size_urands[464]  = 20'd7;
    rd_req_size_urands[465]  = 20'd1;
    rd_req_size_urands[466]  = 20'd10;
    rd_req_size_urands[467]  = 20'd9;
    rd_req_size_urands[468]  = 20'd10;
    rd_req_size_urands[469]  = 20'd1;
    rd_req_size_urands[470]  = 20'd7;
    rd_req_size_urands[471]  = 20'd7;
    rd_req_size_urands[472]  = 20'd5;
    rd_req_size_urands[473]  = 20'd6;
    rd_req_size_urands[474]  = 20'd3;
    rd_req_size_urands[475]  = 20'd10;
    rd_req_size_urands[476]  = 20'd7;
    rd_req_size_urands[477]  = 20'd10;
    rd_req_size_urands[478]  = 20'd6;
    rd_req_size_urands[479]  = 20'd8;
    rd_req_size_urands[480]  = 20'd2;
    rd_req_size_urands[481]  = 20'd5;
    rd_req_size_urands[482]  = 20'd7;
    rd_req_size_urands[483]  = 20'd7;
    rd_req_size_urands[484]  = 20'd3;
    rd_req_size_urands[485]  = 20'd3;
    rd_req_size_urands[486]  = 20'd3;
    rd_req_size_urands[487]  = 20'd6;
    rd_req_size_urands[488]  = 20'd1;
    rd_req_size_urands[489]  = 20'd2;
    rd_req_size_urands[490]  = 20'd1;
    rd_req_size_urands[491]  = 20'd7;
    rd_req_size_urands[492]  = 20'd4;
    rd_req_size_urands[493]  = 20'd10;
    rd_req_size_urands[494]  = 20'd3;
    rd_req_size_urands[495]  = 20'd10;
    rd_req_size_urands[496]  = 20'd7;
    rd_req_size_urands[497]  = 20'd8;
    rd_req_size_urands[498]  = 20'd8;
    rd_req_size_urands[499]  = 20'd7;
    rd_req_size_urands[500]  = 20'd10;
    rd_req_size_urands[501]  = 20'd3;
    rd_req_size_urands[502]  = 20'd3;
    rd_req_size_urands[503]  = 20'd8;
    rd_req_size_urands[504]  = 20'd3;
    rd_req_size_urands[505]  = 20'd6;
    rd_req_size_urands[506]  = 20'd7;
    rd_req_size_urands[507]  = 20'd10;
    rd_req_size_urands[508]  = 20'd4;
    rd_req_size_urands[509]  = 20'd5;
    rd_req_size_urands[510]  = 20'd6;
    rd_req_size_urands[511]  = 20'd4;
    rd_req_size_urands[512]  = 20'd5;
    rd_req_size_urands[513]  = 20'd4;
    rd_req_size_urands[514]  = 20'd2;
    rd_req_size_urands[515]  = 20'd4;
    rd_req_size_urands[516]  = 20'd9;
    rd_req_size_urands[517]  = 20'd3;
    rd_req_size_urands[518]  = 20'd9;
    rd_req_size_urands[519]  = 20'd9;
    rd_req_size_urands[520]  = 20'd6;
    rd_req_size_urands[521]  = 20'd1;
    rd_req_size_urands[522]  = 20'd8;
    rd_req_size_urands[523]  = 20'd7;
    rd_req_size_urands[524]  = 20'd3;
    rd_req_size_urands[525]  = 20'd1;
    rd_req_size_urands[526]  = 20'd10;
    rd_req_size_urands[527]  = 20'd8;
    rd_req_size_urands[528]  = 20'd2;
    rd_req_size_urands[529]  = 20'd9;
    rd_req_size_urands[530]  = 20'd10;
    rd_req_size_urands[531]  = 20'd10;
    rd_req_size_urands[532]  = 20'd5;
    rd_req_size_urands[533]  = 20'd10;
    rd_req_size_urands[534]  = 20'd2;
    rd_req_size_urands[535]  = 20'd2;
    rd_req_size_urands[536]  = 20'd1;
    rd_req_size_urands[537]  = 20'd10;
    rd_req_size_urands[538]  = 20'd3;
    rd_req_size_urands[539]  = 20'd8;
    rd_req_size_urands[540]  = 20'd10;
    rd_req_size_urands[541]  = 20'd1;
    rd_req_size_urands[542]  = 20'd10;
    rd_req_size_urands[543]  = 20'd7;
    rd_req_size_urands[544]  = 20'd1;
    rd_req_size_urands[545]  = 20'd8;
    rd_req_size_urands[546]  = 20'd10;
    rd_req_size_urands[547]  = 20'd9;
    rd_req_size_urands[548]  = 20'd2;
    rd_req_size_urands[549]  = 20'd7;
    rd_req_size_urands[550]  = 20'd3;
    rd_req_size_urands[551]  = 20'd5;
    rd_req_size_urands[552]  = 20'd9;
    rd_req_size_urands[553]  = 20'd1;
    rd_req_size_urands[554]  = 20'd2;
    rd_req_size_urands[555]  = 20'd1;
    rd_req_size_urands[556]  = 20'd9;
    rd_req_size_urands[557]  = 20'd1;
    rd_req_size_urands[558]  = 20'd5;
    rd_req_size_urands[559]  = 20'd6;
    rd_req_size_urands[560]  = 20'd1;
    rd_req_size_urands[561]  = 20'd1;
    rd_req_size_urands[562]  = 20'd6;
    rd_req_size_urands[563]  = 20'd8;
    rd_req_size_urands[564]  = 20'd7;
    rd_req_size_urands[565]  = 20'd2;
    rd_req_size_urands[566]  = 20'd5;
    rd_req_size_urands[567]  = 20'd3;
    rd_req_size_urands[568]  = 20'd7;
    rd_req_size_urands[569]  = 20'd5;
    rd_req_size_urands[570]  = 20'd1;
    rd_req_size_urands[571]  = 20'd5;
    rd_req_size_urands[572]  = 20'd3;
    rd_req_size_urands[573]  = 20'd6;
    rd_req_size_urands[574]  = 20'd9;
    rd_req_size_urands[575]  = 20'd3;
    rd_req_size_urands[576]  = 20'd5;
    rd_req_size_urands[577]  = 20'd8;
    rd_req_size_urands[578]  = 20'd6;
    rd_req_size_urands[579]  = 20'd5;
    rd_req_size_urands[580]  = 20'd2;
    rd_req_size_urands[581]  = 20'd7;
    rd_req_size_urands[582]  = 20'd1;
    rd_req_size_urands[583]  = 20'd10;
    rd_req_size_urands[584]  = 20'd1;
    rd_req_size_urands[585]  = 20'd8;
    rd_req_size_urands[586]  = 20'd9;
    rd_req_size_urands[587]  = 20'd8;
    rd_req_size_urands[588]  = 20'd3;
    rd_req_size_urands[589]  = 20'd7;
    rd_req_size_urands[590]  = 20'd5;
    rd_req_size_urands[591]  = 20'd9;
    rd_req_size_urands[592]  = 20'd8;
    rd_req_size_urands[593]  = 20'd10;
    rd_req_size_urands[594]  = 20'd3;
    rd_req_size_urands[595]  = 20'd3;
    rd_req_size_urands[596]  = 20'd8;
    rd_req_size_urands[597]  = 20'd5;
    rd_req_size_urands[598]  = 20'd10;
    rd_req_size_urands[599]  = 20'd9;
    rd_req_size_urands[600]  = 20'd7;
    rd_req_size_urands[601]  = 20'd2;
    rd_req_size_urands[602]  = 20'd7;
    rd_req_size_urands[603]  = 20'd7;
    rd_req_size_urands[604]  = 20'd5;
    rd_req_size_urands[605]  = 20'd7;
    rd_req_size_urands[606]  = 20'd7;
    rd_req_size_urands[607]  = 20'd10;
    rd_req_size_urands[608]  = 20'd7;
    rd_req_size_urands[609]  = 20'd1;
    rd_req_size_urands[610]  = 20'd2;
    rd_req_size_urands[611]  = 20'd6;
    rd_req_size_urands[612]  = 20'd9;
    rd_req_size_urands[613]  = 20'd2;
    rd_req_size_urands[614]  = 20'd2;
    rd_req_size_urands[615]  = 20'd10;
    rd_req_size_urands[616]  = 20'd1;
    rd_req_size_urands[617]  = 20'd3;
    rd_req_size_urands[618]  = 20'd2;
    rd_req_size_urands[619]  = 20'd10;
    rd_req_size_urands[620]  = 20'd8;
    rd_req_size_urands[621]  = 20'd3;
    rd_req_size_urands[622]  = 20'd4;
    rd_req_size_urands[623]  = 20'd5;
    rd_req_size_urands[624]  = 20'd1;
    rd_req_size_urands[625]  = 20'd4;
    rd_req_size_urands[626]  = 20'd6;
    rd_req_size_urands[627]  = 20'd8;
    rd_req_size_urands[628]  = 20'd1;
    rd_req_size_urands[629]  = 20'd3;
    rd_req_size_urands[630]  = 20'd5;
    rd_req_size_urands[631]  = 20'd7;
    rd_req_size_urands[632]  = 20'd7;
    rd_req_size_urands[633]  = 20'd7;
    rd_req_size_urands[634]  = 20'd1;
    rd_req_size_urands[635]  = 20'd10;
    rd_req_size_urands[636]  = 20'd5;
    rd_req_size_urands[637]  = 20'd8;
    rd_req_size_urands[638]  = 20'd2;
    rd_req_size_urands[639]  = 20'd1;
    rd_req_size_urands[640]  = 20'd1;
    rd_req_size_urands[641]  = 20'd3;
    rd_req_size_urands[642]  = 20'd5;
    rd_req_size_urands[643]  = 20'd1;
    rd_req_size_urands[644]  = 20'd3;
    rd_req_size_urands[645]  = 20'd2;
    rd_req_size_urands[646]  = 20'd9;
    rd_req_size_urands[647]  = 20'd1;
    rd_req_size_urands[648]  = 20'd6;
    rd_req_size_urands[649]  = 20'd7;
    rd_req_size_urands[650]  = 20'd7;
    rd_req_size_urands[651]  = 20'd6;
    rd_req_size_urands[652]  = 20'd4;
    rd_req_size_urands[653]  = 20'd3;
    rd_req_size_urands[654]  = 20'd2;
    rd_req_size_urands[655]  = 20'd10;
    rd_req_size_urands[656]  = 20'd7;
    rd_req_size_urands[657]  = 20'd8;
    rd_req_size_urands[658]  = 20'd3;
    rd_req_size_urands[659]  = 20'd1;
    rd_req_size_urands[660]  = 20'd6;
    rd_req_size_urands[661]  = 20'd4;
    rd_req_size_urands[662]  = 20'd10;
    rd_req_size_urands[663]  = 20'd6;
    rd_req_size_urands[664]  = 20'd1;
    rd_req_size_urands[665]  = 20'd6;
    rd_req_size_urands[666]  = 20'd10;
    rd_req_size_urands[667]  = 20'd10;
    rd_req_size_urands[668]  = 20'd1;
    rd_req_size_urands[669]  = 20'd6;
    rd_req_size_urands[670]  = 20'd4;
    rd_req_size_urands[671]  = 20'd6;
    rd_req_size_urands[672]  = 20'd7;
    rd_req_size_urands[673]  = 20'd2;
    rd_req_size_urands[674]  = 20'd10;
    rd_req_size_urands[675]  = 20'd2;
    rd_req_size_urands[676]  = 20'd2;
    rd_req_size_urands[677]  = 20'd2;
    rd_req_size_urands[678]  = 20'd6;
    rd_req_size_urands[679]  = 20'd1;
    rd_req_size_urands[680]  = 20'd5;
    rd_req_size_urands[681]  = 20'd2;
    rd_req_size_urands[682]  = 20'd1;
    rd_req_size_urands[683]  = 20'd4;
    rd_req_size_urands[684]  = 20'd2;
    rd_req_size_urands[685]  = 20'd7;
    rd_req_size_urands[686]  = 20'd4;
    rd_req_size_urands[687]  = 20'd8;
    rd_req_size_urands[688]  = 20'd4;
    rd_req_size_urands[689]  = 20'd1;
    rd_req_size_urands[690]  = 20'd4;
    rd_req_size_urands[691]  = 20'd1;
    rd_req_size_urands[692]  = 20'd1;
    rd_req_size_urands[693]  = 20'd2;
    rd_req_size_urands[694]  = 20'd6;
    rd_req_size_urands[695]  = 20'd1;
    rd_req_size_urands[696]  = 20'd10;
    rd_req_size_urands[697]  = 20'd7;
    rd_req_size_urands[698]  = 20'd10;
    rd_req_size_urands[699]  = 20'd3;
    rd_req_size_urands[700]  = 20'd5;
    rd_req_size_urands[701]  = 20'd8;
    rd_req_size_urands[702]  = 20'd1;
    rd_req_size_urands[703]  = 20'd5;
    rd_req_size_urands[704]  = 20'd5;
    rd_req_size_urands[705]  = 20'd9;
    rd_req_size_urands[706]  = 20'd9;
    rd_req_size_urands[707]  = 20'd5;
    rd_req_size_urands[708]  = 20'd10;
    rd_req_size_urands[709]  = 20'd7;
    rd_req_size_urands[710]  = 20'd8;
    rd_req_size_urands[711]  = 20'd5;
    rd_req_size_urands[712]  = 20'd4;
    rd_req_size_urands[713]  = 20'd4;
    rd_req_size_urands[714]  = 20'd9;
    rd_req_size_urands[715]  = 20'd6;
    rd_req_size_urands[716]  = 20'd2;
    rd_req_size_urands[717]  = 20'd9;
    rd_req_size_urands[718]  = 20'd6;
    rd_req_size_urands[719]  = 20'd6;
    rd_req_size_urands[720]  = 20'd3;
    rd_req_size_urands[721]  = 20'd7;
    rd_req_size_urands[722]  = 20'd9;
    rd_req_size_urands[723]  = 20'd10;
    rd_req_size_urands[724]  = 20'd7;
    rd_req_size_urands[725]  = 20'd10;
    rd_req_size_urands[726]  = 20'd4;
    rd_req_size_urands[727]  = 20'd1;
    rd_req_size_urands[728]  = 20'd1;
    rd_req_size_urands[729]  = 20'd5;
    rd_req_size_urands[730]  = 20'd9;
    rd_req_size_urands[731]  = 20'd1;
    rd_req_size_urands[732]  = 20'd7;
    rd_req_size_urands[733]  = 20'd1;
    rd_req_size_urands[734]  = 20'd9;
    rd_req_size_urands[735]  = 20'd3;
    rd_req_size_urands[736]  = 20'd6;
    rd_req_size_urands[737]  = 20'd9;
    rd_req_size_urands[738]  = 20'd10;
    rd_req_size_urands[739]  = 20'd10;
    rd_req_size_urands[740]  = 20'd10;
    rd_req_size_urands[741]  = 20'd6;
    rd_req_size_urands[742]  = 20'd3;
    rd_req_size_urands[743]  = 20'd8;
    rd_req_size_urands[744]  = 20'd4;
    rd_req_size_urands[745]  = 20'd1;
    rd_req_size_urands[746]  = 20'd7;
    rd_req_size_urands[747]  = 20'd4;
    rd_req_size_urands[748]  = 20'd10;
    rd_req_size_urands[749]  = 20'd2;
    rd_req_size_urands[750]  = 20'd7;
    rd_req_size_urands[751]  = 20'd2;
    rd_req_size_urands[752]  = 20'd2;
    rd_req_size_urands[753]  = 20'd7;
    rd_req_size_urands[754]  = 20'd2;
    rd_req_size_urands[755]  = 20'd6;
    rd_req_size_urands[756]  = 20'd9;
    rd_req_size_urands[757]  = 20'd9;
    rd_req_size_urands[758]  = 20'd1;
    rd_req_size_urands[759]  = 20'd4;
    rd_req_size_urands[760]  = 20'd3;
    rd_req_size_urands[761]  = 20'd10;
    rd_req_size_urands[762]  = 20'd4;
    rd_req_size_urands[763]  = 20'd1;
    rd_req_size_urands[764]  = 20'd8;
    rd_req_size_urands[765]  = 20'd3;
    rd_req_size_urands[766]  = 20'd5;
    rd_req_size_urands[767]  = 20'd5;
    rd_req_size_urands[768]  = 20'd10;
    rd_req_size_urands[769]  = 20'd6;
    rd_req_size_urands[770]  = 20'd2;
    rd_req_size_urands[771]  = 20'd10;
    rd_req_size_urands[772]  = 20'd10;
    rd_req_size_urands[773]  = 20'd2;
    rd_req_size_urands[774]  = 20'd2;
    rd_req_size_urands[775]  = 20'd1;
    rd_req_size_urands[776]  = 20'd2;
    rd_req_size_urands[777]  = 20'd8;
    rd_req_size_urands[778]  = 20'd2;
    rd_req_size_urands[779]  = 20'd1;
    rd_req_size_urands[780]  = 20'd2;
    rd_req_size_urands[781]  = 20'd5;
    rd_req_size_urands[782]  = 20'd6;
    rd_req_size_urands[783]  = 20'd1;
    rd_req_size_urands[784]  = 20'd2;
    rd_req_size_urands[785]  = 20'd4;
    rd_req_size_urands[786]  = 20'd3;
    rd_req_size_urands[787]  = 20'd1;
    rd_req_size_urands[788]  = 20'd7;
    rd_req_size_urands[789]  = 20'd9;
    rd_req_size_urands[790]  = 20'd4;
    rd_req_size_urands[791]  = 20'd7;
    rd_req_size_urands[792]  = 20'd5;
    rd_req_size_urands[793]  = 20'd10;
    rd_req_size_urands[794]  = 20'd4;
    rd_req_size_urands[795]  = 20'd10;
    rd_req_size_urands[796]  = 20'd4;
    rd_req_size_urands[797]  = 20'd7;
    rd_req_size_urands[798]  = 20'd6;
    rd_req_size_urands[799]  = 20'd4;
    rd_req_size_urands[800]  = 20'd7;
    rd_req_size_urands[801]  = 20'd10;
    rd_req_size_urands[802]  = 20'd8;
    rd_req_size_urands[803]  = 20'd7;
    rd_req_size_urands[804]  = 20'd5;
    rd_req_size_urands[805]  = 20'd4;
    rd_req_size_urands[806]  = 20'd6;
    rd_req_size_urands[807]  = 20'd5;
    rd_req_size_urands[808]  = 20'd6;
    rd_req_size_urands[809]  = 20'd9;
    rd_req_size_urands[810]  = 20'd4;
    rd_req_size_urands[811]  = 20'd3;
    rd_req_size_urands[812]  = 20'd10;
    rd_req_size_urands[813]  = 20'd8;
    rd_req_size_urands[814]  = 20'd8;
    rd_req_size_urands[815]  = 20'd4;
    rd_req_size_urands[816]  = 20'd4;
    rd_req_size_urands[817]  = 20'd2;
    rd_req_size_urands[818]  = 20'd2;
    rd_req_size_urands[819]  = 20'd1;
    rd_req_size_urands[820]  = 20'd3;
    rd_req_size_urands[821]  = 20'd8;
    rd_req_size_urands[822]  = 20'd8;
    rd_req_size_urands[823]  = 20'd5;
    rd_req_size_urands[824]  = 20'd1;
    rd_req_size_urands[825]  = 20'd2;
    rd_req_size_urands[826]  = 20'd6;
    rd_req_size_urands[827]  = 20'd10;
    rd_req_size_urands[828]  = 20'd6;
    rd_req_size_urands[829]  = 20'd4;
    rd_req_size_urands[830]  = 20'd1;
    rd_req_size_urands[831]  = 20'd5;
    rd_req_size_urands[832]  = 20'd3;
    rd_req_size_urands[833]  = 20'd3;
    rd_req_size_urands[834]  = 20'd7;
    rd_req_size_urands[835]  = 20'd7;
    rd_req_size_urands[836]  = 20'd2;
    rd_req_size_urands[837]  = 20'd10;
    rd_req_size_urands[838]  = 20'd5;
    rd_req_size_urands[839]  = 20'd5;
    rd_req_size_urands[840]  = 20'd8;
    rd_req_size_urands[841]  = 20'd2;
    rd_req_size_urands[842]  = 20'd10;
    rd_req_size_urands[843]  = 20'd3;
    rd_req_size_urands[844]  = 20'd9;
    rd_req_size_urands[845]  = 20'd5;
    rd_req_size_urands[846]  = 20'd10;
    rd_req_size_urands[847]  = 20'd3;
    rd_req_size_urands[848]  = 20'd1;
    rd_req_size_urands[849]  = 20'd10;
    rd_req_size_urands[850]  = 20'd2;
    rd_req_size_urands[851]  = 20'd3;
    rd_req_size_urands[852]  = 20'd8;
    rd_req_size_urands[853]  = 20'd10;
    rd_req_size_urands[854]  = 20'd10;
    rd_req_size_urands[855]  = 20'd8;
    rd_req_size_urands[856]  = 20'd2;
    rd_req_size_urands[857]  = 20'd6;
    rd_req_size_urands[858]  = 20'd1;
    rd_req_size_urands[859]  = 20'd1;
    rd_req_size_urands[860]  = 20'd10;
    rd_req_size_urands[861]  = 20'd1;
    rd_req_size_urands[862]  = 20'd2;
    rd_req_size_urands[863]  = 20'd1;
    rd_req_size_urands[864]  = 20'd2;
    rd_req_size_urands[865]  = 20'd3;
    rd_req_size_urands[866]  = 20'd4;
    rd_req_size_urands[867]  = 20'd3;
    rd_req_size_urands[868]  = 20'd1;
    rd_req_size_urands[869]  = 20'd4;
    rd_req_size_urands[870]  = 20'd7;
    rd_req_size_urands[871]  = 20'd7;
    rd_req_size_urands[872]  = 20'd7;
    rd_req_size_urands[873]  = 20'd10;
    rd_req_size_urands[874]  = 20'd7;
    rd_req_size_urands[875]  = 20'd6;
    rd_req_size_urands[876]  = 20'd4;
    rd_req_size_urands[877]  = 20'd9;
    rd_req_size_urands[878]  = 20'd1;
    rd_req_size_urands[879]  = 20'd6;
    rd_req_size_urands[880]  = 20'd10;
    rd_req_size_urands[881]  = 20'd6;
    rd_req_size_urands[882]  = 20'd1;
    rd_req_size_urands[883]  = 20'd9;
    rd_req_size_urands[884]  = 20'd7;
    rd_req_size_urands[885]  = 20'd7;
    rd_req_size_urands[886]  = 20'd5;
    rd_req_size_urands[887]  = 20'd8;
    rd_req_size_urands[888]  = 20'd6;
    rd_req_size_urands[889]  = 20'd1;
    rd_req_size_urands[890]  = 20'd8;
    rd_req_size_urands[891]  = 20'd5;
    rd_req_size_urands[892]  = 20'd2;
    rd_req_size_urands[893]  = 20'd4;
    rd_req_size_urands[894]  = 20'd7;
    rd_req_size_urands[895]  = 20'd9;
    rd_req_size_urands[896]  = 20'd3;
    rd_req_size_urands[897]  = 20'd9;
    rd_req_size_urands[898]  = 20'd8;
    rd_req_size_urands[899]  = 20'd5;
    rd_req_size_urands[900]  = 20'd2;
    rd_req_size_urands[901]  = 20'd6;
    rd_req_size_urands[902]  = 20'd8;
    rd_req_size_urands[903]  = 20'd8;
    rd_req_size_urands[904]  = 20'd3;
    rd_req_size_urands[905]  = 20'd2;
    rd_req_size_urands[906]  = 20'd6;
    rd_req_size_urands[907]  = 20'd1;
    rd_req_size_urands[908]  = 20'd10;
    rd_req_size_urands[909]  = 20'd7;
    rd_req_size_urands[910]  = 20'd6;
    rd_req_size_urands[911]  = 20'd7;
    rd_req_size_urands[912]  = 20'd8;
    rd_req_size_urands[913]  = 20'd5;
    rd_req_size_urands[914]  = 20'd7;
    rd_req_size_urands[915]  = 20'd6;
    rd_req_size_urands[916]  = 20'd10;
    rd_req_size_urands[917]  = 20'd6;
    rd_req_size_urands[918]  = 20'd7;
    rd_req_size_urands[919]  = 20'd2;
    rd_req_size_urands[920]  = 20'd6;
    rd_req_size_urands[921]  = 20'd4;
    rd_req_size_urands[922]  = 20'd3;
    rd_req_size_urands[923]  = 20'd4;
    rd_req_size_urands[924]  = 20'd6;
    rd_req_size_urands[925]  = 20'd4;
    rd_req_size_urands[926]  = 20'd10;
    rd_req_size_urands[927]  = 20'd8;
    rd_req_size_urands[928]  = 20'd10;
    rd_req_size_urands[929]  = 20'd5;
    rd_req_size_urands[930]  = 20'd2;
    rd_req_size_urands[931]  = 20'd6;
    rd_req_size_urands[932]  = 20'd2;
    rd_req_size_urands[933]  = 20'd6;
    rd_req_size_urands[934]  = 20'd10;
    rd_req_size_urands[935]  = 20'd1;
    rd_req_size_urands[936]  = 20'd10;
    rd_req_size_urands[937]  = 20'd1;
    rd_req_size_urands[938]  = 20'd10;
    rd_req_size_urands[939]  = 20'd1;
    rd_req_size_urands[940]  = 20'd8;
    rd_req_size_urands[941]  = 20'd6;
    rd_req_size_urands[942]  = 20'd6;
    rd_req_size_urands[943]  = 20'd2;
    rd_req_size_urands[944]  = 20'd5;
    rd_req_size_urands[945]  = 20'd8;
    rd_req_size_urands[946]  = 20'd9;
    rd_req_size_urands[947]  = 20'd1;
    rd_req_size_urands[948]  = 20'd2;
    rd_req_size_urands[949]  = 20'd3;
    rd_req_size_urands[950]  = 20'd10;
    rd_req_size_urands[951]  = 20'd10;
    rd_req_size_urands[952]  = 20'd3;
    rd_req_size_urands[953]  = 20'd8;
    rd_req_size_urands[954]  = 20'd7;
    rd_req_size_urands[955]  = 20'd6;
    rd_req_size_urands[956]  = 20'd1;
    rd_req_size_urands[957]  = 20'd8;
    rd_req_size_urands[958]  = 20'd6;
    rd_req_size_urands[959]  = 20'd3;
    rd_req_size_urands[960]  = 20'd6;
    rd_req_size_urands[961]  = 20'd10;
    rd_req_size_urands[962]  = 20'd5;
    rd_req_size_urands[963]  = 20'd5;
    rd_req_size_urands[964]  = 20'd2;
    rd_req_size_urands[965]  = 20'd1;
    rd_req_size_urands[966]  = 20'd7;
    rd_req_size_urands[967]  = 20'd1;
    rd_req_size_urands[968]  = 20'd1;
    rd_req_size_urands[969]  = 20'd5;
    rd_req_size_urands[970]  = 20'd9;
    rd_req_size_urands[971]  = 20'd10;
    rd_req_size_urands[972]  = 20'd5;
    rd_req_size_urands[973]  = 20'd4;
    rd_req_size_urands[974]  = 20'd3;
    rd_req_size_urands[975]  = 20'd7;
    rd_req_size_urands[976]  = 20'd6;
    rd_req_size_urands[977]  = 20'd4;
    rd_req_size_urands[978]  = 20'd9;
    rd_req_size_urands[979]  = 20'd8;
    rd_req_size_urands[980]  = 20'd1;
    rd_req_size_urands[981]  = 20'd5;
    rd_req_size_urands[982]  = 20'd9;
    rd_req_size_urands[983]  = 20'd3;
    rd_req_size_urands[984]  = 20'd10;
    rd_req_size_urands[985]  = 20'd7;
    rd_req_size_urands[986]  = 20'd1;
    rd_req_size_urands[987]  = 20'd10;
    rd_req_size_urands[988]  = 20'd6;
    rd_req_size_urands[989]  = 20'd6;
    rd_req_size_urands[990]  = 20'd2;
    rd_req_size_urands[991]  = 20'd3;
    rd_req_size_urands[992]  = 20'd9;
    rd_req_size_urands[993]  = 20'd3;
    rd_req_size_urands[994]  = 20'd10;
    rd_req_size_urands[995]  = 20'd9;
    rd_req_size_urands[996]  = 20'd7;
    rd_req_size_urands[997]  = 20'd4;
    rd_req_size_urands[998]  = 20'd4;
    rd_req_size_urands[999]  = 20'd2;

    rd_req_pu_id_urands[0]    = 32'd3129082488;
    rd_req_pu_id_urands[1]    = 32'd4233799488;
    rd_req_pu_id_urands[2]    = 32'd2043998187;
    rd_req_pu_id_urands[3]    = 32'd340747405;
    rd_req_pu_id_urands[4]    = 32'd3138184934;
    rd_req_pu_id_urands[5]    = 32'd3677552271;
    rd_req_pu_id_urands[6]    = 32'd2596426268;
    rd_req_pu_id_urands[7]    = 32'd3344839173;
    rd_req_pu_id_urands[8]    = 32'd2896930078;
    rd_req_pu_id_urands[9]    = 32'd2531326996;
    rd_req_pu_id_urands[10]   = 32'd2416175395;
    rd_req_pu_id_urands[11]   = 32'd1764656823;
    rd_req_pu_id_urands[12]   = 32'd1628256755;
    rd_req_pu_id_urands[13]   = 32'd2370082769;
    rd_req_pu_id_urands[14]   = 32'd3487384310;
    rd_req_pu_id_urands[15]   = 32'd773819291;
    rd_req_pu_id_urands[16]   = 32'd4161258109;
    rd_req_pu_id_urands[17]   = 32'd2212227160;
    rd_req_pu_id_urands[18]   = 32'd3078389442;
    rd_req_pu_id_urands[19]   = 32'd2643374203;
    rd_req_pu_id_urands[20]   = 32'd267689879;
    rd_req_pu_id_urands[21]   = 32'd231294713;
    rd_req_pu_id_urands[22]   = 32'd4121449187;
    rd_req_pu_id_urands[23]   = 32'd2601380018;
    rd_req_pu_id_urands[24]   = 32'd3461225845;
    rd_req_pu_id_urands[25]   = 32'd4152488359;
    rd_req_pu_id_urands[26]   = 32'd1193978522;
    rd_req_pu_id_urands[27]   = 32'd1146857659;
    rd_req_pu_id_urands[28]   = 32'd214700482;
    rd_req_pu_id_urands[29]   = 32'd3540672149;
    rd_req_pu_id_urands[30]   = 32'd3529466481;
    rd_req_pu_id_urands[31]   = 32'd3611527662;
    rd_req_pu_id_urands[32]   = 32'd3245859674;
    rd_req_pu_id_urands[33]   = 32'd1962037124;
    rd_req_pu_id_urands[34]   = 32'd2200395875;
    rd_req_pu_id_urands[35]   = 32'd1202421432;
    rd_req_pu_id_urands[36]   = 32'd2355167398;
    rd_req_pu_id_urands[37]   = 32'd2780300903;
    rd_req_pu_id_urands[38]   = 32'd1288661937;
    rd_req_pu_id_urands[39]   = 32'd3644338595;
    rd_req_pu_id_urands[40]   = 32'd1967928033;
    rd_req_pu_id_urands[41]   = 32'd2539301044;
    rd_req_pu_id_urands[42]   = 32'd2433317692;
    rd_req_pu_id_urands[43]   = 32'd3867317737;
    rd_req_pu_id_urands[44]   = 32'd1597001887;
    rd_req_pu_id_urands[45]   = 32'd914514006;
    rd_req_pu_id_urands[46]   = 32'd958623613;
    rd_req_pu_id_urands[47]   = 32'd470861552;
    rd_req_pu_id_urands[48]   = 32'd3390771603;
    rd_req_pu_id_urands[49]   = 32'd195888953;
    rd_req_pu_id_urands[50]   = 32'd2741139984;
    rd_req_pu_id_urands[51]   = 32'd2866846900;
    rd_req_pu_id_urands[52]   = 32'd255556378;
    rd_req_pu_id_urands[53]   = 32'd4224879807;
    rd_req_pu_id_urands[54]   = 32'd3065190181;
    rd_req_pu_id_urands[55]   = 32'd3984863931;
    rd_req_pu_id_urands[56]   = 32'd3011296695;
    rd_req_pu_id_urands[57]   = 32'd80238342;
    rd_req_pu_id_urands[58]   = 32'd1110829982;
    rd_req_pu_id_urands[59]   = 32'd3208967053;
    rd_req_pu_id_urands[60]   = 32'd3659677768;
    rd_req_pu_id_urands[61]   = 32'd2774219046;
    rd_req_pu_id_urands[62]   = 32'd44677995;
    rd_req_pu_id_urands[63]   = 32'd1228992547;
    rd_req_pu_id_urands[64]   = 32'd1716164254;
    rd_req_pu_id_urands[65]   = 32'd923938646;
    rd_req_pu_id_urands[66]   = 32'd743339201;
    rd_req_pu_id_urands[67]   = 32'd543816952;
    rd_req_pu_id_urands[68]   = 32'd994005931;
    rd_req_pu_id_urands[69]   = 32'd42199010;
    rd_req_pu_id_urands[70]   = 32'd2612480549;
    rd_req_pu_id_urands[71]   = 32'd2791238727;
    rd_req_pu_id_urands[72]   = 32'd1757710190;
    rd_req_pu_id_urands[73]   = 32'd653383088;
    rd_req_pu_id_urands[74]   = 32'd3714747067;
    rd_req_pu_id_urands[75]   = 32'd1406267126;
    rd_req_pu_id_urands[76]   = 32'd3827192578;
    rd_req_pu_id_urands[77]   = 32'd147290781;
    rd_req_pu_id_urands[78]   = 32'd2973051452;
    rd_req_pu_id_urands[79]   = 32'd996880638;
    rd_req_pu_id_urands[80]   = 32'd2520727909;
    rd_req_pu_id_urands[81]   = 32'd414145251;
    rd_req_pu_id_urands[82]   = 32'd937531594;
    rd_req_pu_id_urands[83]   = 32'd2502894003;
    rd_req_pu_id_urands[84]   = 32'd253911758;
    rd_req_pu_id_urands[85]   = 32'd2007126422;
    rd_req_pu_id_urands[86]   = 32'd3781332960;
    rd_req_pu_id_urands[87]   = 32'd88161344;
    rd_req_pu_id_urands[88]   = 32'd3555859088;
    rd_req_pu_id_urands[89]   = 32'd577808438;
    rd_req_pu_id_urands[90]   = 32'd2021663723;
    rd_req_pu_id_urands[91]   = 32'd1741679526;
    rd_req_pu_id_urands[92]   = 32'd3087186698;
    rd_req_pu_id_urands[93]   = 32'd30782475;
    rd_req_pu_id_urands[94]   = 32'd1702646448;
    rd_req_pu_id_urands[95]   = 32'd1863461156;
    rd_req_pu_id_urands[96]   = 32'd4198977900;
    rd_req_pu_id_urands[97]   = 32'd1168146474;
    rd_req_pu_id_urands[98]   = 32'd709262493;
    rd_req_pu_id_urands[99]   = 32'd2404774797;
    rd_req_pu_id_urands[100]  = 32'd1730210920;
    rd_req_pu_id_urands[101]  = 32'd4232119082;
    rd_req_pu_id_urands[102]  = 32'd3184765224;
    rd_req_pu_id_urands[103]  = 32'd2896869378;
    rd_req_pu_id_urands[104]  = 32'd3345106261;
    rd_req_pu_id_urands[105]  = 32'd2031803818;
    rd_req_pu_id_urands[106]  = 32'd9660104;
    rd_req_pu_id_urands[107]  = 32'd3628782934;
    rd_req_pu_id_urands[108]  = 32'd4046908137;
    rd_req_pu_id_urands[109]  = 32'd4193632945;
    rd_req_pu_id_urands[110]  = 32'd1081977896;
    rd_req_pu_id_urands[111]  = 32'd1366945853;
    rd_req_pu_id_urands[112]  = 32'd3035099323;
    rd_req_pu_id_urands[113]  = 32'd2348335714;
    rd_req_pu_id_urands[114]  = 32'd1044586891;
    rd_req_pu_id_urands[115]  = 32'd2813319318;
    rd_req_pu_id_urands[116]  = 32'd1801630330;
    rd_req_pu_id_urands[117]  = 32'd995885885;
    rd_req_pu_id_urands[118]  = 32'd2942795647;
    rd_req_pu_id_urands[119]  = 32'd1128868904;
    rd_req_pu_id_urands[120]  = 32'd3894255835;
    rd_req_pu_id_urands[121]  = 32'd102909511;
    rd_req_pu_id_urands[122]  = 32'd165581048;
    rd_req_pu_id_urands[123]  = 32'd588506583;
    rd_req_pu_id_urands[124]  = 32'd2157229206;
    rd_req_pu_id_urands[125]  = 32'd3696543103;
    rd_req_pu_id_urands[126]  = 32'd3479013970;
    rd_req_pu_id_urands[127]  = 32'd598563993;
    rd_req_pu_id_urands[128]  = 32'd1041981233;
    rd_req_pu_id_urands[129]  = 32'd3814684218;
    rd_req_pu_id_urands[130]  = 32'd2035371815;
    rd_req_pu_id_urands[131]  = 32'd2202146824;
    rd_req_pu_id_urands[132]  = 32'd796433322;
    rd_req_pu_id_urands[133]  = 32'd1732425433;
    rd_req_pu_id_urands[134]  = 32'd1657022457;
    rd_req_pu_id_urands[135]  = 32'd2336618926;
    rd_req_pu_id_urands[136]  = 32'd1983806553;
    rd_req_pu_id_urands[137]  = 32'd3191016370;
    rd_req_pu_id_urands[138]  = 32'd3818977396;
    rd_req_pu_id_urands[139]  = 32'd2335728663;
    rd_req_pu_id_urands[140]  = 32'd298191374;
    rd_req_pu_id_urands[141]  = 32'd2263925224;
    rd_req_pu_id_urands[142]  = 32'd1353607815;
    rd_req_pu_id_urands[143]  = 32'd1017390368;
    rd_req_pu_id_urands[144]  = 32'd1870039146;
    rd_req_pu_id_urands[145]  = 32'd1583066433;
    rd_req_pu_id_urands[146]  = 32'd1486362290;
    rd_req_pu_id_urands[147]  = 32'd2787982551;
    rd_req_pu_id_urands[148]  = 32'd1151875490;
    rd_req_pu_id_urands[149]  = 32'd534189514;
    rd_req_pu_id_urands[150]  = 32'd2739414834;
    rd_req_pu_id_urands[151]  = 32'd689578312;
    rd_req_pu_id_urands[152]  = 32'd1086322651;
    rd_req_pu_id_urands[153]  = 32'd2405956328;
    rd_req_pu_id_urands[154]  = 32'd3192320991;
    rd_req_pu_id_urands[155]  = 32'd1138267096;
    rd_req_pu_id_urands[156]  = 32'd3492105367;
    rd_req_pu_id_urands[157]  = 32'd4081711681;
    rd_req_pu_id_urands[158]  = 32'd1897253950;
    rd_req_pu_id_urands[159]  = 32'd4098857775;
    rd_req_pu_id_urands[160]  = 32'd4060825460;
    rd_req_pu_id_urands[161]  = 32'd3792842712;
    rd_req_pu_id_urands[162]  = 32'd3140007711;
    rd_req_pu_id_urands[163]  = 32'd1756459501;
    rd_req_pu_id_urands[164]  = 32'd298939365;
    rd_req_pu_id_urands[165]  = 32'd3306440036;
    rd_req_pu_id_urands[166]  = 32'd1707382407;
    rd_req_pu_id_urands[167]  = 32'd3868027034;
    rd_req_pu_id_urands[168]  = 32'd2634409688;
    rd_req_pu_id_urands[169]  = 32'd3897877136;
    rd_req_pu_id_urands[170]  = 32'd3329039680;
    rd_req_pu_id_urands[171]  = 32'd834085996;
    rd_req_pu_id_urands[172]  = 32'd44176760;
    rd_req_pu_id_urands[173]  = 32'd3530896625;
    rd_req_pu_id_urands[174]  = 32'd4021753737;
    rd_req_pu_id_urands[175]  = 32'd34019385;
    rd_req_pu_id_urands[176]  = 32'd2370349865;
    rd_req_pu_id_urands[177]  = 32'd4219795560;
    rd_req_pu_id_urands[178]  = 32'd2302115445;
    rd_req_pu_id_urands[179]  = 32'd714585487;
    rd_req_pu_id_urands[180]  = 32'd3458257118;
    rd_req_pu_id_urands[181]  = 32'd1283182868;
    rd_req_pu_id_urands[182]  = 32'd3454006357;
    rd_req_pu_id_urands[183]  = 32'd2668754115;
    rd_req_pu_id_urands[184]  = 32'd1515313500;
    rd_req_pu_id_urands[185]  = 32'd3276169175;
    rd_req_pu_id_urands[186]  = 32'd4240557633;
    rd_req_pu_id_urands[187]  = 32'd1534023769;
    rd_req_pu_id_urands[188]  = 32'd1427783373;
    rd_req_pu_id_urands[189]  = 32'd933101718;
    rd_req_pu_id_urands[190]  = 32'd3521611325;
    rd_req_pu_id_urands[191]  = 32'd1383209736;
    rd_req_pu_id_urands[192]  = 32'd55953825;
    rd_req_pu_id_urands[193]  = 32'd633440243;
    rd_req_pu_id_urands[194]  = 32'd614026541;
    rd_req_pu_id_urands[195]  = 32'd2047340940;
    rd_req_pu_id_urands[196]  = 32'd3952779987;
    rd_req_pu_id_urands[197]  = 32'd1998622871;
    rd_req_pu_id_urands[198]  = 32'd2392770975;
    rd_req_pu_id_urands[199]  = 32'd1634883654;
    rd_req_pu_id_urands[200]  = 32'd4009730858;
    rd_req_pu_id_urands[201]  = 32'd3043570310;
    rd_req_pu_id_urands[202]  = 32'd3492311087;
    rd_req_pu_id_urands[203]  = 32'd2806238830;
    rd_req_pu_id_urands[204]  = 32'd2537978835;
    rd_req_pu_id_urands[205]  = 32'd2925709332;
    rd_req_pu_id_urands[206]  = 32'd3877844537;
    rd_req_pu_id_urands[207]  = 32'd1371755030;
    rd_req_pu_id_urands[208]  = 32'd850242523;
    rd_req_pu_id_urands[209]  = 32'd2908289741;
    rd_req_pu_id_urands[210]  = 32'd169939246;
    rd_req_pu_id_urands[211]  = 32'd571051759;
    rd_req_pu_id_urands[212]  = 32'd2726026262;
    rd_req_pu_id_urands[213]  = 32'd3996677555;
    rd_req_pu_id_urands[214]  = 32'd2281751212;
    rd_req_pu_id_urands[215]  = 32'd1149843904;
    rd_req_pu_id_urands[216]  = 32'd3047245829;
    rd_req_pu_id_urands[217]  = 32'd656771051;
    rd_req_pu_id_urands[218]  = 32'd839173959;
    rd_req_pu_id_urands[219]  = 32'd2939523921;
    rd_req_pu_id_urands[220]  = 32'd3541736717;
    rd_req_pu_id_urands[221]  = 32'd1269930512;
    rd_req_pu_id_urands[222]  = 32'd1904605186;
    rd_req_pu_id_urands[223]  = 32'd228181188;
    rd_req_pu_id_urands[224]  = 32'd552458724;
    rd_req_pu_id_urands[225]  = 32'd3946852222;
    rd_req_pu_id_urands[226]  = 32'd1587236053;
    rd_req_pu_id_urands[227]  = 32'd766039586;
    rd_req_pu_id_urands[228]  = 32'd16690743;
    rd_req_pu_id_urands[229]  = 32'd1027365865;
    rd_req_pu_id_urands[230]  = 32'd1065384873;
    rd_req_pu_id_urands[231]  = 32'd886996338;
    rd_req_pu_id_urands[232]  = 32'd2398784975;
    rd_req_pu_id_urands[233]  = 32'd698208329;
    rd_req_pu_id_urands[234]  = 32'd3373907162;
    rd_req_pu_id_urands[235]  = 32'd929399088;
    rd_req_pu_id_urands[236]  = 32'd3525071527;
    rd_req_pu_id_urands[237]  = 32'd1727564328;
    rd_req_pu_id_urands[238]  = 32'd940772333;
    rd_req_pu_id_urands[239]  = 32'd533227910;
    rd_req_pu_id_urands[240]  = 32'd4154510356;
    rd_req_pu_id_urands[241]  = 32'd1088188064;
    rd_req_pu_id_urands[242]  = 32'd3970380382;
    rd_req_pu_id_urands[243]  = 32'd985392314;
    rd_req_pu_id_urands[244]  = 32'd1588359449;
    rd_req_pu_id_urands[245]  = 32'd2912296681;
    rd_req_pu_id_urands[246]  = 32'd940569784;
    rd_req_pu_id_urands[247]  = 32'd3092458705;
    rd_req_pu_id_urands[248]  = 32'd2063954417;
    rd_req_pu_id_urands[249]  = 32'd1395283634;
    rd_req_pu_id_urands[250]  = 32'd3230120785;
    rd_req_pu_id_urands[251]  = 32'd1052830128;
    rd_req_pu_id_urands[252]  = 32'd2478178307;
    rd_req_pu_id_urands[253]  = 32'd1261757571;
    rd_req_pu_id_urands[254]  = 32'd698897836;
    rd_req_pu_id_urands[255]  = 32'd898356231;
    rd_req_pu_id_urands[256]  = 32'd513833655;
    rd_req_pu_id_urands[257]  = 32'd1209661414;
    rd_req_pu_id_urands[258]  = 32'd2535607960;
    rd_req_pu_id_urands[259]  = 32'd933079923;
    rd_req_pu_id_urands[260]  = 32'd1329881970;
    rd_req_pu_id_urands[261]  = 32'd558111259;
    rd_req_pu_id_urands[262]  = 32'd3399691756;
    rd_req_pu_id_urands[263]  = 32'd2948276877;
    rd_req_pu_id_urands[264]  = 32'd1249474429;
    rd_req_pu_id_urands[265]  = 32'd1243485222;
    rd_req_pu_id_urands[266]  = 32'd992310209;
    rd_req_pu_id_urands[267]  = 32'd583001025;
    rd_req_pu_id_urands[268]  = 32'd3104671131;
    rd_req_pu_id_urands[269]  = 32'd3232654766;
    rd_req_pu_id_urands[270]  = 32'd951565499;
    rd_req_pu_id_urands[271]  = 32'd3290926394;
    rd_req_pu_id_urands[272]  = 32'd1577452284;
    rd_req_pu_id_urands[273]  = 32'd3749101140;
    rd_req_pu_id_urands[274]  = 32'd66351140;
    rd_req_pu_id_urands[275]  = 32'd1549297767;
    rd_req_pu_id_urands[276]  = 32'd296549009;
    rd_req_pu_id_urands[277]  = 32'd918938091;
    rd_req_pu_id_urands[278]  = 32'd3183059875;
    rd_req_pu_id_urands[279]  = 32'd1795911313;
    rd_req_pu_id_urands[280]  = 32'd1881322694;
    rd_req_pu_id_urands[281]  = 32'd3552152674;
    rd_req_pu_id_urands[282]  = 32'd82277783;
    rd_req_pu_id_urands[283]  = 32'd774481798;
    rd_req_pu_id_urands[284]  = 32'd1503999739;
    rd_req_pu_id_urands[285]  = 32'd3499429173;
    rd_req_pu_id_urands[286]  = 32'd1121864852;
    rd_req_pu_id_urands[287]  = 32'd941256573;
    rd_req_pu_id_urands[288]  = 32'd2920953104;
    rd_req_pu_id_urands[289]  = 32'd1321081708;
    rd_req_pu_id_urands[290]  = 32'd164597839;
    rd_req_pu_id_urands[291]  = 32'd2613709421;
    rd_req_pu_id_urands[292]  = 32'd1840794015;
    rd_req_pu_id_urands[293]  = 32'd2534849669;
    rd_req_pu_id_urands[294]  = 32'd1013388586;
    rd_req_pu_id_urands[295]  = 32'd1319523952;
    rd_req_pu_id_urands[296]  = 32'd1352687645;
    rd_req_pu_id_urands[297]  = 32'd2424907711;
    rd_req_pu_id_urands[298]  = 32'd3391776688;
    rd_req_pu_id_urands[299]  = 32'd4038199222;
    rd_req_pu_id_urands[300]  = 32'd1143732278;
    rd_req_pu_id_urands[301]  = 32'd595315442;
    rd_req_pu_id_urands[302]  = 32'd1570937254;
    rd_req_pu_id_urands[303]  = 32'd341225020;
    rd_req_pu_id_urands[304]  = 32'd4077812177;
    rd_req_pu_id_urands[305]  = 32'd2220717878;
    rd_req_pu_id_urands[306]  = 32'd3108451738;
    rd_req_pu_id_urands[307]  = 32'd3135399907;
    rd_req_pu_id_urands[308]  = 32'd3798229889;
    rd_req_pu_id_urands[309]  = 32'd643896285;
    rd_req_pu_id_urands[310]  = 32'd1409138357;
    rd_req_pu_id_urands[311]  = 32'd1433335830;
    rd_req_pu_id_urands[312]  = 32'd4208514742;
    rd_req_pu_id_urands[313]  = 32'd3087105172;
    rd_req_pu_id_urands[314]  = 32'd1688935774;
    rd_req_pu_id_urands[315]  = 32'd1153224008;
    rd_req_pu_id_urands[316]  = 32'd2220014707;
    rd_req_pu_id_urands[317]  = 32'd1843958659;
    rd_req_pu_id_urands[318]  = 32'd535335540;
    rd_req_pu_id_urands[319]  = 32'd1812293330;
    rd_req_pu_id_urands[320]  = 32'd3043680989;
    rd_req_pu_id_urands[321]  = 32'd252283065;
    rd_req_pu_id_urands[322]  = 32'd2022435330;
    rd_req_pu_id_urands[323]  = 32'd2523550602;
    rd_req_pu_id_urands[324]  = 32'd3536009961;
    rd_req_pu_id_urands[325]  = 32'd784120609;
    rd_req_pu_id_urands[326]  = 32'd3919847511;
    rd_req_pu_id_urands[327]  = 32'd4255400336;
    rd_req_pu_id_urands[328]  = 32'd791614843;
    rd_req_pu_id_urands[329]  = 32'd1374177897;
    rd_req_pu_id_urands[330]  = 32'd2077106225;
    rd_req_pu_id_urands[331]  = 32'd4201306234;
    rd_req_pu_id_urands[332]  = 32'd1552536763;
    rd_req_pu_id_urands[333]  = 32'd3563553687;
    rd_req_pu_id_urands[334]  = 32'd2159021876;
    rd_req_pu_id_urands[335]  = 32'd1468173138;
    rd_req_pu_id_urands[336]  = 32'd3118775615;
    rd_req_pu_id_urands[337]  = 32'd2104063814;
    rd_req_pu_id_urands[338]  = 32'd3700332420;
    rd_req_pu_id_urands[339]  = 32'd3907677645;
    rd_req_pu_id_urands[340]  = 32'd2198674866;
    rd_req_pu_id_urands[341]  = 32'd2942566592;
    rd_req_pu_id_urands[342]  = 32'd4165188328;
    rd_req_pu_id_urands[343]  = 32'd4292265205;
    rd_req_pu_id_urands[344]  = 32'd1175867971;
    rd_req_pu_id_urands[345]  = 32'd2930741731;
    rd_req_pu_id_urands[346]  = 32'd493415739;
    rd_req_pu_id_urands[347]  = 32'd1444908647;
    rd_req_pu_id_urands[348]  = 32'd4172629010;
    rd_req_pu_id_urands[349]  = 32'd65007862;
    rd_req_pu_id_urands[350]  = 32'd3120900465;
    rd_req_pu_id_urands[351]  = 32'd3281897652;
    rd_req_pu_id_urands[352]  = 32'd3209955650;
    rd_req_pu_id_urands[353]  = 32'd756069956;
    rd_req_pu_id_urands[354]  = 32'd886232353;
    rd_req_pu_id_urands[355]  = 32'd3451315228;
    rd_req_pu_id_urands[356]  = 32'd158033983;
    rd_req_pu_id_urands[357]  = 32'd524447908;
    rd_req_pu_id_urands[358]  = 32'd1390604515;
    rd_req_pu_id_urands[359]  = 32'd918396983;
    rd_req_pu_id_urands[360]  = 32'd1879176497;
    rd_req_pu_id_urands[361]  = 32'd1746545241;
    rd_req_pu_id_urands[362]  = 32'd1146149367;
    rd_req_pu_id_urands[363]  = 32'd796434971;
    rd_req_pu_id_urands[364]  = 32'd2464536998;
    rd_req_pu_id_urands[365]  = 32'd5770007;
    rd_req_pu_id_urands[366]  = 32'd2397939347;
    rd_req_pu_id_urands[367]  = 32'd2534328263;
    rd_req_pu_id_urands[368]  = 32'd2894776579;
    rd_req_pu_id_urands[369]  = 32'd1683188123;
    rd_req_pu_id_urands[370]  = 32'd108156412;
    rd_req_pu_id_urands[371]  = 32'd1164611320;
    rd_req_pu_id_urands[372]  = 32'd560557624;
    rd_req_pu_id_urands[373]  = 32'd4117707409;
    rd_req_pu_id_urands[374]  = 32'd291394407;
    rd_req_pu_id_urands[375]  = 32'd3885086170;
    rd_req_pu_id_urands[376]  = 32'd3182785899;
    rd_req_pu_id_urands[377]  = 32'd8598654;
    rd_req_pu_id_urands[378]  = 32'd1374497702;
    rd_req_pu_id_urands[379]  = 32'd873842800;
    rd_req_pu_id_urands[380]  = 32'd1214169388;
    rd_req_pu_id_urands[381]  = 32'd115761588;
    rd_req_pu_id_urands[382]  = 32'd3106040063;
    rd_req_pu_id_urands[383]  = 32'd465373867;
    rd_req_pu_id_urands[384]  = 32'd647263600;
    rd_req_pu_id_urands[385]  = 32'd2186405880;
    rd_req_pu_id_urands[386]  = 32'd3940117315;
    rd_req_pu_id_urands[387]  = 32'd1356468602;
    rd_req_pu_id_urands[388]  = 32'd2416398034;
    rd_req_pu_id_urands[389]  = 32'd4066182207;
    rd_req_pu_id_urands[390]  = 32'd3703291004;
    rd_req_pu_id_urands[391]  = 32'd3791559584;
    rd_req_pu_id_urands[392]  = 32'd739404138;
    rd_req_pu_id_urands[393]  = 32'd1654647129;
    rd_req_pu_id_urands[394]  = 32'd512004208;
    rd_req_pu_id_urands[395]  = 32'd3756702748;
    rd_req_pu_id_urands[396]  = 32'd2867336256;
    rd_req_pu_id_urands[397]  = 32'd922325528;
    rd_req_pu_id_urands[398]  = 32'd338266524;
    rd_req_pu_id_urands[399]  = 32'd3924558095;
    rd_req_pu_id_urands[400]  = 32'd1605220338;
    rd_req_pu_id_urands[401]  = 32'd2749708976;
    rd_req_pu_id_urands[402]  = 32'd193699155;
    rd_req_pu_id_urands[403]  = 32'd1017402843;
    rd_req_pu_id_urands[404]  = 32'd2464138022;
    rd_req_pu_id_urands[405]  = 32'd1187817980;
    rd_req_pu_id_urands[406]  = 32'd3900555209;
    rd_req_pu_id_urands[407]  = 32'd3986895400;
    rd_req_pu_id_urands[408]  = 32'd1197887581;
    rd_req_pu_id_urands[409]  = 32'd3059051152;
    rd_req_pu_id_urands[410]  = 32'd3356692047;
    rd_req_pu_id_urands[411]  = 32'd489212940;
    rd_req_pu_id_urands[412]  = 32'd3106919335;
    rd_req_pu_id_urands[413]  = 32'd2229227104;
    rd_req_pu_id_urands[414]  = 32'd4198888467;
    rd_req_pu_id_urands[415]  = 32'd2997764163;
    rd_req_pu_id_urands[416]  = 32'd88814489;
    rd_req_pu_id_urands[417]  = 32'd3225195500;
    rd_req_pu_id_urands[418]  = 32'd615889130;
    rd_req_pu_id_urands[419]  = 32'd3837727152;
    rd_req_pu_id_urands[420]  = 32'd2751043539;
    rd_req_pu_id_urands[421]  = 32'd3703894029;
    rd_req_pu_id_urands[422]  = 32'd3288067273;
    rd_req_pu_id_urands[423]  = 32'd2802297139;
    rd_req_pu_id_urands[424]  = 32'd2177782301;
    rd_req_pu_id_urands[425]  = 32'd423756398;
    rd_req_pu_id_urands[426]  = 32'd2112118708;
    rd_req_pu_id_urands[427]  = 32'd2925369982;
    rd_req_pu_id_urands[428]  = 32'd1756732247;
    rd_req_pu_id_urands[429]  = 32'd3847782033;
    rd_req_pu_id_urands[430]  = 32'd2844083649;
    rd_req_pu_id_urands[431]  = 32'd1652816483;
    rd_req_pu_id_urands[432]  = 32'd2044438135;
    rd_req_pu_id_urands[433]  = 32'd3176510723;
    rd_req_pu_id_urands[434]  = 32'd1187887536;
    rd_req_pu_id_urands[435]  = 32'd3384731957;
    rd_req_pu_id_urands[436]  = 32'd2925221961;
    rd_req_pu_id_urands[437]  = 32'd1814743098;
    rd_req_pu_id_urands[438]  = 32'd773462620;
    rd_req_pu_id_urands[439]  = 32'd717280951;
    rd_req_pu_id_urands[440]  = 32'd1013927605;
    rd_req_pu_id_urands[441]  = 32'd3232147572;
    rd_req_pu_id_urands[442]  = 32'd1523093770;
    rd_req_pu_id_urands[443]  = 32'd522677819;
    rd_req_pu_id_urands[444]  = 32'd183550134;
    rd_req_pu_id_urands[445]  = 32'd3891897853;
    rd_req_pu_id_urands[446]  = 32'd429379083;
    rd_req_pu_id_urands[447]  = 32'd588930500;
    rd_req_pu_id_urands[448]  = 32'd1140038497;
    rd_req_pu_id_urands[449]  = 32'd1627177038;
    rd_req_pu_id_urands[450]  = 32'd3372835123;
    rd_req_pu_id_urands[451]  = 32'd2030419187;
    rd_req_pu_id_urands[452]  = 32'd4111795113;
    rd_req_pu_id_urands[453]  = 32'd22631747;
    rd_req_pu_id_urands[454]  = 32'd2273758056;
    rd_req_pu_id_urands[455]  = 32'd2375601129;
    rd_req_pu_id_urands[456]  = 32'd667561351;
    rd_req_pu_id_urands[457]  = 32'd688744841;
    rd_req_pu_id_urands[458]  = 32'd3296313487;
    rd_req_pu_id_urands[459]  = 32'd2742835136;
    rd_req_pu_id_urands[460]  = 32'd1152389434;
    rd_req_pu_id_urands[461]  = 32'd4028968290;
    rd_req_pu_id_urands[462]  = 32'd3757772942;
    rd_req_pu_id_urands[463]  = 32'd578592552;
    rd_req_pu_id_urands[464]  = 32'd263440149;
    rd_req_pu_id_urands[465]  = 32'd2146736821;
    rd_req_pu_id_urands[466]  = 32'd760869342;
    rd_req_pu_id_urands[467]  = 32'd1046779794;
    rd_req_pu_id_urands[468]  = 32'd4054671625;
    rd_req_pu_id_urands[469]  = 32'd713936011;
    rd_req_pu_id_urands[470]  = 32'd2483542765;
    rd_req_pu_id_urands[471]  = 32'd2874827643;
    rd_req_pu_id_urands[472]  = 32'd880192085;
    rd_req_pu_id_urands[473]  = 32'd4103467921;
    rd_req_pu_id_urands[474]  = 32'd3240829929;
    rd_req_pu_id_urands[475]  = 32'd792594848;
    rd_req_pu_id_urands[476]  = 32'd2788249497;
    rd_req_pu_id_urands[477]  = 32'd497727877;
    rd_req_pu_id_urands[478]  = 32'd1104075002;
    rd_req_pu_id_urands[479]  = 32'd3372039593;
    rd_req_pu_id_urands[480]  = 32'd1958069706;
    rd_req_pu_id_urands[481]  = 32'd203346201;
    rd_req_pu_id_urands[482]  = 32'd92957797;
    rd_req_pu_id_urands[483]  = 32'd2484745912;
    rd_req_pu_id_urands[484]  = 32'd911621962;
    rd_req_pu_id_urands[485]  = 32'd2325764768;
    rd_req_pu_id_urands[486]  = 32'd15224614;
    rd_req_pu_id_urands[487]  = 32'd3901805380;
    rd_req_pu_id_urands[488]  = 32'd936287007;
    rd_req_pu_id_urands[489]  = 32'd1572980434;
    rd_req_pu_id_urands[490]  = 32'd2564900914;
    rd_req_pu_id_urands[491]  = 32'd1517605760;
    rd_req_pu_id_urands[492]  = 32'd2138085827;
    rd_req_pu_id_urands[493]  = 32'd1504103161;
    rd_req_pu_id_urands[494]  = 32'd2378286107;
    rd_req_pu_id_urands[495]  = 32'd3620367537;
    rd_req_pu_id_urands[496]  = 32'd744899610;
    rd_req_pu_id_urands[497]  = 32'd6351710;
    rd_req_pu_id_urands[498]  = 32'd1694658213;
    rd_req_pu_id_urands[499]  = 32'd869858665;
    rd_req_pu_id_urands[500]  = 32'd3391788345;
    rd_req_pu_id_urands[501]  = 32'd3067679196;
    rd_req_pu_id_urands[502]  = 32'd3691447213;
    rd_req_pu_id_urands[503]  = 32'd686628538;
    rd_req_pu_id_urands[504]  = 32'd249063717;
    rd_req_pu_id_urands[505]  = 32'd985739974;
    rd_req_pu_id_urands[506]  = 32'd465929258;
    rd_req_pu_id_urands[507]  = 32'd1708057641;
    rd_req_pu_id_urands[508]  = 32'd1162111725;
    rd_req_pu_id_urands[509]  = 32'd2580789535;
    rd_req_pu_id_urands[510]  = 32'd3140680024;
    rd_req_pu_id_urands[511]  = 32'd1268556462;
    rd_req_pu_id_urands[512]  = 32'd1678607997;
    rd_req_pu_id_urands[513]  = 32'd746372356;
    rd_req_pu_id_urands[514]  = 32'd3811958534;
    rd_req_pu_id_urands[515]  = 32'd1506867149;
    rd_req_pu_id_urands[516]  = 32'd1954514936;
    rd_req_pu_id_urands[517]  = 32'd1809816733;
    rd_req_pu_id_urands[518]  = 32'd6478824;
    rd_req_pu_id_urands[519]  = 32'd1375461457;
    rd_req_pu_id_urands[520]  = 32'd1731465737;
    rd_req_pu_id_urands[521]  = 32'd3124584909;
    rd_req_pu_id_urands[522]  = 32'd4028281608;
    rd_req_pu_id_urands[523]  = 32'd1226860887;
    rd_req_pu_id_urands[524]  = 32'd1406039487;
    rd_req_pu_id_urands[525]  = 32'd1023540840;
    rd_req_pu_id_urands[526]  = 32'd3898477317;
    rd_req_pu_id_urands[527]  = 32'd3786111702;
    rd_req_pu_id_urands[528]  = 32'd1699314973;
    rd_req_pu_id_urands[529]  = 32'd280522418;
    rd_req_pu_id_urands[530]  = 32'd3130699197;
    rd_req_pu_id_urands[531]  = 32'd4202259903;
    rd_req_pu_id_urands[532]  = 32'd4189090820;
    rd_req_pu_id_urands[533]  = 32'd3813409792;
    rd_req_pu_id_urands[534]  = 32'd2273750177;
    rd_req_pu_id_urands[535]  = 32'd2396289779;
    rd_req_pu_id_urands[536]  = 32'd798721050;
    rd_req_pu_id_urands[537]  = 32'd1826196927;
    rd_req_pu_id_urands[538]  = 32'd3422826178;
    rd_req_pu_id_urands[539]  = 32'd3352613131;
    rd_req_pu_id_urands[540]  = 32'd3989519998;
    rd_req_pu_id_urands[541]  = 32'd1558843222;
    rd_req_pu_id_urands[542]  = 32'd712619808;
    rd_req_pu_id_urands[543]  = 32'd301418011;
    rd_req_pu_id_urands[544]  = 32'd2341128368;
    rd_req_pu_id_urands[545]  = 32'd1255356721;
    rd_req_pu_id_urands[546]  = 32'd3242756466;
    rd_req_pu_id_urands[547]  = 32'd2061447063;
    rd_req_pu_id_urands[548]  = 32'd632525302;
    rd_req_pu_id_urands[549]  = 32'd1738722409;
    rd_req_pu_id_urands[550]  = 32'd857503194;
    rd_req_pu_id_urands[551]  = 32'd3210757802;
    rd_req_pu_id_urands[552]  = 32'd992118435;
    rd_req_pu_id_urands[553]  = 32'd3963993537;
    rd_req_pu_id_urands[554]  = 32'd948213309;
    rd_req_pu_id_urands[555]  = 32'd3291424342;
    rd_req_pu_id_urands[556]  = 32'd1589483988;
    rd_req_pu_id_urands[557]  = 32'd2644436840;
    rd_req_pu_id_urands[558]  = 32'd996032156;
    rd_req_pu_id_urands[559]  = 32'd3446698542;
    rd_req_pu_id_urands[560]  = 32'd483128254;
    rd_req_pu_id_urands[561]  = 32'd3866002375;
    rd_req_pu_id_urands[562]  = 32'd2284539437;
    rd_req_pu_id_urands[563]  = 32'd2887634031;
    rd_req_pu_id_urands[564]  = 32'd1432342905;
    rd_req_pu_id_urands[565]  = 32'd3384414118;
    rd_req_pu_id_urands[566]  = 32'd2460175132;
    rd_req_pu_id_urands[567]  = 32'd2546486485;
    rd_req_pu_id_urands[568]  = 32'd1904028747;
    rd_req_pu_id_urands[569]  = 32'd1715735207;
    rd_req_pu_id_urands[570]  = 32'd3832001187;
    rd_req_pu_id_urands[571]  = 32'd3152155437;
    rd_req_pu_id_urands[572]  = 32'd415476517;
    rd_req_pu_id_urands[573]  = 32'd4106047463;
    rd_req_pu_id_urands[574]  = 32'd3776811680;
    rd_req_pu_id_urands[575]  = 32'd1531944805;
    rd_req_pu_id_urands[576]  = 32'd3794655580;
    rd_req_pu_id_urands[577]  = 32'd2299060660;
    rd_req_pu_id_urands[578]  = 32'd2752482506;
    rd_req_pu_id_urands[579]  = 32'd4041079569;
    rd_req_pu_id_urands[580]  = 32'd2402754733;
    rd_req_pu_id_urands[581]  = 32'd1967300181;
    rd_req_pu_id_urands[582]  = 32'd209097640;
    rd_req_pu_id_urands[583]  = 32'd2378660104;
    rd_req_pu_id_urands[584]  = 32'd448270403;
    rd_req_pu_id_urands[585]  = 32'd2266025069;
    rd_req_pu_id_urands[586]  = 32'd318177675;
    rd_req_pu_id_urands[587]  = 32'd886320929;
    rd_req_pu_id_urands[588]  = 32'd27370506;
    rd_req_pu_id_urands[589]  = 32'd3407908281;
    rd_req_pu_id_urands[590]  = 32'd1065198947;
    rd_req_pu_id_urands[591]  = 32'd3266280116;
    rd_req_pu_id_urands[592]  = 32'd2431904228;
    rd_req_pu_id_urands[593]  = 32'd3755382352;
    rd_req_pu_id_urands[594]  = 32'd944058903;
    rd_req_pu_id_urands[595]  = 32'd4224829752;
    rd_req_pu_id_urands[596]  = 32'd3190048589;
    rd_req_pu_id_urands[597]  = 32'd2775444367;
    rd_req_pu_id_urands[598]  = 32'd340285656;
    rd_req_pu_id_urands[599]  = 32'd1979411180;
    rd_req_pu_id_urands[600]  = 32'd1254609815;
    rd_req_pu_id_urands[601]  = 32'd2632894412;
    rd_req_pu_id_urands[602]  = 32'd488059823;
    rd_req_pu_id_urands[603]  = 32'd1538155523;
    rd_req_pu_id_urands[604]  = 32'd2239481222;
    rd_req_pu_id_urands[605]  = 32'd1535496396;
    rd_req_pu_id_urands[606]  = 32'd3994846080;
    rd_req_pu_id_urands[607]  = 32'd448802341;
    rd_req_pu_id_urands[608]  = 32'd4226104200;
    rd_req_pu_id_urands[609]  = 32'd2966182262;
    rd_req_pu_id_urands[610]  = 32'd3244770000;
    rd_req_pu_id_urands[611]  = 32'd1969065558;
    rd_req_pu_id_urands[612]  = 32'd2851986028;
    rd_req_pu_id_urands[613]  = 32'd2289469255;
    rd_req_pu_id_urands[614]  = 32'd3482218367;
    rd_req_pu_id_urands[615]  = 32'd4135985419;
    rd_req_pu_id_urands[616]  = 32'd3751657568;
    rd_req_pu_id_urands[617]  = 32'd770020575;
    rd_req_pu_id_urands[618]  = 32'd3159128289;
    rd_req_pu_id_urands[619]  = 32'd2859139680;
    rd_req_pu_id_urands[620]  = 32'd2025653776;
    rd_req_pu_id_urands[621]  = 32'd2674085499;
    rd_req_pu_id_urands[622]  = 32'd4001305528;
    rd_req_pu_id_urands[623]  = 32'd3723860345;
    rd_req_pu_id_urands[624]  = 32'd1369223892;
    rd_req_pu_id_urands[625]  = 32'd2736067190;
    rd_req_pu_id_urands[626]  = 32'd1185127811;
    rd_req_pu_id_urands[627]  = 32'd2826958210;
    rd_req_pu_id_urands[628]  = 32'd3996701439;
    rd_req_pu_id_urands[629]  = 32'd2540581715;
    rd_req_pu_id_urands[630]  = 32'd4007315512;
    rd_req_pu_id_urands[631]  = 32'd1139888273;
    rd_req_pu_id_urands[632]  = 32'd1940892978;
    rd_req_pu_id_urands[633]  = 32'd4067733660;
    rd_req_pu_id_urands[634]  = 32'd1133088295;
    rd_req_pu_id_urands[635]  = 32'd1506979789;
    rd_req_pu_id_urands[636]  = 32'd3836961068;
    rd_req_pu_id_urands[637]  = 32'd3864962799;
    rd_req_pu_id_urands[638]  = 32'd2473367392;
    rd_req_pu_id_urands[639]  = 32'd843423656;
    rd_req_pu_id_urands[640]  = 32'd1740741664;
    rd_req_pu_id_urands[641]  = 32'd1183995543;
    rd_req_pu_id_urands[642]  = 32'd217313778;
    rd_req_pu_id_urands[643]  = 32'd2227425702;
    rd_req_pu_id_urands[644]  = 32'd2816058767;
    rd_req_pu_id_urands[645]  = 32'd2895092049;
    rd_req_pu_id_urands[646]  = 32'd2947829331;
    rd_req_pu_id_urands[647]  = 32'd2466963008;
    rd_req_pu_id_urands[648]  = 32'd3162824708;
    rd_req_pu_id_urands[649]  = 32'd3246308633;
    rd_req_pu_id_urands[650]  = 32'd859522832;
    rd_req_pu_id_urands[651]  = 32'd4176369580;
    rd_req_pu_id_urands[652]  = 32'd426116078;
    rd_req_pu_id_urands[653]  = 32'd3837792164;
    rd_req_pu_id_urands[654]  = 32'd100023910;
    rd_req_pu_id_urands[655]  = 32'd4236689852;
    rd_req_pu_id_urands[656]  = 32'd1053168519;
    rd_req_pu_id_urands[657]  = 32'd3227163000;
    rd_req_pu_id_urands[658]  = 32'd3620089453;
    rd_req_pu_id_urands[659]  = 32'd2733025786;
    rd_req_pu_id_urands[660]  = 32'd2240507291;
    rd_req_pu_id_urands[661]  = 32'd2651857428;
    rd_req_pu_id_urands[662]  = 32'd3644837452;
    rd_req_pu_id_urands[663]  = 32'd163816370;
    rd_req_pu_id_urands[664]  = 32'd1746377627;
    rd_req_pu_id_urands[665]  = 32'd3791364364;
    rd_req_pu_id_urands[666]  = 32'd3275209460;
    rd_req_pu_id_urands[667]  = 32'd1002205746;
    rd_req_pu_id_urands[668]  = 32'd565742893;
    rd_req_pu_id_urands[669]  = 32'd2854780061;
    rd_req_pu_id_urands[670]  = 32'd2847444981;
    rd_req_pu_id_urands[671]  = 32'd4225497705;
    rd_req_pu_id_urands[672]  = 32'd2681258330;
    rd_req_pu_id_urands[673]  = 32'd640203782;
    rd_req_pu_id_urands[674]  = 32'd2922577775;
    rd_req_pu_id_urands[675]  = 32'd626323802;
    rd_req_pu_id_urands[676]  = 32'd3478879662;
    rd_req_pu_id_urands[677]  = 32'd1183762138;
    rd_req_pu_id_urands[678]  = 32'd2213475250;
    rd_req_pu_id_urands[679]  = 32'd1932407316;
    rd_req_pu_id_urands[680]  = 32'd1793416208;
    rd_req_pu_id_urands[681]  = 32'd1104888588;
    rd_req_pu_id_urands[682]  = 32'd1181273466;
    rd_req_pu_id_urands[683]  = 32'd3770367113;
    rd_req_pu_id_urands[684]  = 32'd1534915203;
    rd_req_pu_id_urands[685]  = 32'd1897899484;
    rd_req_pu_id_urands[686]  = 32'd3264205684;
    rd_req_pu_id_urands[687]  = 32'd2011316702;
    rd_req_pu_id_urands[688]  = 32'd2820499698;
    rd_req_pu_id_urands[689]  = 32'd515804124;
    rd_req_pu_id_urands[690]  = 32'd2145329834;
    rd_req_pu_id_urands[691]  = 32'd2338797950;
    rd_req_pu_id_urands[692]  = 32'd845498944;
    rd_req_pu_id_urands[693]  = 32'd295717013;
    rd_req_pu_id_urands[694]  = 32'd840910509;
    rd_req_pu_id_urands[695]  = 32'd490594730;
    rd_req_pu_id_urands[696]  = 32'd2160181373;
    rd_req_pu_id_urands[697]  = 32'd2981780776;
    rd_req_pu_id_urands[698]  = 32'd3535941814;
    rd_req_pu_id_urands[699]  = 32'd2992785380;
    rd_req_pu_id_urands[700]  = 32'd3057855597;
    rd_req_pu_id_urands[701]  = 32'd38710253;
    rd_req_pu_id_urands[702]  = 32'd2234286975;
    rd_req_pu_id_urands[703]  = 32'd3204180961;
    rd_req_pu_id_urands[704]  = 32'd4070239506;
    rd_req_pu_id_urands[705]  = 32'd3480327799;
    rd_req_pu_id_urands[706]  = 32'd1504804575;
    rd_req_pu_id_urands[707]  = 32'd3549280109;
    rd_req_pu_id_urands[708]  = 32'd2219273118;
    rd_req_pu_id_urands[709]  = 32'd4206185136;
    rd_req_pu_id_urands[710]  = 32'd2384688915;
    rd_req_pu_id_urands[711]  = 32'd2023164490;
    rd_req_pu_id_urands[712]  = 32'd148576660;
    rd_req_pu_id_urands[713]  = 32'd4237076374;
    rd_req_pu_id_urands[714]  = 32'd144893350;
    rd_req_pu_id_urands[715]  = 32'd3095871817;
    rd_req_pu_id_urands[716]  = 32'd2498928479;
    rd_req_pu_id_urands[717]  = 32'd1558490347;
    rd_req_pu_id_urands[718]  = 32'd2169692153;
    rd_req_pu_id_urands[719]  = 32'd2639948476;
    rd_req_pu_id_urands[720]  = 32'd2074191474;
    rd_req_pu_id_urands[721]  = 32'd3911518463;
    rd_req_pu_id_urands[722]  = 32'd2303437051;
    rd_req_pu_id_urands[723]  = 32'd4201446912;
    rd_req_pu_id_urands[724]  = 32'd2455206431;
    rd_req_pu_id_urands[725]  = 32'd2777129223;
    rd_req_pu_id_urands[726]  = 32'd2319423012;
    rd_req_pu_id_urands[727]  = 32'd4031504842;
    rd_req_pu_id_urands[728]  = 32'd4032738740;
    rd_req_pu_id_urands[729]  = 32'd2470521885;
    rd_req_pu_id_urands[730]  = 32'd2104859651;
    rd_req_pu_id_urands[731]  = 32'd903790725;
    rd_req_pu_id_urands[732]  = 32'd3729337602;
    rd_req_pu_id_urands[733]  = 32'd2963855353;
    rd_req_pu_id_urands[734]  = 32'd3921038108;
    rd_req_pu_id_urands[735]  = 32'd2786685655;
    rd_req_pu_id_urands[736]  = 32'd1054937605;
    rd_req_pu_id_urands[737]  = 32'd410232301;
    rd_req_pu_id_urands[738]  = 32'd3959887719;
    rd_req_pu_id_urands[739]  = 32'd4170028202;
    rd_req_pu_id_urands[740]  = 32'd3607559556;
    rd_req_pu_id_urands[741]  = 32'd2991485570;
    rd_req_pu_id_urands[742]  = 32'd3134547111;
    rd_req_pu_id_urands[743]  = 32'd2077199703;
    rd_req_pu_id_urands[744]  = 32'd2645290693;
    rd_req_pu_id_urands[745]  = 32'd901892081;
    rd_req_pu_id_urands[746]  = 32'd2013538883;
    rd_req_pu_id_urands[747]  = 32'd2836028295;
    rd_req_pu_id_urands[748]  = 32'd2676704286;
    rd_req_pu_id_urands[749]  = 32'd1400961758;
    rd_req_pu_id_urands[750]  = 32'd832433304;
    rd_req_pu_id_urands[751]  = 32'd630486736;
    rd_req_pu_id_urands[752]  = 32'd3826361676;
    rd_req_pu_id_urands[753]  = 32'd4226887172;
    rd_req_pu_id_urands[754]  = 32'd440307736;
    rd_req_pu_id_urands[755]  = 32'd1237495462;
    rd_req_pu_id_urands[756]  = 32'd3949157205;
    rd_req_pu_id_urands[757]  = 32'd998220708;
    rd_req_pu_id_urands[758]  = 32'd2483995463;
    rd_req_pu_id_urands[759]  = 32'd1565621866;
    rd_req_pu_id_urands[760]  = 32'd3698300515;
    rd_req_pu_id_urands[761]  = 32'd1136417566;
    rd_req_pu_id_urands[762]  = 32'd2731857060;
    rd_req_pu_id_urands[763]  = 32'd4039472250;
    rd_req_pu_id_urands[764]  = 32'd1331161025;
    rd_req_pu_id_urands[765]  = 32'd3660567017;
    rd_req_pu_id_urands[766]  = 32'd4177959602;
    rd_req_pu_id_urands[767]  = 32'd1340215921;
    rd_req_pu_id_urands[768]  = 32'd1453707602;
    rd_req_pu_id_urands[769]  = 32'd1588942184;
    rd_req_pu_id_urands[770]  = 32'd4018372254;
    rd_req_pu_id_urands[771]  = 32'd1231754865;
    rd_req_pu_id_urands[772]  = 32'd4273804149;
    rd_req_pu_id_urands[773]  = 32'd4225775633;
    rd_req_pu_id_urands[774]  = 32'd1764162308;
    rd_req_pu_id_urands[775]  = 32'd1712245936;
    rd_req_pu_id_urands[776]  = 32'd271600657;
    rd_req_pu_id_urands[777]  = 32'd3746911726;
    rd_req_pu_id_urands[778]  = 32'd797493631;
    rd_req_pu_id_urands[779]  = 32'd1878624181;
    rd_req_pu_id_urands[780]  = 32'd2687615311;
    rd_req_pu_id_urands[781]  = 32'd2575095767;
    rd_req_pu_id_urands[782]  = 32'd1715711887;
    rd_req_pu_id_urands[783]  = 32'd2576463939;
    rd_req_pu_id_urands[784]  = 32'd4164967327;
    rd_req_pu_id_urands[785]  = 32'd2717490855;
    rd_req_pu_id_urands[786]  = 32'd2167959913;
    rd_req_pu_id_urands[787]  = 32'd1402843919;
    rd_req_pu_id_urands[788]  = 32'd3673833549;
    rd_req_pu_id_urands[789]  = 32'd740707736;
    rd_req_pu_id_urands[790]  = 32'd1939393384;
    rd_req_pu_id_urands[791]  = 32'd1345617167;
    rd_req_pu_id_urands[792]  = 32'd1008080356;
    rd_req_pu_id_urands[793]  = 32'd3497026556;
    rd_req_pu_id_urands[794]  = 32'd2670260538;
    rd_req_pu_id_urands[795]  = 32'd1413375473;
    rd_req_pu_id_urands[796]  = 32'd2279606152;
    rd_req_pu_id_urands[797]  = 32'd3597705098;
    rd_req_pu_id_urands[798]  = 32'd3961055637;
    rd_req_pu_id_urands[799]  = 32'd630644257;
    rd_req_pu_id_urands[800]  = 32'd2187534343;
    rd_req_pu_id_urands[801]  = 32'd949953951;
    rd_req_pu_id_urands[802]  = 32'd1328193797;
    rd_req_pu_id_urands[803]  = 32'd510195170;
    rd_req_pu_id_urands[804]  = 32'd492055056;
    rd_req_pu_id_urands[805]  = 32'd2235481182;
    rd_req_pu_id_urands[806]  = 32'd373300357;
    rd_req_pu_id_urands[807]  = 32'd2635750903;
    rd_req_pu_id_urands[808]  = 32'd2688111236;
    rd_req_pu_id_urands[809]  = 32'd2364559290;
    rd_req_pu_id_urands[810]  = 32'd282092751;
    rd_req_pu_id_urands[811]  = 32'd2566708882;
    rd_req_pu_id_urands[812]  = 32'd2582815419;
    rd_req_pu_id_urands[813]  = 32'd1609975385;
    rd_req_pu_id_urands[814]  = 32'd375798442;
    rd_req_pu_id_urands[815]  = 32'd3003909550;
    rd_req_pu_id_urands[816]  = 32'd1532902285;
    rd_req_pu_id_urands[817]  = 32'd142722424;
    rd_req_pu_id_urands[818]  = 32'd4249748325;
    rd_req_pu_id_urands[819]  = 32'd3739201203;
    rd_req_pu_id_urands[820]  = 32'd452908500;
    rd_req_pu_id_urands[821]  = 32'd167794619;
    rd_req_pu_id_urands[822]  = 32'd1337701049;
    rd_req_pu_id_urands[823]  = 32'd2526766739;
    rd_req_pu_id_urands[824]  = 32'd1150642578;
    rd_req_pu_id_urands[825]  = 32'd4084486046;
    rd_req_pu_id_urands[826]  = 32'd1941888071;
    rd_req_pu_id_urands[827]  = 32'd2976250866;
    rd_req_pu_id_urands[828]  = 32'd1061143550;
    rd_req_pu_id_urands[829]  = 32'd4235345521;
    rd_req_pu_id_urands[830]  = 32'd1537612880;
    rd_req_pu_id_urands[831]  = 32'd2637832717;
    rd_req_pu_id_urands[832]  = 32'd3649754950;
    rd_req_pu_id_urands[833]  = 32'd3464477717;
    rd_req_pu_id_urands[834]  = 32'd2098264329;
    rd_req_pu_id_urands[835]  = 32'd2526971317;
    rd_req_pu_id_urands[836]  = 32'd2305949611;
    rd_req_pu_id_urands[837]  = 32'd1128760871;
    rd_req_pu_id_urands[838]  = 32'd1576792884;
    rd_req_pu_id_urands[839]  = 32'd2189229087;
    rd_req_pu_id_urands[840]  = 32'd685187218;
    rd_req_pu_id_urands[841]  = 32'd3582255774;
    rd_req_pu_id_urands[842]  = 32'd934148564;
    rd_req_pu_id_urands[843]  = 32'd524911140;
    rd_req_pu_id_urands[844]  = 32'd1112534659;
    rd_req_pu_id_urands[845]  = 32'd3575835163;
    rd_req_pu_id_urands[846]  = 32'd3120318799;
    rd_req_pu_id_urands[847]  = 32'd3318930333;
    rd_req_pu_id_urands[848]  = 32'd171270650;
    rd_req_pu_id_urands[849]  = 32'd3644566281;
    rd_req_pu_id_urands[850]  = 32'd924006323;
    rd_req_pu_id_urands[851]  = 32'd2835406197;
    rd_req_pu_id_urands[852]  = 32'd888802297;
    rd_req_pu_id_urands[853]  = 32'd2530671868;
    rd_req_pu_id_urands[854]  = 32'd3631209966;
    rd_req_pu_id_urands[855]  = 32'd4206072862;
    rd_req_pu_id_urands[856]  = 32'd2666076294;
    rd_req_pu_id_urands[857]  = 32'd3988138348;
    rd_req_pu_id_urands[858]  = 32'd1821549799;
    rd_req_pu_id_urands[859]  = 32'd3178411504;
    rd_req_pu_id_urands[860]  = 32'd3254318879;
    rd_req_pu_id_urands[861]  = 32'd3775675336;
    rd_req_pu_id_urands[862]  = 32'd437196017;
    rd_req_pu_id_urands[863]  = 32'd2043333927;
    rd_req_pu_id_urands[864]  = 32'd984994483;
    rd_req_pu_id_urands[865]  = 32'd3440583940;
    rd_req_pu_id_urands[866]  = 32'd3106202822;
    rd_req_pu_id_urands[867]  = 32'd1278327491;
    rd_req_pu_id_urands[868]  = 32'd2001537281;
    rd_req_pu_id_urands[869]  = 32'd4203300164;
    rd_req_pu_id_urands[870]  = 32'd2201541435;
    rd_req_pu_id_urands[871]  = 32'd3810312735;
    rd_req_pu_id_urands[872]  = 32'd2865200591;
    rd_req_pu_id_urands[873]  = 32'd209490524;
    rd_req_pu_id_urands[874]  = 32'd3825946203;
    rd_req_pu_id_urands[875]  = 32'd57505114;
    rd_req_pu_id_urands[876]  = 32'd814858024;
    rd_req_pu_id_urands[877]  = 32'd3649304391;
    rd_req_pu_id_urands[878]  = 32'd37622349;
    rd_req_pu_id_urands[879]  = 32'd982449980;
    rd_req_pu_id_urands[880]  = 32'd3259563914;
    rd_req_pu_id_urands[881]  = 32'd338045757;
    rd_req_pu_id_urands[882]  = 32'd424630610;
    rd_req_pu_id_urands[883]  = 32'd1303973139;
    rd_req_pu_id_urands[884]  = 32'd1043831603;
    rd_req_pu_id_urands[885]  = 32'd4037593848;
    rd_req_pu_id_urands[886]  = 32'd3159648041;
    rd_req_pu_id_urands[887]  = 32'd3507385488;
    rd_req_pu_id_urands[888]  = 32'd2810023525;
    rd_req_pu_id_urands[889]  = 32'd2693760383;
    rd_req_pu_id_urands[890]  = 32'd2232307255;
    rd_req_pu_id_urands[891]  = 32'd2744370010;
    rd_req_pu_id_urands[892]  = 32'd579657422;
    rd_req_pu_id_urands[893]  = 32'd47573348;
    rd_req_pu_id_urands[894]  = 32'd3830127723;
    rd_req_pu_id_urands[895]  = 32'd1657747946;
    rd_req_pu_id_urands[896]  = 32'd3183729777;
    rd_req_pu_id_urands[897]  = 32'd3883045063;
    rd_req_pu_id_urands[898]  = 32'd3856912160;
    rd_req_pu_id_urands[899]  = 32'd3629581770;
    rd_req_pu_id_urands[900]  = 32'd2111297445;
    rd_req_pu_id_urands[901]  = 32'd2138956451;
    rd_req_pu_id_urands[902]  = 32'd3133857662;
    rd_req_pu_id_urands[903]  = 32'd1036322863;
    rd_req_pu_id_urands[904]  = 32'd3320434369;
    rd_req_pu_id_urands[905]  = 32'd196692902;
    rd_req_pu_id_urands[906]  = 32'd3380235644;
    rd_req_pu_id_urands[907]  = 32'd3481443647;
    rd_req_pu_id_urands[908]  = 32'd148833548;
    rd_req_pu_id_urands[909]  = 32'd1348175138;
    rd_req_pu_id_urands[910]  = 32'd3009001446;
    rd_req_pu_id_urands[911]  = 32'd4139503571;
    rd_req_pu_id_urands[912]  = 32'd3025646874;
    rd_req_pu_id_urands[913]  = 32'd3509434158;
    rd_req_pu_id_urands[914]  = 32'd156502223;
    rd_req_pu_id_urands[915]  = 32'd332574249;
    rd_req_pu_id_urands[916]  = 32'd3243904183;
    rd_req_pu_id_urands[917]  = 32'd3921292876;
    rd_req_pu_id_urands[918]  = 32'd4221629027;
    rd_req_pu_id_urands[919]  = 32'd3880859057;
    rd_req_pu_id_urands[920]  = 32'd3293744849;
    rd_req_pu_id_urands[921]  = 32'd1634340076;
    rd_req_pu_id_urands[922]  = 32'd2179145603;
    rd_req_pu_id_urands[923]  = 32'd1484024562;
    rd_req_pu_id_urands[924]  = 32'd4190488881;
    rd_req_pu_id_urands[925]  = 32'd1591157812;
    rd_req_pu_id_urands[926]  = 32'd1686533782;
    rd_req_pu_id_urands[927]  = 32'd3212590064;
    rd_req_pu_id_urands[928]  = 32'd938550216;
    rd_req_pu_id_urands[929]  = 32'd683336721;
    rd_req_pu_id_urands[930]  = 32'd110166749;
    rd_req_pu_id_urands[931]  = 32'd2091016727;
    rd_req_pu_id_urands[932]  = 32'd4097620692;
    rd_req_pu_id_urands[933]  = 32'd2235155360;
    rd_req_pu_id_urands[934]  = 32'd1983158959;
    rd_req_pu_id_urands[935]  = 32'd829807154;
    rd_req_pu_id_urands[936]  = 32'd1125697101;
    rd_req_pu_id_urands[937]  = 32'd562677285;
    rd_req_pu_id_urands[938]  = 32'd2386239342;
    rd_req_pu_id_urands[939]  = 32'd4095929086;
    rd_req_pu_id_urands[940]  = 32'd2137688371;
    rd_req_pu_id_urands[941]  = 32'd1364848683;
    rd_req_pu_id_urands[942]  = 32'd1879170436;
    rd_req_pu_id_urands[943]  = 32'd3971367210;
    rd_req_pu_id_urands[944]  = 32'd1331426926;
    rd_req_pu_id_urands[945]  = 32'd3343041632;
    rd_req_pu_id_urands[946]  = 32'd4175494287;
    rd_req_pu_id_urands[947]  = 32'd2556580846;
    rd_req_pu_id_urands[948]  = 32'd4053504340;
    rd_req_pu_id_urands[949]  = 32'd295468961;
    rd_req_pu_id_urands[950]  = 32'd2547129374;
    rd_req_pu_id_urands[951]  = 32'd2474967380;
    rd_req_pu_id_urands[952]  = 32'd2858518043;
    rd_req_pu_id_urands[953]  = 32'd1990724953;
    rd_req_pu_id_urands[954]  = 32'd1136403849;
    rd_req_pu_id_urands[955]  = 32'd3653662084;
    rd_req_pu_id_urands[956]  = 32'd91118043;
    rd_req_pu_id_urands[957]  = 32'd3640975360;
    rd_req_pu_id_urands[958]  = 32'd1390616595;
    rd_req_pu_id_urands[959]  = 32'd432473529;
    rd_req_pu_id_urands[960]  = 32'd1370901125;
    rd_req_pu_id_urands[961]  = 32'd2427605690;
    rd_req_pu_id_urands[962]  = 32'd3670643968;
    rd_req_pu_id_urands[963]  = 32'd1733198887;
    rd_req_pu_id_urands[964]  = 32'd367354171;
    rd_req_pu_id_urands[965]  = 32'd2147652374;
    rd_req_pu_id_urands[966]  = 32'd902821931;
    rd_req_pu_id_urands[967]  = 32'd1074087962;
    rd_req_pu_id_urands[968]  = 32'd860057731;
    rd_req_pu_id_urands[969]  = 32'd1839152733;
    rd_req_pu_id_urands[970]  = 32'd567495104;
    rd_req_pu_id_urands[971]  = 32'd941835725;
    rd_req_pu_id_urands[972]  = 32'd3638573827;
    rd_req_pu_id_urands[973]  = 32'd4132555665;
    rd_req_pu_id_urands[974]  = 32'd3178253497;
    rd_req_pu_id_urands[975]  = 32'd1103558980;
    rd_req_pu_id_urands[976]  = 32'd2035972843;
    rd_req_pu_id_urands[977]  = 32'd839648079;
    rd_req_pu_id_urands[978]  = 32'd867210096;
    rd_req_pu_id_urands[979]  = 32'd3205784455;
    rd_req_pu_id_urands[980]  = 32'd7222854;
    rd_req_pu_id_urands[981]  = 32'd3834055989;
    rd_req_pu_id_urands[982]  = 32'd975321992;
    rd_req_pu_id_urands[983]  = 32'd2221480095;
    rd_req_pu_id_urands[984]  = 32'd1203366316;
    rd_req_pu_id_urands[985]  = 32'd4082733489;
    rd_req_pu_id_urands[986]  = 32'd2753281454;
    rd_req_pu_id_urands[987]  = 32'd1501855616;
    rd_req_pu_id_urands[988]  = 32'd2585367008;
    rd_req_pu_id_urands[989]  = 32'd799549106;
    rd_req_pu_id_urands[990]  = 32'd3355627479;
    rd_req_pu_id_urands[991]  = 32'd500149957;
    rd_req_pu_id_urands[992]  = 32'd3391662124;
    rd_req_pu_id_urands[993]  = 32'd2051164125;
    rd_req_pu_id_urands[994]  = 32'd1743991407;
    rd_req_pu_id_urands[995]  = 32'd1850092980;
    rd_req_pu_id_urands[996]  = 32'd4049947021;
    rd_req_pu_id_urands[997]  = 32'd19630031;
    rd_req_pu_id_urands[998]  = 32'd1878623210;
    rd_req_pu_id_urands[999]  = 32'd519033017;

    rd_req_d_type_urands[0]    = 1'b0;
    rd_req_d_type_urands[1]    = 1'b0;
    rd_req_d_type_urands[2]    = 1'b1;
    rd_req_d_type_urands[3]    = 1'b1;
    rd_req_d_type_urands[4]    = 1'b1;
    rd_req_d_type_urands[5]    = 1'b1;
    rd_req_d_type_urands[6]    = 1'b1;
    rd_req_d_type_urands[7]    = 1'b0;
    rd_req_d_type_urands[8]    = 1'b1;
    rd_req_d_type_urands[9]    = 1'b1;
    rd_req_d_type_urands[10]   = 1'b0;
    rd_req_d_type_urands[11]   = 1'b1;
    rd_req_d_type_urands[12]   = 1'b0;
    rd_req_d_type_urands[13]   = 1'b1;
    rd_req_d_type_urands[14]   = 1'b0;
    rd_req_d_type_urands[15]   = 1'b1;
    rd_req_d_type_urands[16]   = 1'b0;
    rd_req_d_type_urands[17]   = 1'b0;
    rd_req_d_type_urands[18]   = 1'b0;
    rd_req_d_type_urands[19]   = 1'b1;
    rd_req_d_type_urands[20]   = 1'b0;
    rd_req_d_type_urands[21]   = 1'b0;
    rd_req_d_type_urands[22]   = 1'b0;
    rd_req_d_type_urands[23]   = 1'b1;
    rd_req_d_type_urands[24]   = 1'b0;
    rd_req_d_type_urands[25]   = 1'b0;
    rd_req_d_type_urands[26]   = 1'b0;
    rd_req_d_type_urands[27]   = 1'b0;
    rd_req_d_type_urands[28]   = 1'b0;
    rd_req_d_type_urands[29]   = 1'b1;
    rd_req_d_type_urands[30]   = 1'b1;
    rd_req_d_type_urands[31]   = 1'b1;
    rd_req_d_type_urands[32]   = 1'b0;
    rd_req_d_type_urands[33]   = 1'b0;
    rd_req_d_type_urands[34]   = 1'b1;
    rd_req_d_type_urands[35]   = 1'b0;
    rd_req_d_type_urands[36]   = 1'b0;
    rd_req_d_type_urands[37]   = 1'b1;
    rd_req_d_type_urands[38]   = 1'b0;
    rd_req_d_type_urands[39]   = 1'b0;
    rd_req_d_type_urands[40]   = 1'b1;
    rd_req_d_type_urands[41]   = 1'b0;
    rd_req_d_type_urands[42]   = 1'b0;
    rd_req_d_type_urands[43]   = 1'b1;
    rd_req_d_type_urands[44]   = 1'b1;
    rd_req_d_type_urands[45]   = 1'b0;
    rd_req_d_type_urands[46]   = 1'b1;
    rd_req_d_type_urands[47]   = 1'b0;
    rd_req_d_type_urands[48]   = 1'b1;
    rd_req_d_type_urands[49]   = 1'b1;
    rd_req_d_type_urands[50]   = 1'b0;
    rd_req_d_type_urands[51]   = 1'b1;
    rd_req_d_type_urands[52]   = 1'b0;
    rd_req_d_type_urands[53]   = 1'b0;
    rd_req_d_type_urands[54]   = 1'b0;
    rd_req_d_type_urands[55]   = 1'b0;
    rd_req_d_type_urands[56]   = 1'b1;
    rd_req_d_type_urands[57]   = 1'b1;
    rd_req_d_type_urands[58]   = 1'b0;
    rd_req_d_type_urands[59]   = 1'b0;
    rd_req_d_type_urands[60]   = 1'b1;
    rd_req_d_type_urands[61]   = 1'b1;
    rd_req_d_type_urands[62]   = 1'b1;
    rd_req_d_type_urands[63]   = 1'b1;
    rd_req_d_type_urands[64]   = 1'b0;
    rd_req_d_type_urands[65]   = 1'b1;
    rd_req_d_type_urands[66]   = 1'b1;
    rd_req_d_type_urands[67]   = 1'b1;
    rd_req_d_type_urands[68]   = 1'b0;
    rd_req_d_type_urands[69]   = 1'b1;
    rd_req_d_type_urands[70]   = 1'b0;
    rd_req_d_type_urands[71]   = 1'b1;
    rd_req_d_type_urands[72]   = 1'b1;
    rd_req_d_type_urands[73]   = 1'b1;
    rd_req_d_type_urands[74]   = 1'b1;
    rd_req_d_type_urands[75]   = 1'b0;
    rd_req_d_type_urands[76]   = 1'b0;
    rd_req_d_type_urands[77]   = 1'b1;
    rd_req_d_type_urands[78]   = 1'b1;
    rd_req_d_type_urands[79]   = 1'b1;
    rd_req_d_type_urands[80]   = 1'b0;
    rd_req_d_type_urands[81]   = 1'b1;
    rd_req_d_type_urands[82]   = 1'b0;
    rd_req_d_type_urands[83]   = 1'b0;
    rd_req_d_type_urands[84]   = 1'b0;
    rd_req_d_type_urands[85]   = 1'b1;
    rd_req_d_type_urands[86]   = 1'b0;
    rd_req_d_type_urands[87]   = 1'b0;
    rd_req_d_type_urands[88]   = 1'b1;
    rd_req_d_type_urands[89]   = 1'b0;
    rd_req_d_type_urands[90]   = 1'b0;
    rd_req_d_type_urands[91]   = 1'b1;
    rd_req_d_type_urands[92]   = 1'b0;
    rd_req_d_type_urands[93]   = 1'b0;
    rd_req_d_type_urands[94]   = 1'b0;
    rd_req_d_type_urands[95]   = 1'b1;
    rd_req_d_type_urands[96]   = 1'b0;
    rd_req_d_type_urands[97]   = 1'b1;
    rd_req_d_type_urands[98]   = 1'b0;
    rd_req_d_type_urands[99]   = 1'b1;
    rd_req_d_type_urands[100]  = 1'b1;
    rd_req_d_type_urands[101]  = 1'b1;
    rd_req_d_type_urands[102]  = 1'b1;
    rd_req_d_type_urands[103]  = 1'b0;
    rd_req_d_type_urands[104]  = 1'b0;
    rd_req_d_type_urands[105]  = 1'b1;
    rd_req_d_type_urands[106]  = 1'b0;
    rd_req_d_type_urands[107]  = 1'b0;
    rd_req_d_type_urands[108]  = 1'b1;
    rd_req_d_type_urands[109]  = 1'b0;
    rd_req_d_type_urands[110]  = 1'b1;
    rd_req_d_type_urands[111]  = 1'b0;
    rd_req_d_type_urands[112]  = 1'b0;
    rd_req_d_type_urands[113]  = 1'b0;
    rd_req_d_type_urands[114]  = 1'b1;
    rd_req_d_type_urands[115]  = 1'b1;
    rd_req_d_type_urands[116]  = 1'b1;
    rd_req_d_type_urands[117]  = 1'b0;
    rd_req_d_type_urands[118]  = 1'b1;
    rd_req_d_type_urands[119]  = 1'b1;
    rd_req_d_type_urands[120]  = 1'b1;
    rd_req_d_type_urands[121]  = 1'b0;
    rd_req_d_type_urands[122]  = 1'b1;
    rd_req_d_type_urands[123]  = 1'b1;
    rd_req_d_type_urands[124]  = 1'b0;
    rd_req_d_type_urands[125]  = 1'b1;
    rd_req_d_type_urands[126]  = 1'b1;
    rd_req_d_type_urands[127]  = 1'b1;
    rd_req_d_type_urands[128]  = 1'b0;
    rd_req_d_type_urands[129]  = 1'b0;
    rd_req_d_type_urands[130]  = 1'b0;
    rd_req_d_type_urands[131]  = 1'b0;
    rd_req_d_type_urands[132]  = 1'b1;
    rd_req_d_type_urands[133]  = 1'b0;
    rd_req_d_type_urands[134]  = 1'b1;
    rd_req_d_type_urands[135]  = 1'b0;
    rd_req_d_type_urands[136]  = 1'b0;
    rd_req_d_type_urands[137]  = 1'b1;
    rd_req_d_type_urands[138]  = 1'b1;
    rd_req_d_type_urands[139]  = 1'b0;
    rd_req_d_type_urands[140]  = 1'b0;
    rd_req_d_type_urands[141]  = 1'b0;
    rd_req_d_type_urands[142]  = 1'b1;
    rd_req_d_type_urands[143]  = 1'b0;
    rd_req_d_type_urands[144]  = 1'b0;
    rd_req_d_type_urands[145]  = 1'b0;
    rd_req_d_type_urands[146]  = 1'b1;
    rd_req_d_type_urands[147]  = 1'b0;
    rd_req_d_type_urands[148]  = 1'b0;
    rd_req_d_type_urands[149]  = 1'b1;
    rd_req_d_type_urands[150]  = 1'b0;
    rd_req_d_type_urands[151]  = 1'b0;
    rd_req_d_type_urands[152]  = 1'b1;
    rd_req_d_type_urands[153]  = 1'b0;
    rd_req_d_type_urands[154]  = 1'b1;
    rd_req_d_type_urands[155]  = 1'b1;
    rd_req_d_type_urands[156]  = 1'b1;
    rd_req_d_type_urands[157]  = 1'b1;
    rd_req_d_type_urands[158]  = 1'b0;
    rd_req_d_type_urands[159]  = 1'b0;
    rd_req_d_type_urands[160]  = 1'b1;
    rd_req_d_type_urands[161]  = 1'b1;
    rd_req_d_type_urands[162]  = 1'b0;
    rd_req_d_type_urands[163]  = 1'b0;
    rd_req_d_type_urands[164]  = 1'b1;
    rd_req_d_type_urands[165]  = 1'b1;
    rd_req_d_type_urands[166]  = 1'b1;
    rd_req_d_type_urands[167]  = 1'b1;
    rd_req_d_type_urands[168]  = 1'b0;
    rd_req_d_type_urands[169]  = 1'b0;
    rd_req_d_type_urands[170]  = 1'b0;
    rd_req_d_type_urands[171]  = 1'b0;
    rd_req_d_type_urands[172]  = 1'b0;
    rd_req_d_type_urands[173]  = 1'b1;
    rd_req_d_type_urands[174]  = 1'b0;
    rd_req_d_type_urands[175]  = 1'b1;
    rd_req_d_type_urands[176]  = 1'b1;
    rd_req_d_type_urands[177]  = 1'b1;
    rd_req_d_type_urands[178]  = 1'b1;
    rd_req_d_type_urands[179]  = 1'b1;
    rd_req_d_type_urands[180]  = 1'b1;
    rd_req_d_type_urands[181]  = 1'b1;
    rd_req_d_type_urands[182]  = 1'b0;
    rd_req_d_type_urands[183]  = 1'b1;
    rd_req_d_type_urands[184]  = 1'b1;
    rd_req_d_type_urands[185]  = 1'b0;
    rd_req_d_type_urands[186]  = 1'b0;
    rd_req_d_type_urands[187]  = 1'b1;
    rd_req_d_type_urands[188]  = 1'b1;
    rd_req_d_type_urands[189]  = 1'b1;
    rd_req_d_type_urands[190]  = 1'b0;
    rd_req_d_type_urands[191]  = 1'b1;
    rd_req_d_type_urands[192]  = 1'b1;
    rd_req_d_type_urands[193]  = 1'b1;
    rd_req_d_type_urands[194]  = 1'b1;
    rd_req_d_type_urands[195]  = 1'b0;
    rd_req_d_type_urands[196]  = 1'b1;
    rd_req_d_type_urands[197]  = 1'b1;
    rd_req_d_type_urands[198]  = 1'b1;
    rd_req_d_type_urands[199]  = 1'b0;
    rd_req_d_type_urands[200]  = 1'b1;
    rd_req_d_type_urands[201]  = 1'b1;
    rd_req_d_type_urands[202]  = 1'b1;
    rd_req_d_type_urands[203]  = 1'b1;
    rd_req_d_type_urands[204]  = 1'b0;
    rd_req_d_type_urands[205]  = 1'b1;
    rd_req_d_type_urands[206]  = 1'b1;
    rd_req_d_type_urands[207]  = 1'b0;
    rd_req_d_type_urands[208]  = 1'b0;
    rd_req_d_type_urands[209]  = 1'b0;
    rd_req_d_type_urands[210]  = 1'b1;
    rd_req_d_type_urands[211]  = 1'b0;
    rd_req_d_type_urands[212]  = 1'b1;
    rd_req_d_type_urands[213]  = 1'b0;
    rd_req_d_type_urands[214]  = 1'b1;
    rd_req_d_type_urands[215]  = 1'b0;
    rd_req_d_type_urands[216]  = 1'b0;
    rd_req_d_type_urands[217]  = 1'b1;
    rd_req_d_type_urands[218]  = 1'b0;
    rd_req_d_type_urands[219]  = 1'b0;
    rd_req_d_type_urands[220]  = 1'b0;
    rd_req_d_type_urands[221]  = 1'b1;
    rd_req_d_type_urands[222]  = 1'b0;
    rd_req_d_type_urands[223]  = 1'b1;
    rd_req_d_type_urands[224]  = 1'b0;
    rd_req_d_type_urands[225]  = 1'b1;
    rd_req_d_type_urands[226]  = 1'b1;
    rd_req_d_type_urands[227]  = 1'b1;
    rd_req_d_type_urands[228]  = 1'b1;
    rd_req_d_type_urands[229]  = 1'b1;
    rd_req_d_type_urands[230]  = 1'b1;
    rd_req_d_type_urands[231]  = 1'b1;
    rd_req_d_type_urands[232]  = 1'b1;
    rd_req_d_type_urands[233]  = 1'b1;
    rd_req_d_type_urands[234]  = 1'b1;
    rd_req_d_type_urands[235]  = 1'b1;
    rd_req_d_type_urands[236]  = 1'b0;
    rd_req_d_type_urands[237]  = 1'b0;
    rd_req_d_type_urands[238]  = 1'b0;
    rd_req_d_type_urands[239]  = 1'b1;
    rd_req_d_type_urands[240]  = 1'b1;
    rd_req_d_type_urands[241]  = 1'b1;
    rd_req_d_type_urands[242]  = 1'b0;
    rd_req_d_type_urands[243]  = 1'b1;
    rd_req_d_type_urands[244]  = 1'b1;
    rd_req_d_type_urands[245]  = 1'b0;
    rd_req_d_type_urands[246]  = 1'b1;
    rd_req_d_type_urands[247]  = 1'b1;
    rd_req_d_type_urands[248]  = 1'b0;
    rd_req_d_type_urands[249]  = 1'b1;
    rd_req_d_type_urands[250]  = 1'b0;
    rd_req_d_type_urands[251]  = 1'b1;
    rd_req_d_type_urands[252]  = 1'b0;
    rd_req_d_type_urands[253]  = 1'b0;
    rd_req_d_type_urands[254]  = 1'b0;
    rd_req_d_type_urands[255]  = 1'b0;
    rd_req_d_type_urands[256]  = 1'b0;
    rd_req_d_type_urands[257]  = 1'b1;
    rd_req_d_type_urands[258]  = 1'b0;
    rd_req_d_type_urands[259]  = 1'b0;
    rd_req_d_type_urands[260]  = 1'b1;
    rd_req_d_type_urands[261]  = 1'b1;
    rd_req_d_type_urands[262]  = 1'b0;
    rd_req_d_type_urands[263]  = 1'b0;
    rd_req_d_type_urands[264]  = 1'b0;
    rd_req_d_type_urands[265]  = 1'b1;
    rd_req_d_type_urands[266]  = 1'b0;
    rd_req_d_type_urands[267]  = 1'b1;
    rd_req_d_type_urands[268]  = 1'b1;
    rd_req_d_type_urands[269]  = 1'b0;
    rd_req_d_type_urands[270]  = 1'b1;
    rd_req_d_type_urands[271]  = 1'b0;
    rd_req_d_type_urands[272]  = 1'b0;
    rd_req_d_type_urands[273]  = 1'b0;
    rd_req_d_type_urands[274]  = 1'b1;
    rd_req_d_type_urands[275]  = 1'b1;
    rd_req_d_type_urands[276]  = 1'b1;
    rd_req_d_type_urands[277]  = 1'b1;
    rd_req_d_type_urands[278]  = 1'b0;
    rd_req_d_type_urands[279]  = 1'b0;
    rd_req_d_type_urands[280]  = 1'b0;
    rd_req_d_type_urands[281]  = 1'b1;
    rd_req_d_type_urands[282]  = 1'b0;
    rd_req_d_type_urands[283]  = 1'b0;
    rd_req_d_type_urands[284]  = 1'b0;
    rd_req_d_type_urands[285]  = 1'b0;
    rd_req_d_type_urands[286]  = 1'b0;
    rd_req_d_type_urands[287]  = 1'b1;
    rd_req_d_type_urands[288]  = 1'b0;
    rd_req_d_type_urands[289]  = 1'b1;
    rd_req_d_type_urands[290]  = 1'b0;
    rd_req_d_type_urands[291]  = 1'b1;
    rd_req_d_type_urands[292]  = 1'b0;
    rd_req_d_type_urands[293]  = 1'b1;
    rd_req_d_type_urands[294]  = 1'b0;
    rd_req_d_type_urands[295]  = 1'b0;
    rd_req_d_type_urands[296]  = 1'b0;
    rd_req_d_type_urands[297]  = 1'b0;
    rd_req_d_type_urands[298]  = 1'b1;
    rd_req_d_type_urands[299]  = 1'b0;
    rd_req_d_type_urands[300]  = 1'b0;
    rd_req_d_type_urands[301]  = 1'b0;
    rd_req_d_type_urands[302]  = 1'b1;
    rd_req_d_type_urands[303]  = 1'b0;
    rd_req_d_type_urands[304]  = 1'b0;
    rd_req_d_type_urands[305]  = 1'b0;
    rd_req_d_type_urands[306]  = 1'b1;
    rd_req_d_type_urands[307]  = 1'b1;
    rd_req_d_type_urands[308]  = 1'b1;
    rd_req_d_type_urands[309]  = 1'b0;
    rd_req_d_type_urands[310]  = 1'b0;
    rd_req_d_type_urands[311]  = 1'b0;
    rd_req_d_type_urands[312]  = 1'b0;
    rd_req_d_type_urands[313]  = 1'b1;
    rd_req_d_type_urands[314]  = 1'b0;
    rd_req_d_type_urands[315]  = 1'b1;
    rd_req_d_type_urands[316]  = 1'b1;
    rd_req_d_type_urands[317]  = 1'b1;
    rd_req_d_type_urands[318]  = 1'b1;
    rd_req_d_type_urands[319]  = 1'b1;
    rd_req_d_type_urands[320]  = 1'b0;
    rd_req_d_type_urands[321]  = 1'b0;
    rd_req_d_type_urands[322]  = 1'b1;
    rd_req_d_type_urands[323]  = 1'b0;
    rd_req_d_type_urands[324]  = 1'b0;
    rd_req_d_type_urands[325]  = 1'b0;
    rd_req_d_type_urands[326]  = 1'b1;
    rd_req_d_type_urands[327]  = 1'b1;
    rd_req_d_type_urands[328]  = 1'b0;
    rd_req_d_type_urands[329]  = 1'b0;
    rd_req_d_type_urands[330]  = 1'b1;
    rd_req_d_type_urands[331]  = 1'b1;
    rd_req_d_type_urands[332]  = 1'b0;
    rd_req_d_type_urands[333]  = 1'b0;
    rd_req_d_type_urands[334]  = 1'b1;
    rd_req_d_type_urands[335]  = 1'b1;
    rd_req_d_type_urands[336]  = 1'b0;
    rd_req_d_type_urands[337]  = 1'b1;
    rd_req_d_type_urands[338]  = 1'b1;
    rd_req_d_type_urands[339]  = 1'b1;
    rd_req_d_type_urands[340]  = 1'b0;
    rd_req_d_type_urands[341]  = 1'b1;
    rd_req_d_type_urands[342]  = 1'b0;
    rd_req_d_type_urands[343]  = 1'b0;
    rd_req_d_type_urands[344]  = 1'b1;
    rd_req_d_type_urands[345]  = 1'b1;
    rd_req_d_type_urands[346]  = 1'b0;
    rd_req_d_type_urands[347]  = 1'b1;
    rd_req_d_type_urands[348]  = 1'b1;
    rd_req_d_type_urands[349]  = 1'b0;
    rd_req_d_type_urands[350]  = 1'b0;
    rd_req_d_type_urands[351]  = 1'b0;
    rd_req_d_type_urands[352]  = 1'b1;
    rd_req_d_type_urands[353]  = 1'b1;
    rd_req_d_type_urands[354]  = 1'b0;
    rd_req_d_type_urands[355]  = 1'b0;
    rd_req_d_type_urands[356]  = 1'b0;
    rd_req_d_type_urands[357]  = 1'b1;
    rd_req_d_type_urands[358]  = 1'b0;
    rd_req_d_type_urands[359]  = 1'b0;
    rd_req_d_type_urands[360]  = 1'b1;
    rd_req_d_type_urands[361]  = 1'b1;
    rd_req_d_type_urands[362]  = 1'b0;
    rd_req_d_type_urands[363]  = 1'b1;
    rd_req_d_type_urands[364]  = 1'b1;
    rd_req_d_type_urands[365]  = 1'b0;
    rd_req_d_type_urands[366]  = 1'b0;
    rd_req_d_type_urands[367]  = 1'b0;
    rd_req_d_type_urands[368]  = 1'b1;
    rd_req_d_type_urands[369]  = 1'b0;
    rd_req_d_type_urands[370]  = 1'b0;
    rd_req_d_type_urands[371]  = 1'b1;
    rd_req_d_type_urands[372]  = 1'b1;
    rd_req_d_type_urands[373]  = 1'b0;
    rd_req_d_type_urands[374]  = 1'b0;
    rd_req_d_type_urands[375]  = 1'b0;
    rd_req_d_type_urands[376]  = 1'b1;
    rd_req_d_type_urands[377]  = 1'b1;
    rd_req_d_type_urands[378]  = 1'b0;
    rd_req_d_type_urands[379]  = 1'b1;
    rd_req_d_type_urands[380]  = 1'b0;
    rd_req_d_type_urands[381]  = 1'b1;
    rd_req_d_type_urands[382]  = 1'b0;
    rd_req_d_type_urands[383]  = 1'b1;
    rd_req_d_type_urands[384]  = 1'b1;
    rd_req_d_type_urands[385]  = 1'b1;
    rd_req_d_type_urands[386]  = 1'b1;
    rd_req_d_type_urands[387]  = 1'b1;
    rd_req_d_type_urands[388]  = 1'b0;
    rd_req_d_type_urands[389]  = 1'b0;
    rd_req_d_type_urands[390]  = 1'b0;
    rd_req_d_type_urands[391]  = 1'b0;
    rd_req_d_type_urands[392]  = 1'b1;
    rd_req_d_type_urands[393]  = 1'b0;
    rd_req_d_type_urands[394]  = 1'b0;
    rd_req_d_type_urands[395]  = 1'b1;
    rd_req_d_type_urands[396]  = 1'b1;
    rd_req_d_type_urands[397]  = 1'b1;
    rd_req_d_type_urands[398]  = 1'b1;
    rd_req_d_type_urands[399]  = 1'b0;
    rd_req_d_type_urands[400]  = 1'b0;
    rd_req_d_type_urands[401]  = 1'b0;
    rd_req_d_type_urands[402]  = 1'b1;
    rd_req_d_type_urands[403]  = 1'b0;
    rd_req_d_type_urands[404]  = 1'b1;
    rd_req_d_type_urands[405]  = 1'b1;
    rd_req_d_type_urands[406]  = 1'b0;
    rd_req_d_type_urands[407]  = 1'b0;
    rd_req_d_type_urands[408]  = 1'b1;
    rd_req_d_type_urands[409]  = 1'b1;
    rd_req_d_type_urands[410]  = 1'b1;
    rd_req_d_type_urands[411]  = 1'b0;
    rd_req_d_type_urands[412]  = 1'b0;
    rd_req_d_type_urands[413]  = 1'b1;
    rd_req_d_type_urands[414]  = 1'b1;
    rd_req_d_type_urands[415]  = 1'b1;
    rd_req_d_type_urands[416]  = 1'b0;
    rd_req_d_type_urands[417]  = 1'b0;
    rd_req_d_type_urands[418]  = 1'b0;
    rd_req_d_type_urands[419]  = 1'b0;
    rd_req_d_type_urands[420]  = 1'b1;
    rd_req_d_type_urands[421]  = 1'b1;
    rd_req_d_type_urands[422]  = 1'b0;
    rd_req_d_type_urands[423]  = 1'b1;
    rd_req_d_type_urands[424]  = 1'b0;
    rd_req_d_type_urands[425]  = 1'b1;
    rd_req_d_type_urands[426]  = 1'b0;
    rd_req_d_type_urands[427]  = 1'b1;
    rd_req_d_type_urands[428]  = 1'b0;
    rd_req_d_type_urands[429]  = 1'b1;
    rd_req_d_type_urands[430]  = 1'b1;
    rd_req_d_type_urands[431]  = 1'b0;
    rd_req_d_type_urands[432]  = 1'b0;
    rd_req_d_type_urands[433]  = 1'b0;
    rd_req_d_type_urands[434]  = 1'b0;
    rd_req_d_type_urands[435]  = 1'b0;
    rd_req_d_type_urands[436]  = 1'b1;
    rd_req_d_type_urands[437]  = 1'b1;
    rd_req_d_type_urands[438]  = 1'b1;
    rd_req_d_type_urands[439]  = 1'b1;
    rd_req_d_type_urands[440]  = 1'b0;
    rd_req_d_type_urands[441]  = 1'b0;
    rd_req_d_type_urands[442]  = 1'b0;
    rd_req_d_type_urands[443]  = 1'b0;
    rd_req_d_type_urands[444]  = 1'b0;
    rd_req_d_type_urands[445]  = 1'b1;
    rd_req_d_type_urands[446]  = 1'b1;
    rd_req_d_type_urands[447]  = 1'b0;
    rd_req_d_type_urands[448]  = 1'b0;
    rd_req_d_type_urands[449]  = 1'b1;
    rd_req_d_type_urands[450]  = 1'b0;
    rd_req_d_type_urands[451]  = 1'b0;
    rd_req_d_type_urands[452]  = 1'b0;
    rd_req_d_type_urands[453]  = 1'b1;
    rd_req_d_type_urands[454]  = 1'b1;
    rd_req_d_type_urands[455]  = 1'b1;
    rd_req_d_type_urands[456]  = 1'b1;
    rd_req_d_type_urands[457]  = 1'b0;
    rd_req_d_type_urands[458]  = 1'b0;
    rd_req_d_type_urands[459]  = 1'b1;
    rd_req_d_type_urands[460]  = 1'b1;
    rd_req_d_type_urands[461]  = 1'b1;
    rd_req_d_type_urands[462]  = 1'b0;
    rd_req_d_type_urands[463]  = 1'b0;
    rd_req_d_type_urands[464]  = 1'b0;
    rd_req_d_type_urands[465]  = 1'b0;
    rd_req_d_type_urands[466]  = 1'b0;
    rd_req_d_type_urands[467]  = 1'b0;
    rd_req_d_type_urands[468]  = 1'b0;
    rd_req_d_type_urands[469]  = 1'b0;
    rd_req_d_type_urands[470]  = 1'b1;
    rd_req_d_type_urands[471]  = 1'b1;
    rd_req_d_type_urands[472]  = 1'b0;
    rd_req_d_type_urands[473]  = 1'b0;
    rd_req_d_type_urands[474]  = 1'b1;
    rd_req_d_type_urands[475]  = 1'b1;
    rd_req_d_type_urands[476]  = 1'b1;
    rd_req_d_type_urands[477]  = 1'b1;
    rd_req_d_type_urands[478]  = 1'b1;
    rd_req_d_type_urands[479]  = 1'b0;
    rd_req_d_type_urands[480]  = 1'b1;
    rd_req_d_type_urands[481]  = 1'b1;
    rd_req_d_type_urands[482]  = 1'b1;
    rd_req_d_type_urands[483]  = 1'b1;
    rd_req_d_type_urands[484]  = 1'b1;
    rd_req_d_type_urands[485]  = 1'b1;
    rd_req_d_type_urands[486]  = 1'b0;
    rd_req_d_type_urands[487]  = 1'b1;
    rd_req_d_type_urands[488]  = 1'b1;
    rd_req_d_type_urands[489]  = 1'b1;
    rd_req_d_type_urands[490]  = 1'b0;
    rd_req_d_type_urands[491]  = 1'b1;
    rd_req_d_type_urands[492]  = 1'b0;
    rd_req_d_type_urands[493]  = 1'b0;
    rd_req_d_type_urands[494]  = 1'b1;
    rd_req_d_type_urands[495]  = 1'b0;
    rd_req_d_type_urands[496]  = 1'b1;
    rd_req_d_type_urands[497]  = 1'b1;
    rd_req_d_type_urands[498]  = 1'b0;
    rd_req_d_type_urands[499]  = 1'b1;
    rd_req_d_type_urands[500]  = 1'b1;
    rd_req_d_type_urands[501]  = 1'b1;
    rd_req_d_type_urands[502]  = 1'b0;
    rd_req_d_type_urands[503]  = 1'b1;
    rd_req_d_type_urands[504]  = 1'b1;
    rd_req_d_type_urands[505]  = 1'b1;
    rd_req_d_type_urands[506]  = 1'b1;
    rd_req_d_type_urands[507]  = 1'b1;
    rd_req_d_type_urands[508]  = 1'b0;
    rd_req_d_type_urands[509]  = 1'b1;
    rd_req_d_type_urands[510]  = 1'b0;
    rd_req_d_type_urands[511]  = 1'b0;
    rd_req_d_type_urands[512]  = 1'b0;
    rd_req_d_type_urands[513]  = 1'b0;
    rd_req_d_type_urands[514]  = 1'b1;
    rd_req_d_type_urands[515]  = 1'b0;
    rd_req_d_type_urands[516]  = 1'b1;
    rd_req_d_type_urands[517]  = 1'b1;
    rd_req_d_type_urands[518]  = 1'b1;
    rd_req_d_type_urands[519]  = 1'b0;
    rd_req_d_type_urands[520]  = 1'b0;
    rd_req_d_type_urands[521]  = 1'b0;
    rd_req_d_type_urands[522]  = 1'b0;
    rd_req_d_type_urands[523]  = 1'b1;
    rd_req_d_type_urands[524]  = 1'b0;
    rd_req_d_type_urands[525]  = 1'b0;
    rd_req_d_type_urands[526]  = 1'b0;
    rd_req_d_type_urands[527]  = 1'b1;
    rd_req_d_type_urands[528]  = 1'b1;
    rd_req_d_type_urands[529]  = 1'b1;
    rd_req_d_type_urands[530]  = 1'b0;
    rd_req_d_type_urands[531]  = 1'b1;
    rd_req_d_type_urands[532]  = 1'b1;
    rd_req_d_type_urands[533]  = 1'b0;
    rd_req_d_type_urands[534]  = 1'b0;
    rd_req_d_type_urands[535]  = 1'b1;
    rd_req_d_type_urands[536]  = 1'b1;
    rd_req_d_type_urands[537]  = 1'b1;
    rd_req_d_type_urands[538]  = 1'b1;
    rd_req_d_type_urands[539]  = 1'b0;
    rd_req_d_type_urands[540]  = 1'b0;
    rd_req_d_type_urands[541]  = 1'b1;
    rd_req_d_type_urands[542]  = 1'b0;
    rd_req_d_type_urands[543]  = 1'b0;
    rd_req_d_type_urands[544]  = 1'b0;
    rd_req_d_type_urands[545]  = 1'b1;
    rd_req_d_type_urands[546]  = 1'b0;
    rd_req_d_type_urands[547]  = 1'b0;
    rd_req_d_type_urands[548]  = 1'b1;
    rd_req_d_type_urands[549]  = 1'b1;
    rd_req_d_type_urands[550]  = 1'b1;
    rd_req_d_type_urands[551]  = 1'b1;
    rd_req_d_type_urands[552]  = 1'b1;
    rd_req_d_type_urands[553]  = 1'b1;
    rd_req_d_type_urands[554]  = 1'b1;
    rd_req_d_type_urands[555]  = 1'b1;
    rd_req_d_type_urands[556]  = 1'b0;
    rd_req_d_type_urands[557]  = 1'b0;
    rd_req_d_type_urands[558]  = 1'b1;
    rd_req_d_type_urands[559]  = 1'b0;
    rd_req_d_type_urands[560]  = 1'b0;
    rd_req_d_type_urands[561]  = 1'b1;
    rd_req_d_type_urands[562]  = 1'b0;
    rd_req_d_type_urands[563]  = 1'b0;
    rd_req_d_type_urands[564]  = 1'b0;
    rd_req_d_type_urands[565]  = 1'b0;
    rd_req_d_type_urands[566]  = 1'b0;
    rd_req_d_type_urands[567]  = 1'b0;
    rd_req_d_type_urands[568]  = 1'b1;
    rd_req_d_type_urands[569]  = 1'b0;
    rd_req_d_type_urands[570]  = 1'b0;
    rd_req_d_type_urands[571]  = 1'b0;
    rd_req_d_type_urands[572]  = 1'b0;
    rd_req_d_type_urands[573]  = 1'b1;
    rd_req_d_type_urands[574]  = 1'b0;
    rd_req_d_type_urands[575]  = 1'b1;
    rd_req_d_type_urands[576]  = 1'b0;
    rd_req_d_type_urands[577]  = 1'b1;
    rd_req_d_type_urands[578]  = 1'b0;
    rd_req_d_type_urands[579]  = 1'b1;
    rd_req_d_type_urands[580]  = 1'b1;
    rd_req_d_type_urands[581]  = 1'b0;
    rd_req_d_type_urands[582]  = 1'b1;
    rd_req_d_type_urands[583]  = 1'b0;
    rd_req_d_type_urands[584]  = 1'b1;
    rd_req_d_type_urands[585]  = 1'b0;
    rd_req_d_type_urands[586]  = 1'b1;
    rd_req_d_type_urands[587]  = 1'b0;
    rd_req_d_type_urands[588]  = 1'b0;
    rd_req_d_type_urands[589]  = 1'b1;
    rd_req_d_type_urands[590]  = 1'b1;
    rd_req_d_type_urands[591]  = 1'b1;
    rd_req_d_type_urands[592]  = 1'b1;
    rd_req_d_type_urands[593]  = 1'b0;
    rd_req_d_type_urands[594]  = 1'b1;
    rd_req_d_type_urands[595]  = 1'b1;
    rd_req_d_type_urands[596]  = 1'b0;
    rd_req_d_type_urands[597]  = 1'b0;
    rd_req_d_type_urands[598]  = 1'b0;
    rd_req_d_type_urands[599]  = 1'b1;
    rd_req_d_type_urands[600]  = 1'b1;
    rd_req_d_type_urands[601]  = 1'b1;
    rd_req_d_type_urands[602]  = 1'b0;
    rd_req_d_type_urands[603]  = 1'b1;
    rd_req_d_type_urands[604]  = 1'b0;
    rd_req_d_type_urands[605]  = 1'b1;
    rd_req_d_type_urands[606]  = 1'b1;
    rd_req_d_type_urands[607]  = 1'b1;
    rd_req_d_type_urands[608]  = 1'b1;
    rd_req_d_type_urands[609]  = 1'b1;
    rd_req_d_type_urands[610]  = 1'b0;
    rd_req_d_type_urands[611]  = 1'b1;
    rd_req_d_type_urands[612]  = 1'b0;
    rd_req_d_type_urands[613]  = 1'b0;
    rd_req_d_type_urands[614]  = 1'b0;
    rd_req_d_type_urands[615]  = 1'b0;
    rd_req_d_type_urands[616]  = 1'b1;
    rd_req_d_type_urands[617]  = 1'b0;
    rd_req_d_type_urands[618]  = 1'b0;
    rd_req_d_type_urands[619]  = 1'b1;
    rd_req_d_type_urands[620]  = 1'b1;
    rd_req_d_type_urands[621]  = 1'b1;
    rd_req_d_type_urands[622]  = 1'b1;
    rd_req_d_type_urands[623]  = 1'b1;
    rd_req_d_type_urands[624]  = 1'b1;
    rd_req_d_type_urands[625]  = 1'b1;
    rd_req_d_type_urands[626]  = 1'b0;
    rd_req_d_type_urands[627]  = 1'b0;
    rd_req_d_type_urands[628]  = 1'b1;
    rd_req_d_type_urands[629]  = 1'b0;
    rd_req_d_type_urands[630]  = 1'b1;
    rd_req_d_type_urands[631]  = 1'b0;
    rd_req_d_type_urands[632]  = 1'b0;
    rd_req_d_type_urands[633]  = 1'b1;
    rd_req_d_type_urands[634]  = 1'b0;
    rd_req_d_type_urands[635]  = 1'b0;
    rd_req_d_type_urands[636]  = 1'b0;
    rd_req_d_type_urands[637]  = 1'b1;
    rd_req_d_type_urands[638]  = 1'b0;
    rd_req_d_type_urands[639]  = 1'b1;
    rd_req_d_type_urands[640]  = 1'b1;
    rd_req_d_type_urands[641]  = 1'b0;
    rd_req_d_type_urands[642]  = 1'b1;
    rd_req_d_type_urands[643]  = 1'b1;
    rd_req_d_type_urands[644]  = 1'b1;
    rd_req_d_type_urands[645]  = 1'b1;
    rd_req_d_type_urands[646]  = 1'b1;
    rd_req_d_type_urands[647]  = 1'b0;
    rd_req_d_type_urands[648]  = 1'b1;
    rd_req_d_type_urands[649]  = 1'b1;
    rd_req_d_type_urands[650]  = 1'b1;
    rd_req_d_type_urands[651]  = 1'b0;
    rd_req_d_type_urands[652]  = 1'b0;
    rd_req_d_type_urands[653]  = 1'b0;
    rd_req_d_type_urands[654]  = 1'b0;
    rd_req_d_type_urands[655]  = 1'b0;
    rd_req_d_type_urands[656]  = 1'b1;
    rd_req_d_type_urands[657]  = 1'b0;
    rd_req_d_type_urands[658]  = 1'b1;
    rd_req_d_type_urands[659]  = 1'b1;
    rd_req_d_type_urands[660]  = 1'b0;
    rd_req_d_type_urands[661]  = 1'b0;
    rd_req_d_type_urands[662]  = 1'b0;
    rd_req_d_type_urands[663]  = 1'b0;
    rd_req_d_type_urands[664]  = 1'b1;
    rd_req_d_type_urands[665]  = 1'b1;
    rd_req_d_type_urands[666]  = 1'b1;
    rd_req_d_type_urands[667]  = 1'b1;
    rd_req_d_type_urands[668]  = 1'b0;
    rd_req_d_type_urands[669]  = 1'b1;
    rd_req_d_type_urands[670]  = 1'b1;
    rd_req_d_type_urands[671]  = 1'b0;
    rd_req_d_type_urands[672]  = 1'b1;
    rd_req_d_type_urands[673]  = 1'b0;
    rd_req_d_type_urands[674]  = 1'b0;
    rd_req_d_type_urands[675]  = 1'b0;
    rd_req_d_type_urands[676]  = 1'b1;
    rd_req_d_type_urands[677]  = 1'b0;
    rd_req_d_type_urands[678]  = 1'b0;
    rd_req_d_type_urands[679]  = 1'b1;
    rd_req_d_type_urands[680]  = 1'b1;
    rd_req_d_type_urands[681]  = 1'b0;
    rd_req_d_type_urands[682]  = 1'b0;
    rd_req_d_type_urands[683]  = 1'b1;
    rd_req_d_type_urands[684]  = 1'b0;
    rd_req_d_type_urands[685]  = 1'b0;
    rd_req_d_type_urands[686]  = 1'b0;
    rd_req_d_type_urands[687]  = 1'b0;
    rd_req_d_type_urands[688]  = 1'b0;
    rd_req_d_type_urands[689]  = 1'b1;
    rd_req_d_type_urands[690]  = 1'b1;
    rd_req_d_type_urands[691]  = 1'b1;
    rd_req_d_type_urands[692]  = 1'b1;
    rd_req_d_type_urands[693]  = 1'b0;
    rd_req_d_type_urands[694]  = 1'b1;
    rd_req_d_type_urands[695]  = 1'b1;
    rd_req_d_type_urands[696]  = 1'b0;
    rd_req_d_type_urands[697]  = 1'b1;
    rd_req_d_type_urands[698]  = 1'b0;
    rd_req_d_type_urands[699]  = 1'b1;
    rd_req_d_type_urands[700]  = 1'b0;
    rd_req_d_type_urands[701]  = 1'b1;
    rd_req_d_type_urands[702]  = 1'b1;
    rd_req_d_type_urands[703]  = 1'b1;
    rd_req_d_type_urands[704]  = 1'b0;
    rd_req_d_type_urands[705]  = 1'b1;
    rd_req_d_type_urands[706]  = 1'b0;
    rd_req_d_type_urands[707]  = 1'b0;
    rd_req_d_type_urands[708]  = 1'b0;
    rd_req_d_type_urands[709]  = 1'b0;
    rd_req_d_type_urands[710]  = 1'b1;
    rd_req_d_type_urands[711]  = 1'b1;
    rd_req_d_type_urands[712]  = 1'b1;
    rd_req_d_type_urands[713]  = 1'b1;
    rd_req_d_type_urands[714]  = 1'b1;
    rd_req_d_type_urands[715]  = 1'b1;
    rd_req_d_type_urands[716]  = 1'b0;
    rd_req_d_type_urands[717]  = 1'b0;
    rd_req_d_type_urands[718]  = 1'b0;
    rd_req_d_type_urands[719]  = 1'b0;
    rd_req_d_type_urands[720]  = 1'b0;
    rd_req_d_type_urands[721]  = 1'b0;
    rd_req_d_type_urands[722]  = 1'b0;
    rd_req_d_type_urands[723]  = 1'b1;
    rd_req_d_type_urands[724]  = 1'b1;
    rd_req_d_type_urands[725]  = 1'b1;
    rd_req_d_type_urands[726]  = 1'b0;
    rd_req_d_type_urands[727]  = 1'b0;
    rd_req_d_type_urands[728]  = 1'b0;
    rd_req_d_type_urands[729]  = 1'b0;
    rd_req_d_type_urands[730]  = 1'b1;
    rd_req_d_type_urands[731]  = 1'b1;
    rd_req_d_type_urands[732]  = 1'b0;
    rd_req_d_type_urands[733]  = 1'b0;
    rd_req_d_type_urands[734]  = 1'b0;
    rd_req_d_type_urands[735]  = 1'b1;
    rd_req_d_type_urands[736]  = 1'b1;
    rd_req_d_type_urands[737]  = 1'b1;
    rd_req_d_type_urands[738]  = 1'b1;
    rd_req_d_type_urands[739]  = 1'b0;
    rd_req_d_type_urands[740]  = 1'b1;
    rd_req_d_type_urands[741]  = 1'b1;
    rd_req_d_type_urands[742]  = 1'b1;
    rd_req_d_type_urands[743]  = 1'b1;
    rd_req_d_type_urands[744]  = 1'b1;
    rd_req_d_type_urands[745]  = 1'b1;
    rd_req_d_type_urands[746]  = 1'b1;
    rd_req_d_type_urands[747]  = 1'b0;
    rd_req_d_type_urands[748]  = 1'b0;
    rd_req_d_type_urands[749]  = 1'b0;
    rd_req_d_type_urands[750]  = 1'b0;
    rd_req_d_type_urands[751]  = 1'b1;
    rd_req_d_type_urands[752]  = 1'b1;
    rd_req_d_type_urands[753]  = 1'b0;
    rd_req_d_type_urands[754]  = 1'b0;
    rd_req_d_type_urands[755]  = 1'b1;
    rd_req_d_type_urands[756]  = 1'b1;
    rd_req_d_type_urands[757]  = 1'b0;
    rd_req_d_type_urands[758]  = 1'b0;
    rd_req_d_type_urands[759]  = 1'b0;
    rd_req_d_type_urands[760]  = 1'b0;
    rd_req_d_type_urands[761]  = 1'b1;
    rd_req_d_type_urands[762]  = 1'b0;
    rd_req_d_type_urands[763]  = 1'b1;
    rd_req_d_type_urands[764]  = 1'b0;
    rd_req_d_type_urands[765]  = 1'b0;
    rd_req_d_type_urands[766]  = 1'b1;
    rd_req_d_type_urands[767]  = 1'b0;
    rd_req_d_type_urands[768]  = 1'b1;
    rd_req_d_type_urands[769]  = 1'b0;
    rd_req_d_type_urands[770]  = 1'b1;
    rd_req_d_type_urands[771]  = 1'b0;
    rd_req_d_type_urands[772]  = 1'b0;
    rd_req_d_type_urands[773]  = 1'b0;
    rd_req_d_type_urands[774]  = 1'b1;
    rd_req_d_type_urands[775]  = 1'b0;
    rd_req_d_type_urands[776]  = 1'b0;
    rd_req_d_type_urands[777]  = 1'b0;
    rd_req_d_type_urands[778]  = 1'b1;
    rd_req_d_type_urands[779]  = 1'b0;
    rd_req_d_type_urands[780]  = 1'b1;
    rd_req_d_type_urands[781]  = 1'b1;
    rd_req_d_type_urands[782]  = 1'b1;
    rd_req_d_type_urands[783]  = 1'b1;
    rd_req_d_type_urands[784]  = 1'b1;
    rd_req_d_type_urands[785]  = 1'b0;
    rd_req_d_type_urands[786]  = 1'b1;
    rd_req_d_type_urands[787]  = 1'b1;
    rd_req_d_type_urands[788]  = 1'b1;
    rd_req_d_type_urands[789]  = 1'b0;
    rd_req_d_type_urands[790]  = 1'b1;
    rd_req_d_type_urands[791]  = 1'b0;
    rd_req_d_type_urands[792]  = 1'b1;
    rd_req_d_type_urands[793]  = 1'b0;
    rd_req_d_type_urands[794]  = 1'b1;
    rd_req_d_type_urands[795]  = 1'b1;
    rd_req_d_type_urands[796]  = 1'b1;
    rd_req_d_type_urands[797]  = 1'b0;
    rd_req_d_type_urands[798]  = 1'b1;
    rd_req_d_type_urands[799]  = 1'b1;
    rd_req_d_type_urands[800]  = 1'b1;
    rd_req_d_type_urands[801]  = 1'b0;
    rd_req_d_type_urands[802]  = 1'b0;
    rd_req_d_type_urands[803]  = 1'b0;
    rd_req_d_type_urands[804]  = 1'b0;
    rd_req_d_type_urands[805]  = 1'b1;
    rd_req_d_type_urands[806]  = 1'b0;
    rd_req_d_type_urands[807]  = 1'b0;
    rd_req_d_type_urands[808]  = 1'b0;
    rd_req_d_type_urands[809]  = 1'b1;
    rd_req_d_type_urands[810]  = 1'b1;
    rd_req_d_type_urands[811]  = 1'b1;
    rd_req_d_type_urands[812]  = 1'b1;
    rd_req_d_type_urands[813]  = 1'b0;
    rd_req_d_type_urands[814]  = 1'b1;
    rd_req_d_type_urands[815]  = 1'b0;
    rd_req_d_type_urands[816]  = 1'b1;
    rd_req_d_type_urands[817]  = 1'b0;
    rd_req_d_type_urands[818]  = 1'b1;
    rd_req_d_type_urands[819]  = 1'b1;
    rd_req_d_type_urands[820]  = 1'b0;
    rd_req_d_type_urands[821]  = 1'b0;
    rd_req_d_type_urands[822]  = 1'b1;
    rd_req_d_type_urands[823]  = 1'b0;
    rd_req_d_type_urands[824]  = 1'b0;
    rd_req_d_type_urands[825]  = 1'b1;
    rd_req_d_type_urands[826]  = 1'b1;
    rd_req_d_type_urands[827]  = 1'b0;
    rd_req_d_type_urands[828]  = 1'b1;
    rd_req_d_type_urands[829]  = 1'b1;
    rd_req_d_type_urands[830]  = 1'b1;
    rd_req_d_type_urands[831]  = 1'b0;
    rd_req_d_type_urands[832]  = 1'b1;
    rd_req_d_type_urands[833]  = 1'b1;
    rd_req_d_type_urands[834]  = 1'b1;
    rd_req_d_type_urands[835]  = 1'b1;
    rd_req_d_type_urands[836]  = 1'b1;
    rd_req_d_type_urands[837]  = 1'b1;
    rd_req_d_type_urands[838]  = 1'b0;
    rd_req_d_type_urands[839]  = 1'b1;
    rd_req_d_type_urands[840]  = 1'b1;
    rd_req_d_type_urands[841]  = 1'b0;
    rd_req_d_type_urands[842]  = 1'b0;
    rd_req_d_type_urands[843]  = 1'b0;
    rd_req_d_type_urands[844]  = 1'b0;
    rd_req_d_type_urands[845]  = 1'b0;
    rd_req_d_type_urands[846]  = 1'b1;
    rd_req_d_type_urands[847]  = 1'b0;
    rd_req_d_type_urands[848]  = 1'b1;
    rd_req_d_type_urands[849]  = 1'b1;
    rd_req_d_type_urands[850]  = 1'b1;
    rd_req_d_type_urands[851]  = 1'b0;
    rd_req_d_type_urands[852]  = 1'b1;
    rd_req_d_type_urands[853]  = 1'b0;
    rd_req_d_type_urands[854]  = 1'b1;
    rd_req_d_type_urands[855]  = 1'b1;
    rd_req_d_type_urands[856]  = 1'b1;
    rd_req_d_type_urands[857]  = 1'b1;
    rd_req_d_type_urands[858]  = 1'b1;
    rd_req_d_type_urands[859]  = 1'b1;
    rd_req_d_type_urands[860]  = 1'b1;
    rd_req_d_type_urands[861]  = 1'b1;
    rd_req_d_type_urands[862]  = 1'b0;
    rd_req_d_type_urands[863]  = 1'b1;
    rd_req_d_type_urands[864]  = 1'b1;
    rd_req_d_type_urands[865]  = 1'b0;
    rd_req_d_type_urands[866]  = 1'b1;
    rd_req_d_type_urands[867]  = 1'b0;
    rd_req_d_type_urands[868]  = 1'b0;
    rd_req_d_type_urands[869]  = 1'b1;
    rd_req_d_type_urands[870]  = 1'b1;
    rd_req_d_type_urands[871]  = 1'b1;
    rd_req_d_type_urands[872]  = 1'b1;
    rd_req_d_type_urands[873]  = 1'b1;
    rd_req_d_type_urands[874]  = 1'b1;
    rd_req_d_type_urands[875]  = 1'b0;
    rd_req_d_type_urands[876]  = 1'b0;
    rd_req_d_type_urands[877]  = 1'b1;
    rd_req_d_type_urands[878]  = 1'b1;
    rd_req_d_type_urands[879]  = 1'b1;
    rd_req_d_type_urands[880]  = 1'b0;
    rd_req_d_type_urands[881]  = 1'b1;
    rd_req_d_type_urands[882]  = 1'b1;
    rd_req_d_type_urands[883]  = 1'b0;
    rd_req_d_type_urands[884]  = 1'b0;
    rd_req_d_type_urands[885]  = 1'b0;
    rd_req_d_type_urands[886]  = 1'b1;
    rd_req_d_type_urands[887]  = 1'b0;
    rd_req_d_type_urands[888]  = 1'b1;
    rd_req_d_type_urands[889]  = 1'b0;
    rd_req_d_type_urands[890]  = 1'b0;
    rd_req_d_type_urands[891]  = 1'b1;
    rd_req_d_type_urands[892]  = 1'b1;
    rd_req_d_type_urands[893]  = 1'b0;
    rd_req_d_type_urands[894]  = 1'b0;
    rd_req_d_type_urands[895]  = 1'b1;
    rd_req_d_type_urands[896]  = 1'b1;
    rd_req_d_type_urands[897]  = 1'b0;
    rd_req_d_type_urands[898]  = 1'b1;
    rd_req_d_type_urands[899]  = 1'b1;
    rd_req_d_type_urands[900]  = 1'b0;
    rd_req_d_type_urands[901]  = 1'b1;
    rd_req_d_type_urands[902]  = 1'b0;
    rd_req_d_type_urands[903]  = 1'b1;
    rd_req_d_type_urands[904]  = 1'b0;
    rd_req_d_type_urands[905]  = 1'b1;
    rd_req_d_type_urands[906]  = 1'b0;
    rd_req_d_type_urands[907]  = 1'b1;
    rd_req_d_type_urands[908]  = 1'b1;
    rd_req_d_type_urands[909]  = 1'b0;
    rd_req_d_type_urands[910]  = 1'b0;
    rd_req_d_type_urands[911]  = 1'b0;
    rd_req_d_type_urands[912]  = 1'b0;
    rd_req_d_type_urands[913]  = 1'b1;
    rd_req_d_type_urands[914]  = 1'b1;
    rd_req_d_type_urands[915]  = 1'b1;
    rd_req_d_type_urands[916]  = 1'b0;
    rd_req_d_type_urands[917]  = 1'b0;
    rd_req_d_type_urands[918]  = 1'b0;
    rd_req_d_type_urands[919]  = 1'b1;
    rd_req_d_type_urands[920]  = 1'b1;
    rd_req_d_type_urands[921]  = 1'b1;
    rd_req_d_type_urands[922]  = 1'b1;
    rd_req_d_type_urands[923]  = 1'b1;
    rd_req_d_type_urands[924]  = 1'b0;
    rd_req_d_type_urands[925]  = 1'b0;
    rd_req_d_type_urands[926]  = 1'b0;
    rd_req_d_type_urands[927]  = 1'b1;
    rd_req_d_type_urands[928]  = 1'b1;
    rd_req_d_type_urands[929]  = 1'b0;
    rd_req_d_type_urands[930]  = 1'b1;
    rd_req_d_type_urands[931]  = 1'b1;
    rd_req_d_type_urands[932]  = 1'b1;
    rd_req_d_type_urands[933]  = 1'b1;
    rd_req_d_type_urands[934]  = 1'b1;
    rd_req_d_type_urands[935]  = 1'b1;
    rd_req_d_type_urands[936]  = 1'b1;
    rd_req_d_type_urands[937]  = 1'b1;
    rd_req_d_type_urands[938]  = 1'b0;
    rd_req_d_type_urands[939]  = 1'b0;
    rd_req_d_type_urands[940]  = 1'b0;
    rd_req_d_type_urands[941]  = 1'b0;
    rd_req_d_type_urands[942]  = 1'b1;
    rd_req_d_type_urands[943]  = 1'b0;
    rd_req_d_type_urands[944]  = 1'b0;
    rd_req_d_type_urands[945]  = 1'b0;
    rd_req_d_type_urands[946]  = 1'b0;
    rd_req_d_type_urands[947]  = 1'b1;
    rd_req_d_type_urands[948]  = 1'b1;
    rd_req_d_type_urands[949]  = 1'b1;
    rd_req_d_type_urands[950]  = 1'b0;
    rd_req_d_type_urands[951]  = 1'b0;
    rd_req_d_type_urands[952]  = 1'b1;
    rd_req_d_type_urands[953]  = 1'b0;
    rd_req_d_type_urands[954]  = 1'b1;
    rd_req_d_type_urands[955]  = 1'b1;
    rd_req_d_type_urands[956]  = 1'b1;
    rd_req_d_type_urands[957]  = 1'b1;
    rd_req_d_type_urands[958]  = 1'b1;
    rd_req_d_type_urands[959]  = 1'b1;
    rd_req_d_type_urands[960]  = 1'b1;
    rd_req_d_type_urands[961]  = 1'b0;
    rd_req_d_type_urands[962]  = 1'b0;
    rd_req_d_type_urands[963]  = 1'b1;
    rd_req_d_type_urands[964]  = 1'b0;
    rd_req_d_type_urands[965]  = 1'b0;
    rd_req_d_type_urands[966]  = 1'b0;
    rd_req_d_type_urands[967]  = 1'b1;
    rd_req_d_type_urands[968]  = 1'b0;
    rd_req_d_type_urands[969]  = 1'b0;
    rd_req_d_type_urands[970]  = 1'b1;
    rd_req_d_type_urands[971]  = 1'b0;
    rd_req_d_type_urands[972]  = 1'b0;
    rd_req_d_type_urands[973]  = 1'b1;
    rd_req_d_type_urands[974]  = 1'b1;
    rd_req_d_type_urands[975]  = 1'b1;
    rd_req_d_type_urands[976]  = 1'b0;
    rd_req_d_type_urands[977]  = 1'b1;
    rd_req_d_type_urands[978]  = 1'b0;
    rd_req_d_type_urands[979]  = 1'b0;
    rd_req_d_type_urands[980]  = 1'b1;
    rd_req_d_type_urands[981]  = 1'b1;
    rd_req_d_type_urands[982]  = 1'b0;
    rd_req_d_type_urands[983]  = 1'b1;
    rd_req_d_type_urands[984]  = 1'b0;
    rd_req_d_type_urands[985]  = 1'b0;
    rd_req_d_type_urands[986]  = 1'b0;
    rd_req_d_type_urands[987]  = 1'b1;
    rd_req_d_type_urands[988]  = 1'b1;
    rd_req_d_type_urands[989]  = 1'b0;
    rd_req_d_type_urands[990]  = 1'b1;
    rd_req_d_type_urands[991]  = 1'b1;
    rd_req_d_type_urands[992]  = 1'b1;
    rd_req_d_type_urands[993]  = 1'b1;
    rd_req_d_type_urands[994]  = 1'b1;
    rd_req_d_type_urands[995]  = 1'b0;
    rd_req_d_type_urands[996]  = 1'b0;
    rd_req_d_type_urands[997]  = 1'b0;
    rd_req_d_type_urands[998]  = 1'b0;
    rd_req_d_type_urands[999]  = 1'b1;

    inbuf_empty_rands[0]    = 1'b1;
    inbuf_empty_rands[1]    = 1'b1;
    inbuf_empty_rands[2]    = 1'b1;
    inbuf_empty_rands[3]    = 1'b0;
    inbuf_empty_rands[4]    = 1'b1;
    inbuf_empty_rands[5]    = 1'b0;
    inbuf_empty_rands[6]    = 1'b0;
    inbuf_empty_rands[7]    = 1'b1;
    inbuf_empty_rands[8]    = 1'b1;
    inbuf_empty_rands[9]    = 1'b0;
    inbuf_empty_rands[10]   = 1'b1;
    inbuf_empty_rands[11]   = 1'b0;
    inbuf_empty_rands[12]   = 1'b1;
    inbuf_empty_rands[13]   = 1'b0;
    inbuf_empty_rands[14]   = 1'b0;
    inbuf_empty_rands[15]   = 1'b1;
    inbuf_empty_rands[16]   = 1'b0;
    inbuf_empty_rands[17]   = 1'b1;
    inbuf_empty_rands[18]   = 1'b1;
    inbuf_empty_rands[19]   = 1'b0;
    inbuf_empty_rands[20]   = 1'b0;
    inbuf_empty_rands[21]   = 1'b0;
    inbuf_empty_rands[22]   = 1'b1;
    inbuf_empty_rands[23]   = 1'b1;
    inbuf_empty_rands[24]   = 1'b0;
    inbuf_empty_rands[25]   = 1'b1;
    inbuf_empty_rands[26]   = 1'b0;
    inbuf_empty_rands[27]   = 1'b0;
    inbuf_empty_rands[28]   = 1'b1;
    inbuf_empty_rands[29]   = 1'b1;
    inbuf_empty_rands[30]   = 1'b0;
    inbuf_empty_rands[31]   = 1'b1;
    inbuf_empty_rands[32]   = 1'b0;
    inbuf_empty_rands[33]   = 1'b0;
    inbuf_empty_rands[34]   = 1'b1;
    inbuf_empty_rands[35]   = 1'b0;
    inbuf_empty_rands[36]   = 1'b1;
    inbuf_empty_rands[37]   = 1'b1;
    inbuf_empty_rands[38]   = 1'b0;
    inbuf_empty_rands[39]   = 1'b1;
    inbuf_empty_rands[40]   = 1'b0;
    inbuf_empty_rands[41]   = 1'b1;
    inbuf_empty_rands[42]   = 1'b1;
    inbuf_empty_rands[43]   = 1'b0;
    inbuf_empty_rands[44]   = 1'b0;
    inbuf_empty_rands[45]   = 1'b0;
    inbuf_empty_rands[46]   = 1'b1;
    inbuf_empty_rands[47]   = 1'b1;
    inbuf_empty_rands[48]   = 1'b1;
    inbuf_empty_rands[49]   = 1'b1;
    inbuf_empty_rands[50]   = 1'b1;
    inbuf_empty_rands[51]   = 1'b1;
    inbuf_empty_rands[52]   = 1'b1;
    inbuf_empty_rands[53]   = 1'b0;
    inbuf_empty_rands[54]   = 1'b0;
    inbuf_empty_rands[55]   = 1'b0;
    inbuf_empty_rands[56]   = 1'b1;
    inbuf_empty_rands[57]   = 1'b0;
    inbuf_empty_rands[58]   = 1'b1;
    inbuf_empty_rands[59]   = 1'b0;
    inbuf_empty_rands[60]   = 1'b0;
    inbuf_empty_rands[61]   = 1'b0;
    inbuf_empty_rands[62]   = 1'b1;
    inbuf_empty_rands[63]   = 1'b0;
    inbuf_empty_rands[64]   = 1'b0;
    inbuf_empty_rands[65]   = 1'b0;
    inbuf_empty_rands[66]   = 1'b0;
    inbuf_empty_rands[67]   = 1'b1;
    inbuf_empty_rands[68]   = 1'b0;
    inbuf_empty_rands[69]   = 1'b0;
    inbuf_empty_rands[70]   = 1'b0;
    inbuf_empty_rands[71]   = 1'b0;
    inbuf_empty_rands[72]   = 1'b1;
    inbuf_empty_rands[73]   = 1'b0;
    inbuf_empty_rands[74]   = 1'b0;
    inbuf_empty_rands[75]   = 1'b0;
    inbuf_empty_rands[76]   = 1'b1;
    inbuf_empty_rands[77]   = 1'b1;
    inbuf_empty_rands[78]   = 1'b0;
    inbuf_empty_rands[79]   = 1'b0;
    inbuf_empty_rands[80]   = 1'b0;
    inbuf_empty_rands[81]   = 1'b1;
    inbuf_empty_rands[82]   = 1'b1;
    inbuf_empty_rands[83]   = 1'b1;
    inbuf_empty_rands[84]   = 1'b0;
    inbuf_empty_rands[85]   = 1'b0;
    inbuf_empty_rands[86]   = 1'b0;
    inbuf_empty_rands[87]   = 1'b1;
    inbuf_empty_rands[88]   = 1'b0;
    inbuf_empty_rands[89]   = 1'b0;
    inbuf_empty_rands[90]   = 1'b1;
    inbuf_empty_rands[91]   = 1'b0;
    inbuf_empty_rands[92]   = 1'b0;
    inbuf_empty_rands[93]   = 1'b0;
    inbuf_empty_rands[94]   = 1'b1;
    inbuf_empty_rands[95]   = 1'b0;
    inbuf_empty_rands[96]   = 1'b0;
    inbuf_empty_rands[97]   = 1'b0;
    inbuf_empty_rands[98]   = 1'b1;
    inbuf_empty_rands[99]   = 1'b0;
    inbuf_empty_rands[100]  = 1'b1;
    inbuf_empty_rands[101]  = 1'b1;
    inbuf_empty_rands[102]  = 1'b0;
    inbuf_empty_rands[103]  = 1'b0;
    inbuf_empty_rands[104]  = 1'b0;
    inbuf_empty_rands[105]  = 1'b1;
    inbuf_empty_rands[106]  = 1'b1;
    inbuf_empty_rands[107]  = 1'b1;
    inbuf_empty_rands[108]  = 1'b1;
    inbuf_empty_rands[109]  = 1'b0;
    inbuf_empty_rands[110]  = 1'b0;
    inbuf_empty_rands[111]  = 1'b0;
    inbuf_empty_rands[112]  = 1'b0;
    inbuf_empty_rands[113]  = 1'b1;
    inbuf_empty_rands[114]  = 1'b0;
    inbuf_empty_rands[115]  = 1'b1;
    inbuf_empty_rands[116]  = 1'b0;
    inbuf_empty_rands[117]  = 1'b0;
    inbuf_empty_rands[118]  = 1'b1;
    inbuf_empty_rands[119]  = 1'b1;
    inbuf_empty_rands[120]  = 1'b1;
    inbuf_empty_rands[121]  = 1'b1;
    inbuf_empty_rands[122]  = 1'b1;
    inbuf_empty_rands[123]  = 1'b1;
    inbuf_empty_rands[124]  = 1'b0;
    inbuf_empty_rands[125]  = 1'b0;
    inbuf_empty_rands[126]  = 1'b0;
    inbuf_empty_rands[127]  = 1'b0;
    inbuf_empty_rands[128]  = 1'b0;
    inbuf_empty_rands[129]  = 1'b1;
    inbuf_empty_rands[130]  = 1'b1;
    inbuf_empty_rands[131]  = 1'b1;
    inbuf_empty_rands[132]  = 1'b1;
    inbuf_empty_rands[133]  = 1'b1;
    inbuf_empty_rands[134]  = 1'b0;
    inbuf_empty_rands[135]  = 1'b1;
    inbuf_empty_rands[136]  = 1'b0;
    inbuf_empty_rands[137]  = 1'b0;
    inbuf_empty_rands[138]  = 1'b1;
    inbuf_empty_rands[139]  = 1'b0;
    inbuf_empty_rands[140]  = 1'b0;
    inbuf_empty_rands[141]  = 1'b0;
    inbuf_empty_rands[142]  = 1'b1;
    inbuf_empty_rands[143]  = 1'b0;
    inbuf_empty_rands[144]  = 1'b0;
    inbuf_empty_rands[145]  = 1'b0;
    inbuf_empty_rands[146]  = 1'b0;
    inbuf_empty_rands[147]  = 1'b1;
    inbuf_empty_rands[148]  = 1'b1;
    inbuf_empty_rands[149]  = 1'b1;
    inbuf_empty_rands[150]  = 1'b0;
    inbuf_empty_rands[151]  = 1'b0;
    inbuf_empty_rands[152]  = 1'b1;
    inbuf_empty_rands[153]  = 1'b1;
    inbuf_empty_rands[154]  = 1'b1;
    inbuf_empty_rands[155]  = 1'b1;
    inbuf_empty_rands[156]  = 1'b1;
    inbuf_empty_rands[157]  = 1'b1;
    inbuf_empty_rands[158]  = 1'b1;
    inbuf_empty_rands[159]  = 1'b0;
    inbuf_empty_rands[160]  = 1'b0;
    inbuf_empty_rands[161]  = 1'b1;
    inbuf_empty_rands[162]  = 1'b1;
    inbuf_empty_rands[163]  = 1'b0;
    inbuf_empty_rands[164]  = 1'b0;
    inbuf_empty_rands[165]  = 1'b0;
    inbuf_empty_rands[166]  = 1'b0;
    inbuf_empty_rands[167]  = 1'b1;
    inbuf_empty_rands[168]  = 1'b1;
    inbuf_empty_rands[169]  = 1'b1;
    inbuf_empty_rands[170]  = 1'b0;
    inbuf_empty_rands[171]  = 1'b0;
    inbuf_empty_rands[172]  = 1'b1;
    inbuf_empty_rands[173]  = 1'b0;
    inbuf_empty_rands[174]  = 1'b0;
    inbuf_empty_rands[175]  = 1'b1;
    inbuf_empty_rands[176]  = 1'b0;
    inbuf_empty_rands[177]  = 1'b1;
    inbuf_empty_rands[178]  = 1'b0;
    inbuf_empty_rands[179]  = 1'b1;
    inbuf_empty_rands[180]  = 1'b0;
    inbuf_empty_rands[181]  = 1'b1;
    inbuf_empty_rands[182]  = 1'b1;
    inbuf_empty_rands[183]  = 1'b1;
    inbuf_empty_rands[184]  = 1'b0;
    inbuf_empty_rands[185]  = 1'b1;
    inbuf_empty_rands[186]  = 1'b0;
    inbuf_empty_rands[187]  = 1'b1;
    inbuf_empty_rands[188]  = 1'b1;
    inbuf_empty_rands[189]  = 1'b1;
    inbuf_empty_rands[190]  = 1'b1;
    inbuf_empty_rands[191]  = 1'b0;
    inbuf_empty_rands[192]  = 1'b0;
    inbuf_empty_rands[193]  = 1'b1;
    inbuf_empty_rands[194]  = 1'b1;
    inbuf_empty_rands[195]  = 1'b0;
    inbuf_empty_rands[196]  = 1'b1;
    inbuf_empty_rands[197]  = 1'b0;
    inbuf_empty_rands[198]  = 1'b0;
    inbuf_empty_rands[199]  = 1'b0;
    inbuf_empty_rands[200]  = 1'b1;
    inbuf_empty_rands[201]  = 1'b0;
    inbuf_empty_rands[202]  = 1'b0;
    inbuf_empty_rands[203]  = 1'b1;
    inbuf_empty_rands[204]  = 1'b0;
    inbuf_empty_rands[205]  = 1'b1;
    inbuf_empty_rands[206]  = 1'b1;
    inbuf_empty_rands[207]  = 1'b1;
    inbuf_empty_rands[208]  = 1'b1;
    inbuf_empty_rands[209]  = 1'b0;
    inbuf_empty_rands[210]  = 1'b0;
    inbuf_empty_rands[211]  = 1'b0;
    inbuf_empty_rands[212]  = 1'b0;
    inbuf_empty_rands[213]  = 1'b1;
    inbuf_empty_rands[214]  = 1'b0;
    inbuf_empty_rands[215]  = 1'b0;
    inbuf_empty_rands[216]  = 1'b0;
    inbuf_empty_rands[217]  = 1'b1;
    inbuf_empty_rands[218]  = 1'b0;
    inbuf_empty_rands[219]  = 1'b0;
    inbuf_empty_rands[220]  = 1'b0;
    inbuf_empty_rands[221]  = 1'b1;
    inbuf_empty_rands[222]  = 1'b0;
    inbuf_empty_rands[223]  = 1'b0;
    inbuf_empty_rands[224]  = 1'b0;
    inbuf_empty_rands[225]  = 1'b1;
    inbuf_empty_rands[226]  = 1'b0;
    inbuf_empty_rands[227]  = 1'b1;
    inbuf_empty_rands[228]  = 1'b0;
    inbuf_empty_rands[229]  = 1'b1;
    inbuf_empty_rands[230]  = 1'b0;
    inbuf_empty_rands[231]  = 1'b1;
    inbuf_empty_rands[232]  = 1'b0;
    inbuf_empty_rands[233]  = 1'b1;
    inbuf_empty_rands[234]  = 1'b0;
    inbuf_empty_rands[235]  = 1'b1;
    inbuf_empty_rands[236]  = 1'b1;
    inbuf_empty_rands[237]  = 1'b0;
    inbuf_empty_rands[238]  = 1'b1;
    inbuf_empty_rands[239]  = 1'b0;
    inbuf_empty_rands[240]  = 1'b1;
    inbuf_empty_rands[241]  = 1'b0;
    inbuf_empty_rands[242]  = 1'b1;
    inbuf_empty_rands[243]  = 1'b0;
    inbuf_empty_rands[244]  = 1'b1;
    inbuf_empty_rands[245]  = 1'b0;
    inbuf_empty_rands[246]  = 1'b1;
    inbuf_empty_rands[247]  = 1'b0;
    inbuf_empty_rands[248]  = 1'b0;
    inbuf_empty_rands[249]  = 1'b1;
    inbuf_empty_rands[250]  = 1'b1;
    inbuf_empty_rands[251]  = 1'b0;
    inbuf_empty_rands[252]  = 1'b1;
    inbuf_empty_rands[253]  = 1'b1;
    inbuf_empty_rands[254]  = 1'b1;
    inbuf_empty_rands[255]  = 1'b0;
    inbuf_empty_rands[256]  = 1'b0;
    inbuf_empty_rands[257]  = 1'b1;
    inbuf_empty_rands[258]  = 1'b0;
    inbuf_empty_rands[259]  = 1'b1;
    inbuf_empty_rands[260]  = 1'b0;
    inbuf_empty_rands[261]  = 1'b1;
    inbuf_empty_rands[262]  = 1'b1;
    inbuf_empty_rands[263]  = 1'b1;
    inbuf_empty_rands[264]  = 1'b0;
    inbuf_empty_rands[265]  = 1'b0;
    inbuf_empty_rands[266]  = 1'b1;
    inbuf_empty_rands[267]  = 1'b0;
    inbuf_empty_rands[268]  = 1'b0;
    inbuf_empty_rands[269]  = 1'b0;
    inbuf_empty_rands[270]  = 1'b0;
    inbuf_empty_rands[271]  = 1'b1;
    inbuf_empty_rands[272]  = 1'b1;
    inbuf_empty_rands[273]  = 1'b0;
    inbuf_empty_rands[274]  = 1'b0;
    inbuf_empty_rands[275]  = 1'b1;
    inbuf_empty_rands[276]  = 1'b0;
    inbuf_empty_rands[277]  = 1'b0;
    inbuf_empty_rands[278]  = 1'b1;
    inbuf_empty_rands[279]  = 1'b1;
    inbuf_empty_rands[280]  = 1'b0;
    inbuf_empty_rands[281]  = 1'b0;
    inbuf_empty_rands[282]  = 1'b0;
    inbuf_empty_rands[283]  = 1'b1;
    inbuf_empty_rands[284]  = 1'b0;
    inbuf_empty_rands[285]  = 1'b0;
    inbuf_empty_rands[286]  = 1'b1;
    inbuf_empty_rands[287]  = 1'b0;
    inbuf_empty_rands[288]  = 1'b1;
    inbuf_empty_rands[289]  = 1'b1;
    inbuf_empty_rands[290]  = 1'b0;
    inbuf_empty_rands[291]  = 1'b0;
    inbuf_empty_rands[292]  = 1'b1;
    inbuf_empty_rands[293]  = 1'b1;
    inbuf_empty_rands[294]  = 1'b0;
    inbuf_empty_rands[295]  = 1'b1;
    inbuf_empty_rands[296]  = 1'b0;
    inbuf_empty_rands[297]  = 1'b1;
    inbuf_empty_rands[298]  = 1'b0;
    inbuf_empty_rands[299]  = 1'b0;
    inbuf_empty_rands[300]  = 1'b1;
    inbuf_empty_rands[301]  = 1'b1;
    inbuf_empty_rands[302]  = 1'b0;
    inbuf_empty_rands[303]  = 1'b0;
    inbuf_empty_rands[304]  = 1'b1;
    inbuf_empty_rands[305]  = 1'b0;
    inbuf_empty_rands[306]  = 1'b0;
    inbuf_empty_rands[307]  = 1'b1;
    inbuf_empty_rands[308]  = 1'b1;
    inbuf_empty_rands[309]  = 1'b1;
    inbuf_empty_rands[310]  = 1'b1;
    inbuf_empty_rands[311]  = 1'b1;
    inbuf_empty_rands[312]  = 1'b1;
    inbuf_empty_rands[313]  = 1'b0;
    inbuf_empty_rands[314]  = 1'b0;
    inbuf_empty_rands[315]  = 1'b0;
    inbuf_empty_rands[316]  = 1'b0;
    inbuf_empty_rands[317]  = 1'b1;
    inbuf_empty_rands[318]  = 1'b1;
    inbuf_empty_rands[319]  = 1'b1;
    inbuf_empty_rands[320]  = 1'b1;
    inbuf_empty_rands[321]  = 1'b0;
    inbuf_empty_rands[322]  = 1'b0;
    inbuf_empty_rands[323]  = 1'b1;
    inbuf_empty_rands[324]  = 1'b0;
    inbuf_empty_rands[325]  = 1'b0;
    inbuf_empty_rands[326]  = 1'b1;
    inbuf_empty_rands[327]  = 1'b0;
    inbuf_empty_rands[328]  = 1'b1;
    inbuf_empty_rands[329]  = 1'b0;
    inbuf_empty_rands[330]  = 1'b0;
    inbuf_empty_rands[331]  = 1'b1;
    inbuf_empty_rands[332]  = 1'b1;
    inbuf_empty_rands[333]  = 1'b0;
    inbuf_empty_rands[334]  = 1'b1;
    inbuf_empty_rands[335]  = 1'b0;
    inbuf_empty_rands[336]  = 1'b0;
    inbuf_empty_rands[337]  = 1'b1;
    inbuf_empty_rands[338]  = 1'b0;
    inbuf_empty_rands[339]  = 1'b0;
    inbuf_empty_rands[340]  = 1'b1;
    inbuf_empty_rands[341]  = 1'b1;
    inbuf_empty_rands[342]  = 1'b1;
    inbuf_empty_rands[343]  = 1'b0;
    inbuf_empty_rands[344]  = 1'b0;
    inbuf_empty_rands[345]  = 1'b0;
    inbuf_empty_rands[346]  = 1'b0;
    inbuf_empty_rands[347]  = 1'b1;
    inbuf_empty_rands[348]  = 1'b0;
    inbuf_empty_rands[349]  = 1'b1;
    inbuf_empty_rands[350]  = 1'b1;
    inbuf_empty_rands[351]  = 1'b0;
    inbuf_empty_rands[352]  = 1'b0;
    inbuf_empty_rands[353]  = 1'b1;
    inbuf_empty_rands[354]  = 1'b0;
    inbuf_empty_rands[355]  = 1'b1;
    inbuf_empty_rands[356]  = 1'b1;
    inbuf_empty_rands[357]  = 1'b1;
    inbuf_empty_rands[358]  = 1'b1;
    inbuf_empty_rands[359]  = 1'b0;
    inbuf_empty_rands[360]  = 1'b0;
    inbuf_empty_rands[361]  = 1'b0;
    inbuf_empty_rands[362]  = 1'b0;
    inbuf_empty_rands[363]  = 1'b0;
    inbuf_empty_rands[364]  = 1'b1;
    inbuf_empty_rands[365]  = 1'b1;
    inbuf_empty_rands[366]  = 1'b0;
    inbuf_empty_rands[367]  = 1'b0;
    inbuf_empty_rands[368]  = 1'b0;
    inbuf_empty_rands[369]  = 1'b0;
    inbuf_empty_rands[370]  = 1'b1;
    inbuf_empty_rands[371]  = 1'b0;
    inbuf_empty_rands[372]  = 1'b1;
    inbuf_empty_rands[373]  = 1'b0;
    inbuf_empty_rands[374]  = 1'b0;
    inbuf_empty_rands[375]  = 1'b0;
    inbuf_empty_rands[376]  = 1'b1;
    inbuf_empty_rands[377]  = 1'b0;
    inbuf_empty_rands[378]  = 1'b0;
    inbuf_empty_rands[379]  = 1'b1;
    inbuf_empty_rands[380]  = 1'b1;
    inbuf_empty_rands[381]  = 1'b0;
    inbuf_empty_rands[382]  = 1'b0;
    inbuf_empty_rands[383]  = 1'b1;
    inbuf_empty_rands[384]  = 1'b1;
    inbuf_empty_rands[385]  = 1'b0;
    inbuf_empty_rands[386]  = 1'b1;
    inbuf_empty_rands[387]  = 1'b1;
    inbuf_empty_rands[388]  = 1'b0;
    inbuf_empty_rands[389]  = 1'b0;
    inbuf_empty_rands[390]  = 1'b0;
    inbuf_empty_rands[391]  = 1'b0;
    inbuf_empty_rands[392]  = 1'b0;
    inbuf_empty_rands[393]  = 1'b1;
    inbuf_empty_rands[394]  = 1'b0;
    inbuf_empty_rands[395]  = 1'b0;
    inbuf_empty_rands[396]  = 1'b0;
    inbuf_empty_rands[397]  = 1'b0;
    inbuf_empty_rands[398]  = 1'b1;
    inbuf_empty_rands[399]  = 1'b1;
    inbuf_empty_rands[400]  = 1'b0;
    inbuf_empty_rands[401]  = 1'b0;
    inbuf_empty_rands[402]  = 1'b1;
    inbuf_empty_rands[403]  = 1'b0;
    inbuf_empty_rands[404]  = 1'b1;
    inbuf_empty_rands[405]  = 1'b1;
    inbuf_empty_rands[406]  = 1'b1;
    inbuf_empty_rands[407]  = 1'b1;
    inbuf_empty_rands[408]  = 1'b0;
    inbuf_empty_rands[409]  = 1'b0;
    inbuf_empty_rands[410]  = 1'b1;
    inbuf_empty_rands[411]  = 1'b0;
    inbuf_empty_rands[412]  = 1'b0;
    inbuf_empty_rands[413]  = 1'b1;
    inbuf_empty_rands[414]  = 1'b0;
    inbuf_empty_rands[415]  = 1'b1;
    inbuf_empty_rands[416]  = 1'b1;
    inbuf_empty_rands[417]  = 1'b1;
    inbuf_empty_rands[418]  = 1'b0;
    inbuf_empty_rands[419]  = 1'b0;
    inbuf_empty_rands[420]  = 1'b1;
    inbuf_empty_rands[421]  = 1'b0;
    inbuf_empty_rands[422]  = 1'b1;
    inbuf_empty_rands[423]  = 1'b1;
    inbuf_empty_rands[424]  = 1'b0;
    inbuf_empty_rands[425]  = 1'b1;
    inbuf_empty_rands[426]  = 1'b1;
    inbuf_empty_rands[427]  = 1'b0;
    inbuf_empty_rands[428]  = 1'b0;
    inbuf_empty_rands[429]  = 1'b1;
    inbuf_empty_rands[430]  = 1'b1;
    inbuf_empty_rands[431]  = 1'b1;
    inbuf_empty_rands[432]  = 1'b1;
    inbuf_empty_rands[433]  = 1'b1;
    inbuf_empty_rands[434]  = 1'b0;
    inbuf_empty_rands[435]  = 1'b0;
    inbuf_empty_rands[436]  = 1'b1;
    inbuf_empty_rands[437]  = 1'b1;
    inbuf_empty_rands[438]  = 1'b0;
    inbuf_empty_rands[439]  = 1'b1;
    inbuf_empty_rands[440]  = 1'b0;
    inbuf_empty_rands[441]  = 1'b0;
    inbuf_empty_rands[442]  = 1'b1;
    inbuf_empty_rands[443]  = 1'b1;
    inbuf_empty_rands[444]  = 1'b1;
    inbuf_empty_rands[445]  = 1'b1;
    inbuf_empty_rands[446]  = 1'b0;
    inbuf_empty_rands[447]  = 1'b0;
    inbuf_empty_rands[448]  = 1'b1;
    inbuf_empty_rands[449]  = 1'b0;
    inbuf_empty_rands[450]  = 1'b0;
    inbuf_empty_rands[451]  = 1'b0;
    inbuf_empty_rands[452]  = 1'b1;
    inbuf_empty_rands[453]  = 1'b1;
    inbuf_empty_rands[454]  = 1'b0;
    inbuf_empty_rands[455]  = 1'b1;
    inbuf_empty_rands[456]  = 1'b1;
    inbuf_empty_rands[457]  = 1'b0;
    inbuf_empty_rands[458]  = 1'b1;
    inbuf_empty_rands[459]  = 1'b0;
    inbuf_empty_rands[460]  = 1'b1;
    inbuf_empty_rands[461]  = 1'b0;
    inbuf_empty_rands[462]  = 1'b1;
    inbuf_empty_rands[463]  = 1'b0;
    inbuf_empty_rands[464]  = 1'b1;
    inbuf_empty_rands[465]  = 1'b1;
    inbuf_empty_rands[466]  = 1'b0;
    inbuf_empty_rands[467]  = 1'b0;
    inbuf_empty_rands[468]  = 1'b1;
    inbuf_empty_rands[469]  = 1'b0;
    inbuf_empty_rands[470]  = 1'b1;
    inbuf_empty_rands[471]  = 1'b1;
    inbuf_empty_rands[472]  = 1'b0;
    inbuf_empty_rands[473]  = 1'b1;
    inbuf_empty_rands[474]  = 1'b1;
    inbuf_empty_rands[475]  = 1'b0;
    inbuf_empty_rands[476]  = 1'b1;
    inbuf_empty_rands[477]  = 1'b1;
    inbuf_empty_rands[478]  = 1'b0;
    inbuf_empty_rands[479]  = 1'b1;
    inbuf_empty_rands[480]  = 1'b1;
    inbuf_empty_rands[481]  = 1'b0;
    inbuf_empty_rands[482]  = 1'b0;
    inbuf_empty_rands[483]  = 1'b1;
    inbuf_empty_rands[484]  = 1'b1;
    inbuf_empty_rands[485]  = 1'b0;
    inbuf_empty_rands[486]  = 1'b1;
    inbuf_empty_rands[487]  = 1'b0;
    inbuf_empty_rands[488]  = 1'b1;
    inbuf_empty_rands[489]  = 1'b1;
    inbuf_empty_rands[490]  = 1'b0;
    inbuf_empty_rands[491]  = 1'b1;
    inbuf_empty_rands[492]  = 1'b0;
    inbuf_empty_rands[493]  = 1'b1;
    inbuf_empty_rands[494]  = 1'b1;
    inbuf_empty_rands[495]  = 1'b0;
    inbuf_empty_rands[496]  = 1'b1;
    inbuf_empty_rands[497]  = 1'b0;
    inbuf_empty_rands[498]  = 1'b1;
    inbuf_empty_rands[499]  = 1'b1;
    inbuf_empty_rands[500]  = 1'b1;
    inbuf_empty_rands[501]  = 1'b1;
    inbuf_empty_rands[502]  = 1'b1;
    inbuf_empty_rands[503]  = 1'b0;
    inbuf_empty_rands[504]  = 1'b0;
    inbuf_empty_rands[505]  = 1'b0;
    inbuf_empty_rands[506]  = 1'b0;
    inbuf_empty_rands[507]  = 1'b1;
    inbuf_empty_rands[508]  = 1'b1;
    inbuf_empty_rands[509]  = 1'b1;
    inbuf_empty_rands[510]  = 1'b0;
    inbuf_empty_rands[511]  = 1'b1;
    inbuf_empty_rands[512]  = 1'b0;
    inbuf_empty_rands[513]  = 1'b0;
    inbuf_empty_rands[514]  = 1'b0;
    inbuf_empty_rands[515]  = 1'b1;
    inbuf_empty_rands[516]  = 1'b1;
    inbuf_empty_rands[517]  = 1'b1;
    inbuf_empty_rands[518]  = 1'b1;
    inbuf_empty_rands[519]  = 1'b1;
    inbuf_empty_rands[520]  = 1'b1;
    inbuf_empty_rands[521]  = 1'b1;
    inbuf_empty_rands[522]  = 1'b1;
    inbuf_empty_rands[523]  = 1'b1;
    inbuf_empty_rands[524]  = 1'b0;
    inbuf_empty_rands[525]  = 1'b1;
    inbuf_empty_rands[526]  = 1'b0;
    inbuf_empty_rands[527]  = 1'b1;
    inbuf_empty_rands[528]  = 1'b1;
    inbuf_empty_rands[529]  = 1'b1;
    inbuf_empty_rands[530]  = 1'b1;
    inbuf_empty_rands[531]  = 1'b0;
    inbuf_empty_rands[532]  = 1'b1;
    inbuf_empty_rands[533]  = 1'b0;
    inbuf_empty_rands[534]  = 1'b1;
    inbuf_empty_rands[535]  = 1'b1;
    inbuf_empty_rands[536]  = 1'b0;
    inbuf_empty_rands[537]  = 1'b1;
    inbuf_empty_rands[538]  = 1'b0;
    inbuf_empty_rands[539]  = 1'b1;
    inbuf_empty_rands[540]  = 1'b0;
    inbuf_empty_rands[541]  = 1'b1;
    inbuf_empty_rands[542]  = 1'b1;
    inbuf_empty_rands[543]  = 1'b0;
    inbuf_empty_rands[544]  = 1'b1;
    inbuf_empty_rands[545]  = 1'b1;
    inbuf_empty_rands[546]  = 1'b0;
    inbuf_empty_rands[547]  = 1'b0;
    inbuf_empty_rands[548]  = 1'b1;
    inbuf_empty_rands[549]  = 1'b1;
    inbuf_empty_rands[550]  = 1'b1;
    inbuf_empty_rands[551]  = 1'b0;
    inbuf_empty_rands[552]  = 1'b1;
    inbuf_empty_rands[553]  = 1'b1;
    inbuf_empty_rands[554]  = 1'b0;
    inbuf_empty_rands[555]  = 1'b1;
    inbuf_empty_rands[556]  = 1'b1;
    inbuf_empty_rands[557]  = 1'b0;
    inbuf_empty_rands[558]  = 1'b1;
    inbuf_empty_rands[559]  = 1'b1;
    inbuf_empty_rands[560]  = 1'b0;
    inbuf_empty_rands[561]  = 1'b1;
    inbuf_empty_rands[562]  = 1'b0;
    inbuf_empty_rands[563]  = 1'b1;
    inbuf_empty_rands[564]  = 1'b0;
    inbuf_empty_rands[565]  = 1'b0;
    inbuf_empty_rands[566]  = 1'b1;
    inbuf_empty_rands[567]  = 1'b1;
    inbuf_empty_rands[568]  = 1'b1;
    inbuf_empty_rands[569]  = 1'b0;
    inbuf_empty_rands[570]  = 1'b0;
    inbuf_empty_rands[571]  = 1'b0;
    inbuf_empty_rands[572]  = 1'b0;
    inbuf_empty_rands[573]  = 1'b1;
    inbuf_empty_rands[574]  = 1'b1;
    inbuf_empty_rands[575]  = 1'b0;
    inbuf_empty_rands[576]  = 1'b0;
    inbuf_empty_rands[577]  = 1'b0;
    inbuf_empty_rands[578]  = 1'b1;
    inbuf_empty_rands[579]  = 1'b0;
    inbuf_empty_rands[580]  = 1'b0;
    inbuf_empty_rands[581]  = 1'b0;
    inbuf_empty_rands[582]  = 1'b0;
    inbuf_empty_rands[583]  = 1'b0;
    inbuf_empty_rands[584]  = 1'b1;
    inbuf_empty_rands[585]  = 1'b1;
    inbuf_empty_rands[586]  = 1'b0;
    inbuf_empty_rands[587]  = 1'b0;
    inbuf_empty_rands[588]  = 1'b0;
    inbuf_empty_rands[589]  = 1'b0;
    inbuf_empty_rands[590]  = 1'b1;
    inbuf_empty_rands[591]  = 1'b1;
    inbuf_empty_rands[592]  = 1'b0;
    inbuf_empty_rands[593]  = 1'b0;
    inbuf_empty_rands[594]  = 1'b0;
    inbuf_empty_rands[595]  = 1'b1;
    inbuf_empty_rands[596]  = 1'b1;
    inbuf_empty_rands[597]  = 1'b0;
    inbuf_empty_rands[598]  = 1'b1;
    inbuf_empty_rands[599]  = 1'b0;
    inbuf_empty_rands[600]  = 1'b0;
    inbuf_empty_rands[601]  = 1'b0;
    inbuf_empty_rands[602]  = 1'b1;
    inbuf_empty_rands[603]  = 1'b1;
    inbuf_empty_rands[604]  = 1'b1;
    inbuf_empty_rands[605]  = 1'b1;
    inbuf_empty_rands[606]  = 1'b1;
    inbuf_empty_rands[607]  = 1'b0;
    inbuf_empty_rands[608]  = 1'b0;
    inbuf_empty_rands[609]  = 1'b0;
    inbuf_empty_rands[610]  = 1'b0;
    inbuf_empty_rands[611]  = 1'b0;
    inbuf_empty_rands[612]  = 1'b1;
    inbuf_empty_rands[613]  = 1'b0;
    inbuf_empty_rands[614]  = 1'b1;
    inbuf_empty_rands[615]  = 1'b1;
    inbuf_empty_rands[616]  = 1'b1;
    inbuf_empty_rands[617]  = 1'b1;
    inbuf_empty_rands[618]  = 1'b1;
    inbuf_empty_rands[619]  = 1'b1;
    inbuf_empty_rands[620]  = 1'b0;
    inbuf_empty_rands[621]  = 1'b0;
    inbuf_empty_rands[622]  = 1'b1;
    inbuf_empty_rands[623]  = 1'b0;
    inbuf_empty_rands[624]  = 1'b0;
    inbuf_empty_rands[625]  = 1'b1;
    inbuf_empty_rands[626]  = 1'b0;
    inbuf_empty_rands[627]  = 1'b1;
    inbuf_empty_rands[628]  = 1'b0;
    inbuf_empty_rands[629]  = 1'b1;
    inbuf_empty_rands[630]  = 1'b1;
    inbuf_empty_rands[631]  = 1'b0;
    inbuf_empty_rands[632]  = 1'b0;
    inbuf_empty_rands[633]  = 1'b1;
    inbuf_empty_rands[634]  = 1'b1;
    inbuf_empty_rands[635]  = 1'b1;
    inbuf_empty_rands[636]  = 1'b1;
    inbuf_empty_rands[637]  = 1'b0;
    inbuf_empty_rands[638]  = 1'b1;
    inbuf_empty_rands[639]  = 1'b0;
    inbuf_empty_rands[640]  = 1'b1;
    inbuf_empty_rands[641]  = 1'b0;
    inbuf_empty_rands[642]  = 1'b1;
    inbuf_empty_rands[643]  = 1'b0;
    inbuf_empty_rands[644]  = 1'b0;
    inbuf_empty_rands[645]  = 1'b0;
    inbuf_empty_rands[646]  = 1'b0;
    inbuf_empty_rands[647]  = 1'b1;
    inbuf_empty_rands[648]  = 1'b1;
    inbuf_empty_rands[649]  = 1'b0;
    inbuf_empty_rands[650]  = 1'b1;
    inbuf_empty_rands[651]  = 1'b0;
    inbuf_empty_rands[652]  = 1'b1;
    inbuf_empty_rands[653]  = 1'b1;
    inbuf_empty_rands[654]  = 1'b1;
    inbuf_empty_rands[655]  = 1'b1;
    inbuf_empty_rands[656]  = 1'b0;
    inbuf_empty_rands[657]  = 1'b0;
    inbuf_empty_rands[658]  = 1'b0;
    inbuf_empty_rands[659]  = 1'b1;
    inbuf_empty_rands[660]  = 1'b1;
    inbuf_empty_rands[661]  = 1'b1;
    inbuf_empty_rands[662]  = 1'b1;
    inbuf_empty_rands[663]  = 1'b0;
    inbuf_empty_rands[664]  = 1'b0;
    inbuf_empty_rands[665]  = 1'b1;
    inbuf_empty_rands[666]  = 1'b1;
    inbuf_empty_rands[667]  = 1'b0;
    inbuf_empty_rands[668]  = 1'b1;
    inbuf_empty_rands[669]  = 1'b0;
    inbuf_empty_rands[670]  = 1'b1;
    inbuf_empty_rands[671]  = 1'b0;
    inbuf_empty_rands[672]  = 1'b0;
    inbuf_empty_rands[673]  = 1'b1;
    inbuf_empty_rands[674]  = 1'b0;
    inbuf_empty_rands[675]  = 1'b0;
    inbuf_empty_rands[676]  = 1'b1;
    inbuf_empty_rands[677]  = 1'b0;
    inbuf_empty_rands[678]  = 1'b1;
    inbuf_empty_rands[679]  = 1'b1;
    inbuf_empty_rands[680]  = 1'b0;
    inbuf_empty_rands[681]  = 1'b1;
    inbuf_empty_rands[682]  = 1'b0;
    inbuf_empty_rands[683]  = 1'b1;
    inbuf_empty_rands[684]  = 1'b1;
    inbuf_empty_rands[685]  = 1'b1;
    inbuf_empty_rands[686]  = 1'b1;
    inbuf_empty_rands[687]  = 1'b1;
    inbuf_empty_rands[688]  = 1'b1;
    inbuf_empty_rands[689]  = 1'b1;
    inbuf_empty_rands[690]  = 1'b0;
    inbuf_empty_rands[691]  = 1'b0;
    inbuf_empty_rands[692]  = 1'b1;
    inbuf_empty_rands[693]  = 1'b0;
    inbuf_empty_rands[694]  = 1'b1;
    inbuf_empty_rands[695]  = 1'b0;
    inbuf_empty_rands[696]  = 1'b1;
    inbuf_empty_rands[697]  = 1'b1;
    inbuf_empty_rands[698]  = 1'b0;
    inbuf_empty_rands[699]  = 1'b1;
    inbuf_empty_rands[700]  = 1'b1;
    inbuf_empty_rands[701]  = 1'b1;
    inbuf_empty_rands[702]  = 1'b0;
    inbuf_empty_rands[703]  = 1'b0;
    inbuf_empty_rands[704]  = 1'b1;
    inbuf_empty_rands[705]  = 1'b1;
    inbuf_empty_rands[706]  = 1'b1;
    inbuf_empty_rands[707]  = 1'b1;
    inbuf_empty_rands[708]  = 1'b1;
    inbuf_empty_rands[709]  = 1'b0;
    inbuf_empty_rands[710]  = 1'b1;
    inbuf_empty_rands[711]  = 1'b0;
    inbuf_empty_rands[712]  = 1'b1;
    inbuf_empty_rands[713]  = 1'b0;
    inbuf_empty_rands[714]  = 1'b0;
    inbuf_empty_rands[715]  = 1'b1;
    inbuf_empty_rands[716]  = 1'b1;
    inbuf_empty_rands[717]  = 1'b1;
    inbuf_empty_rands[718]  = 1'b1;
    inbuf_empty_rands[719]  = 1'b0;
    inbuf_empty_rands[720]  = 1'b0;
    inbuf_empty_rands[721]  = 1'b0;
    inbuf_empty_rands[722]  = 1'b1;
    inbuf_empty_rands[723]  = 1'b0;
    inbuf_empty_rands[724]  = 1'b0;
    inbuf_empty_rands[725]  = 1'b1;
    inbuf_empty_rands[726]  = 1'b1;
    inbuf_empty_rands[727]  = 1'b0;
    inbuf_empty_rands[728]  = 1'b1;
    inbuf_empty_rands[729]  = 1'b1;
    inbuf_empty_rands[730]  = 1'b0;
    inbuf_empty_rands[731]  = 1'b0;
    inbuf_empty_rands[732]  = 1'b0;
    inbuf_empty_rands[733]  = 1'b1;
    inbuf_empty_rands[734]  = 1'b1;
    inbuf_empty_rands[735]  = 1'b1;
    inbuf_empty_rands[736]  = 1'b0;
    inbuf_empty_rands[737]  = 1'b1;
    inbuf_empty_rands[738]  = 1'b0;
    inbuf_empty_rands[739]  = 1'b0;
    inbuf_empty_rands[740]  = 1'b0;
    inbuf_empty_rands[741]  = 1'b1;
    inbuf_empty_rands[742]  = 1'b0;
    inbuf_empty_rands[743]  = 1'b0;
    inbuf_empty_rands[744]  = 1'b0;
    inbuf_empty_rands[745]  = 1'b0;
    inbuf_empty_rands[746]  = 1'b1;
    inbuf_empty_rands[747]  = 1'b1;
    inbuf_empty_rands[748]  = 1'b1;
    inbuf_empty_rands[749]  = 1'b0;
    inbuf_empty_rands[750]  = 1'b1;
    inbuf_empty_rands[751]  = 1'b0;
    inbuf_empty_rands[752]  = 1'b0;
    inbuf_empty_rands[753]  = 1'b1;
    inbuf_empty_rands[754]  = 1'b0;
    inbuf_empty_rands[755]  = 1'b0;
    inbuf_empty_rands[756]  = 1'b1;
    inbuf_empty_rands[757]  = 1'b1;
    inbuf_empty_rands[758]  = 1'b0;
    inbuf_empty_rands[759]  = 1'b0;
    inbuf_empty_rands[760]  = 1'b1;
    inbuf_empty_rands[761]  = 1'b1;
    inbuf_empty_rands[762]  = 1'b0;
    inbuf_empty_rands[763]  = 1'b0;
    inbuf_empty_rands[764]  = 1'b1;
    inbuf_empty_rands[765]  = 1'b0;
    inbuf_empty_rands[766]  = 1'b1;
    inbuf_empty_rands[767]  = 1'b1;
    inbuf_empty_rands[768]  = 1'b1;
    inbuf_empty_rands[769]  = 1'b0;
    inbuf_empty_rands[770]  = 1'b0;
    inbuf_empty_rands[771]  = 1'b1;
    inbuf_empty_rands[772]  = 1'b0;
    inbuf_empty_rands[773]  = 1'b1;
    inbuf_empty_rands[774]  = 1'b1;
    inbuf_empty_rands[775]  = 1'b1;
    inbuf_empty_rands[776]  = 1'b0;
    inbuf_empty_rands[777]  = 1'b1;
    inbuf_empty_rands[778]  = 1'b1;
    inbuf_empty_rands[779]  = 1'b0;
    inbuf_empty_rands[780]  = 1'b0;
    inbuf_empty_rands[781]  = 1'b1;
    inbuf_empty_rands[782]  = 1'b1;
    inbuf_empty_rands[783]  = 1'b1;
    inbuf_empty_rands[784]  = 1'b0;
    inbuf_empty_rands[785]  = 1'b1;
    inbuf_empty_rands[786]  = 1'b1;
    inbuf_empty_rands[787]  = 1'b0;
    inbuf_empty_rands[788]  = 1'b0;
    inbuf_empty_rands[789]  = 1'b0;
    inbuf_empty_rands[790]  = 1'b0;
    inbuf_empty_rands[791]  = 1'b1;
    inbuf_empty_rands[792]  = 1'b0;
    inbuf_empty_rands[793]  = 1'b1;
    inbuf_empty_rands[794]  = 1'b0;
    inbuf_empty_rands[795]  = 1'b0;
    inbuf_empty_rands[796]  = 1'b1;
    inbuf_empty_rands[797]  = 1'b1;
    inbuf_empty_rands[798]  = 1'b1;
    inbuf_empty_rands[799]  = 1'b0;
    inbuf_empty_rands[800]  = 1'b0;
    inbuf_empty_rands[801]  = 1'b1;
    inbuf_empty_rands[802]  = 1'b0;
    inbuf_empty_rands[803]  = 1'b1;
    inbuf_empty_rands[804]  = 1'b1;
    inbuf_empty_rands[805]  = 1'b0;
    inbuf_empty_rands[806]  = 1'b0;
    inbuf_empty_rands[807]  = 1'b0;
    inbuf_empty_rands[808]  = 1'b0;
    inbuf_empty_rands[809]  = 1'b1;
    inbuf_empty_rands[810]  = 1'b1;
    inbuf_empty_rands[811]  = 1'b1;
    inbuf_empty_rands[812]  = 1'b0;
    inbuf_empty_rands[813]  = 1'b1;
    inbuf_empty_rands[814]  = 1'b0;
    inbuf_empty_rands[815]  = 1'b1;
    inbuf_empty_rands[816]  = 1'b1;
    inbuf_empty_rands[817]  = 1'b1;
    inbuf_empty_rands[818]  = 1'b0;
    inbuf_empty_rands[819]  = 1'b1;
    inbuf_empty_rands[820]  = 1'b0;
    inbuf_empty_rands[821]  = 1'b1;
    inbuf_empty_rands[822]  = 1'b0;
    inbuf_empty_rands[823]  = 1'b1;
    inbuf_empty_rands[824]  = 1'b0;
    inbuf_empty_rands[825]  = 1'b1;
    inbuf_empty_rands[826]  = 1'b1;
    inbuf_empty_rands[827]  = 1'b1;
    inbuf_empty_rands[828]  = 1'b1;
    inbuf_empty_rands[829]  = 1'b1;
    inbuf_empty_rands[830]  = 1'b1;
    inbuf_empty_rands[831]  = 1'b1;
    inbuf_empty_rands[832]  = 1'b0;
    inbuf_empty_rands[833]  = 1'b1;
    inbuf_empty_rands[834]  = 1'b0;
    inbuf_empty_rands[835]  = 1'b1;
    inbuf_empty_rands[836]  = 1'b1;
    inbuf_empty_rands[837]  = 1'b0;
    inbuf_empty_rands[838]  = 1'b1;
    inbuf_empty_rands[839]  = 1'b1;
    inbuf_empty_rands[840]  = 1'b0;
    inbuf_empty_rands[841]  = 1'b0;
    inbuf_empty_rands[842]  = 1'b0;
    inbuf_empty_rands[843]  = 1'b0;
    inbuf_empty_rands[844]  = 1'b1;
    inbuf_empty_rands[845]  = 1'b0;
    inbuf_empty_rands[846]  = 1'b0;
    inbuf_empty_rands[847]  = 1'b0;
    inbuf_empty_rands[848]  = 1'b0;
    inbuf_empty_rands[849]  = 1'b1;
    inbuf_empty_rands[850]  = 1'b1;
    inbuf_empty_rands[851]  = 1'b1;
    inbuf_empty_rands[852]  = 1'b0;
    inbuf_empty_rands[853]  = 1'b1;
    inbuf_empty_rands[854]  = 1'b1;
    inbuf_empty_rands[855]  = 1'b0;
    inbuf_empty_rands[856]  = 1'b1;
    inbuf_empty_rands[857]  = 1'b0;
    inbuf_empty_rands[858]  = 1'b1;
    inbuf_empty_rands[859]  = 1'b1;
    inbuf_empty_rands[860]  = 1'b1;
    inbuf_empty_rands[861]  = 1'b1;
    inbuf_empty_rands[862]  = 1'b1;
    inbuf_empty_rands[863]  = 1'b0;
    inbuf_empty_rands[864]  = 1'b1;
    inbuf_empty_rands[865]  = 1'b1;
    inbuf_empty_rands[866]  = 1'b0;
    inbuf_empty_rands[867]  = 1'b0;
    inbuf_empty_rands[868]  = 1'b0;
    inbuf_empty_rands[869]  = 1'b1;
    inbuf_empty_rands[870]  = 1'b1;
    inbuf_empty_rands[871]  = 1'b0;
    inbuf_empty_rands[872]  = 1'b1;
    inbuf_empty_rands[873]  = 1'b0;
    inbuf_empty_rands[874]  = 1'b1;
    inbuf_empty_rands[875]  = 1'b1;
    inbuf_empty_rands[876]  = 1'b1;
    inbuf_empty_rands[877]  = 1'b1;
    inbuf_empty_rands[878]  = 1'b0;
    inbuf_empty_rands[879]  = 1'b1;
    inbuf_empty_rands[880]  = 1'b0;
    inbuf_empty_rands[881]  = 1'b0;
    inbuf_empty_rands[882]  = 1'b1;
    inbuf_empty_rands[883]  = 1'b0;
    inbuf_empty_rands[884]  = 1'b0;
    inbuf_empty_rands[885]  = 1'b1;
    inbuf_empty_rands[886]  = 1'b1;
    inbuf_empty_rands[887]  = 1'b0;
    inbuf_empty_rands[888]  = 1'b0;
    inbuf_empty_rands[889]  = 1'b1;
    inbuf_empty_rands[890]  = 1'b0;
    inbuf_empty_rands[891]  = 1'b0;
    inbuf_empty_rands[892]  = 1'b0;
    inbuf_empty_rands[893]  = 1'b0;
    inbuf_empty_rands[894]  = 1'b1;
    inbuf_empty_rands[895]  = 1'b1;
    inbuf_empty_rands[896]  = 1'b1;
    inbuf_empty_rands[897]  = 1'b0;
    inbuf_empty_rands[898]  = 1'b1;
    inbuf_empty_rands[899]  = 1'b1;
    inbuf_empty_rands[900]  = 1'b1;
    inbuf_empty_rands[901]  = 1'b1;
    inbuf_empty_rands[902]  = 1'b1;
    inbuf_empty_rands[903]  = 1'b0;
    inbuf_empty_rands[904]  = 1'b0;
    inbuf_empty_rands[905]  = 1'b0;
    inbuf_empty_rands[906]  = 1'b0;
    inbuf_empty_rands[907]  = 1'b0;
    inbuf_empty_rands[908]  = 1'b1;
    inbuf_empty_rands[909]  = 1'b0;
    inbuf_empty_rands[910]  = 1'b1;
    inbuf_empty_rands[911]  = 1'b0;
    inbuf_empty_rands[912]  = 1'b1;
    inbuf_empty_rands[913]  = 1'b1;
    inbuf_empty_rands[914]  = 1'b0;
    inbuf_empty_rands[915]  = 1'b1;
    inbuf_empty_rands[916]  = 1'b1;
    inbuf_empty_rands[917]  = 1'b0;
    inbuf_empty_rands[918]  = 1'b0;
    inbuf_empty_rands[919]  = 1'b1;
    inbuf_empty_rands[920]  = 1'b0;
    inbuf_empty_rands[921]  = 1'b0;
    inbuf_empty_rands[922]  = 1'b1;
    inbuf_empty_rands[923]  = 1'b1;
    inbuf_empty_rands[924]  = 1'b1;
    inbuf_empty_rands[925]  = 1'b1;
    inbuf_empty_rands[926]  = 1'b0;
    inbuf_empty_rands[927]  = 1'b0;
    inbuf_empty_rands[928]  = 1'b1;
    inbuf_empty_rands[929]  = 1'b0;
    inbuf_empty_rands[930]  = 1'b1;
    inbuf_empty_rands[931]  = 1'b1;
    inbuf_empty_rands[932]  = 1'b1;
    inbuf_empty_rands[933]  = 1'b0;
    inbuf_empty_rands[934]  = 1'b0;
    inbuf_empty_rands[935]  = 1'b1;
    inbuf_empty_rands[936]  = 1'b1;
    inbuf_empty_rands[937]  = 1'b1;
    inbuf_empty_rands[938]  = 1'b1;
    inbuf_empty_rands[939]  = 1'b0;
    inbuf_empty_rands[940]  = 1'b1;
    inbuf_empty_rands[941]  = 1'b1;
    inbuf_empty_rands[942]  = 1'b1;
    inbuf_empty_rands[943]  = 1'b1;
    inbuf_empty_rands[944]  = 1'b0;
    inbuf_empty_rands[945]  = 1'b0;
    inbuf_empty_rands[946]  = 1'b1;
    inbuf_empty_rands[947]  = 1'b0;
    inbuf_empty_rands[948]  = 1'b0;
    inbuf_empty_rands[949]  = 1'b0;
    inbuf_empty_rands[950]  = 1'b0;
    inbuf_empty_rands[951]  = 1'b0;
    inbuf_empty_rands[952]  = 1'b1;
    inbuf_empty_rands[953]  = 1'b0;
    inbuf_empty_rands[954]  = 1'b1;
    inbuf_empty_rands[955]  = 1'b1;
    inbuf_empty_rands[956]  = 1'b1;
    inbuf_empty_rands[957]  = 1'b1;
    inbuf_empty_rands[958]  = 1'b0;
    inbuf_empty_rands[959]  = 1'b1;
    inbuf_empty_rands[960]  = 1'b0;
    inbuf_empty_rands[961]  = 1'b0;
    inbuf_empty_rands[962]  = 1'b0;
    inbuf_empty_rands[963]  = 1'b1;
    inbuf_empty_rands[964]  = 1'b1;
    inbuf_empty_rands[965]  = 1'b1;
    inbuf_empty_rands[966]  = 1'b0;
    inbuf_empty_rands[967]  = 1'b0;
    inbuf_empty_rands[968]  = 1'b0;
    inbuf_empty_rands[969]  = 1'b1;
    inbuf_empty_rands[970]  = 1'b0;
    inbuf_empty_rands[971]  = 1'b0;
    inbuf_empty_rands[972]  = 1'b1;
    inbuf_empty_rands[973]  = 1'b1;
    inbuf_empty_rands[974]  = 1'b0;
    inbuf_empty_rands[975]  = 1'b0;
    inbuf_empty_rands[976]  = 1'b0;
    inbuf_empty_rands[977]  = 1'b1;
    inbuf_empty_rands[978]  = 1'b1;
    inbuf_empty_rands[979]  = 1'b1;
    inbuf_empty_rands[980]  = 1'b0;
    inbuf_empty_rands[981]  = 1'b1;
    inbuf_empty_rands[982]  = 1'b0;
    inbuf_empty_rands[983]  = 1'b0;
    inbuf_empty_rands[984]  = 1'b1;
    inbuf_empty_rands[985]  = 1'b0;
    inbuf_empty_rands[986]  = 1'b0;
    inbuf_empty_rands[987]  = 1'b1;
    inbuf_empty_rands[988]  = 1'b0;
    inbuf_empty_rands[989]  = 1'b1;
    inbuf_empty_rands[990]  = 1'b0;
    inbuf_empty_rands[991]  = 1'b1;
    inbuf_empty_rands[992]  = 1'b0;
    inbuf_empty_rands[993]  = 1'b1;
    inbuf_empty_rands[994]  = 1'b0;
    inbuf_empty_rands[995]  = 1'b0;
    inbuf_empty_rands[996]  = 1'b0;
    inbuf_empty_rands[997]  = 1'b0;
    inbuf_empty_rands[998]  = 1'b0;
    inbuf_empty_rands[999]  = 1'b1;
    //inbuf_empty_rands[1000] = 1'b1;

    buffer_full_rands[0]    = 1'b1;
    buffer_full_rands[1]    = 1'b1;
    buffer_full_rands[2]    = 1'b1;
    buffer_full_rands[3]    = 1'b1;
    buffer_full_rands[4]    = 1'b1;
    buffer_full_rands[5]    = 1'b1;
    buffer_full_rands[6]    = 1'b0;
    buffer_full_rands[7]    = 1'b0;
    buffer_full_rands[8]    = 1'b1;
    buffer_full_rands[9]    = 1'b1;
    buffer_full_rands[10]   = 1'b1;
    buffer_full_rands[11]   = 1'b0;
    buffer_full_rands[12]   = 1'b0;
    buffer_full_rands[13]   = 1'b0;
    buffer_full_rands[14]   = 1'b0;
    buffer_full_rands[15]   = 1'b0;
    buffer_full_rands[16]   = 1'b1;
    buffer_full_rands[17]   = 1'b0;
    buffer_full_rands[18]   = 1'b0;
    buffer_full_rands[19]   = 1'b1;
    buffer_full_rands[20]   = 1'b0;
    buffer_full_rands[21]   = 1'b0;
    buffer_full_rands[22]   = 1'b1;
    buffer_full_rands[23]   = 1'b1;
    buffer_full_rands[24]   = 1'b1;
    buffer_full_rands[25]   = 1'b0;
    buffer_full_rands[26]   = 1'b0;
    buffer_full_rands[27]   = 1'b0;
    buffer_full_rands[28]   = 1'b1;
    buffer_full_rands[29]   = 1'b0;
    buffer_full_rands[30]   = 1'b0;
    buffer_full_rands[31]   = 1'b0;
    buffer_full_rands[32]   = 1'b1;
    buffer_full_rands[33]   = 1'b1;
    buffer_full_rands[34]   = 1'b1;
    buffer_full_rands[35]   = 1'b1;
    buffer_full_rands[36]   = 1'b1;
    buffer_full_rands[37]   = 1'b1;
    buffer_full_rands[38]   = 1'b0;
    buffer_full_rands[39]   = 1'b0;
    buffer_full_rands[40]   = 1'b0;
    buffer_full_rands[41]   = 1'b1;
    buffer_full_rands[42]   = 1'b0;
    buffer_full_rands[43]   = 1'b1;
    buffer_full_rands[44]   = 1'b0;
    buffer_full_rands[45]   = 1'b1;
    buffer_full_rands[46]   = 1'b0;
    buffer_full_rands[47]   = 1'b0;
    buffer_full_rands[48]   = 1'b0;
    buffer_full_rands[49]   = 1'b0;
    buffer_full_rands[50]   = 1'b1;
    buffer_full_rands[51]   = 1'b0;
    buffer_full_rands[52]   = 1'b1;
    buffer_full_rands[53]   = 1'b0;
    buffer_full_rands[54]   = 1'b1;
    buffer_full_rands[55]   = 1'b1;
    buffer_full_rands[56]   = 1'b1;
    buffer_full_rands[57]   = 1'b0;
    buffer_full_rands[58]   = 1'b0;
    buffer_full_rands[59]   = 1'b0;
    buffer_full_rands[60]   = 1'b1;
    buffer_full_rands[61]   = 1'b1;
    buffer_full_rands[62]   = 1'b1;
    buffer_full_rands[63]   = 1'b1;
    buffer_full_rands[64]   = 1'b1;
    buffer_full_rands[65]   = 1'b0;
    buffer_full_rands[66]   = 1'b1;
    buffer_full_rands[67]   = 1'b0;
    buffer_full_rands[68]   = 1'b0;
    buffer_full_rands[69]   = 1'b0;
    buffer_full_rands[70]   = 1'b1;
    buffer_full_rands[71]   = 1'b1;
    buffer_full_rands[72]   = 1'b1;
    buffer_full_rands[73]   = 1'b1;
    buffer_full_rands[74]   = 1'b0;
    buffer_full_rands[75]   = 1'b0;
    buffer_full_rands[76]   = 1'b0;
    buffer_full_rands[77]   = 1'b0;
    buffer_full_rands[78]   = 1'b1;
    buffer_full_rands[79]   = 1'b0;
    buffer_full_rands[80]   = 1'b0;
    buffer_full_rands[81]   = 1'b0;
    buffer_full_rands[82]   = 1'b0;
    buffer_full_rands[83]   = 1'b1;
    buffer_full_rands[84]   = 1'b0;
    buffer_full_rands[85]   = 1'b0;
    buffer_full_rands[86]   = 1'b0;
    buffer_full_rands[87]   = 1'b1;
    buffer_full_rands[88]   = 1'b0;
    buffer_full_rands[89]   = 1'b0;
    buffer_full_rands[90]   = 1'b0;
    buffer_full_rands[91]   = 1'b0;
    buffer_full_rands[92]   = 1'b1;
    buffer_full_rands[93]   = 1'b1;
    buffer_full_rands[94]   = 1'b1;
    buffer_full_rands[95]   = 1'b1;
    buffer_full_rands[96]   = 1'b1;
    buffer_full_rands[97]   = 1'b0;
    buffer_full_rands[98]   = 1'b1;
    buffer_full_rands[99]   = 1'b1;
    buffer_full_rands[100]  = 1'b0;
    buffer_full_rands[101]  = 1'b1;
    buffer_full_rands[102]  = 1'b0;
    buffer_full_rands[103]  = 1'b0;
    buffer_full_rands[104]  = 1'b0;
    buffer_full_rands[105]  = 1'b0;
    buffer_full_rands[106]  = 1'b1;
    buffer_full_rands[107]  = 1'b0;
    buffer_full_rands[108]  = 1'b0;
    buffer_full_rands[109]  = 1'b0;
    buffer_full_rands[110]  = 1'b1;
    buffer_full_rands[111]  = 1'b0;
    buffer_full_rands[112]  = 1'b0;
    buffer_full_rands[113]  = 1'b0;
    buffer_full_rands[114]  = 1'b0;
    buffer_full_rands[115]  = 1'b1;
    buffer_full_rands[116]  = 1'b0;
    buffer_full_rands[117]  = 1'b1;
    buffer_full_rands[118]  = 1'b0;
    buffer_full_rands[119]  = 1'b1;
    buffer_full_rands[120]  = 1'b0;
    buffer_full_rands[121]  = 1'b1;
    buffer_full_rands[122]  = 1'b0;
    buffer_full_rands[123]  = 1'b1;
    buffer_full_rands[124]  = 1'b1;
    buffer_full_rands[125]  = 1'b0;
    buffer_full_rands[126]  = 1'b0;
    buffer_full_rands[127]  = 1'b1;
    buffer_full_rands[128]  = 1'b0;
    buffer_full_rands[129]  = 1'b0;
    buffer_full_rands[130]  = 1'b1;
    buffer_full_rands[131]  = 1'b1;
    buffer_full_rands[132]  = 1'b0;
    buffer_full_rands[133]  = 1'b0;
    buffer_full_rands[134]  = 1'b0;
    buffer_full_rands[135]  = 1'b1;
    buffer_full_rands[136]  = 1'b1;
    buffer_full_rands[137]  = 1'b1;
    buffer_full_rands[138]  = 1'b0;
    buffer_full_rands[139]  = 1'b0;
    buffer_full_rands[140]  = 1'b1;
    buffer_full_rands[141]  = 1'b0;
    buffer_full_rands[142]  = 1'b1;
    buffer_full_rands[143]  = 1'b0;
    buffer_full_rands[144]  = 1'b0;
    buffer_full_rands[145]  = 1'b0;
    buffer_full_rands[146]  = 1'b0;
    buffer_full_rands[147]  = 1'b0;
    buffer_full_rands[148]  = 1'b0;
    buffer_full_rands[149]  = 1'b0;
    buffer_full_rands[150]  = 1'b1;
    buffer_full_rands[151]  = 1'b0;
    buffer_full_rands[152]  = 1'b1;
    buffer_full_rands[153]  = 1'b0;
    buffer_full_rands[154]  = 1'b1;
    buffer_full_rands[155]  = 1'b1;
    buffer_full_rands[156]  = 1'b1;
    buffer_full_rands[157]  = 1'b1;
    buffer_full_rands[158]  = 1'b1;
    buffer_full_rands[159]  = 1'b0;
    buffer_full_rands[160]  = 1'b1;
    buffer_full_rands[161]  = 1'b0;
    buffer_full_rands[162]  = 1'b0;
    buffer_full_rands[163]  = 1'b0;
    buffer_full_rands[164]  = 1'b0;
    buffer_full_rands[165]  = 1'b0;
    buffer_full_rands[166]  = 1'b1;
    buffer_full_rands[167]  = 1'b0;
    buffer_full_rands[168]  = 1'b0;
    buffer_full_rands[169]  = 1'b0;
    buffer_full_rands[170]  = 1'b1;
    buffer_full_rands[171]  = 1'b0;
    buffer_full_rands[172]  = 1'b1;
    buffer_full_rands[173]  = 1'b1;
    buffer_full_rands[174]  = 1'b0;
    buffer_full_rands[175]  = 1'b1;
    buffer_full_rands[176]  = 1'b0;
    buffer_full_rands[177]  = 1'b1;
    buffer_full_rands[178]  = 1'b1;
    buffer_full_rands[179]  = 1'b0;
    buffer_full_rands[180]  = 1'b0;
    buffer_full_rands[181]  = 1'b0;
    buffer_full_rands[182]  = 1'b1;
    buffer_full_rands[183]  = 1'b0;
    buffer_full_rands[184]  = 1'b0;
    buffer_full_rands[185]  = 1'b0;
    buffer_full_rands[186]  = 1'b1;
    buffer_full_rands[187]  = 1'b1;
    buffer_full_rands[188]  = 1'b1;
    buffer_full_rands[189]  = 1'b0;
    buffer_full_rands[190]  = 1'b0;
    buffer_full_rands[191]  = 1'b0;
    buffer_full_rands[192]  = 1'b1;
    buffer_full_rands[193]  = 1'b0;
    buffer_full_rands[194]  = 1'b1;
    buffer_full_rands[195]  = 1'b1;
    buffer_full_rands[196]  = 1'b1;
    buffer_full_rands[197]  = 1'b0;
    buffer_full_rands[198]  = 1'b1;
    buffer_full_rands[199]  = 1'b1;
    buffer_full_rands[200]  = 1'b0;
    buffer_full_rands[201]  = 1'b1;
    buffer_full_rands[202]  = 1'b0;
    buffer_full_rands[203]  = 1'b1;
    buffer_full_rands[204]  = 1'b1;
    buffer_full_rands[205]  = 1'b1;
    buffer_full_rands[206]  = 1'b0;
    buffer_full_rands[207]  = 1'b1;
    buffer_full_rands[208]  = 1'b0;
    buffer_full_rands[209]  = 1'b1;
    buffer_full_rands[210]  = 1'b1;
    buffer_full_rands[211]  = 1'b0;
    buffer_full_rands[212]  = 1'b1;
    buffer_full_rands[213]  = 1'b1;
    buffer_full_rands[214]  = 1'b1;
    buffer_full_rands[215]  = 1'b0;
    buffer_full_rands[216]  = 1'b1;
    buffer_full_rands[217]  = 1'b0;
    buffer_full_rands[218]  = 1'b1;
    buffer_full_rands[219]  = 1'b0;
    buffer_full_rands[220]  = 1'b0;
    buffer_full_rands[221]  = 1'b1;
    buffer_full_rands[222]  = 1'b0;
    buffer_full_rands[223]  = 1'b1;
    buffer_full_rands[224]  = 1'b0;
    buffer_full_rands[225]  = 1'b0;
    buffer_full_rands[226]  = 1'b1;
    buffer_full_rands[227]  = 1'b0;
    buffer_full_rands[228]  = 1'b1;
    buffer_full_rands[229]  = 1'b1;
    buffer_full_rands[230]  = 1'b0;
    buffer_full_rands[231]  = 1'b1;
    buffer_full_rands[232]  = 1'b1;
    buffer_full_rands[233]  = 1'b1;
    buffer_full_rands[234]  = 1'b1;
    buffer_full_rands[235]  = 1'b1;
    buffer_full_rands[236]  = 1'b1;
    buffer_full_rands[237]  = 1'b0;
    buffer_full_rands[238]  = 1'b1;
    buffer_full_rands[239]  = 1'b1;
    buffer_full_rands[240]  = 1'b0;
    buffer_full_rands[241]  = 1'b0;
    buffer_full_rands[242]  = 1'b0;
    buffer_full_rands[243]  = 1'b0;
    buffer_full_rands[244]  = 1'b1;
    buffer_full_rands[245]  = 1'b1;
    buffer_full_rands[246]  = 1'b1;
    buffer_full_rands[247]  = 1'b0;
    buffer_full_rands[248]  = 1'b1;
    buffer_full_rands[249]  = 1'b0;
    buffer_full_rands[250]  = 1'b1;
    buffer_full_rands[251]  = 1'b1;
    buffer_full_rands[252]  = 1'b1;
    buffer_full_rands[253]  = 1'b0;
    buffer_full_rands[254]  = 1'b1;
    buffer_full_rands[255]  = 1'b0;
    buffer_full_rands[256]  = 1'b1;
    buffer_full_rands[257]  = 1'b1;
    buffer_full_rands[258]  = 1'b1;
    buffer_full_rands[259]  = 1'b1;
    buffer_full_rands[260]  = 1'b0;
    buffer_full_rands[261]  = 1'b1;
    buffer_full_rands[262]  = 1'b1;
    buffer_full_rands[263]  = 1'b1;
    buffer_full_rands[264]  = 1'b0;
    buffer_full_rands[265]  = 1'b0;
    buffer_full_rands[266]  = 1'b0;
    buffer_full_rands[267]  = 1'b0;
    buffer_full_rands[268]  = 1'b0;
    buffer_full_rands[269]  = 1'b1;
    buffer_full_rands[270]  = 1'b1;
    buffer_full_rands[271]  = 1'b0;
    buffer_full_rands[272]  = 1'b1;
    buffer_full_rands[273]  = 1'b1;
    buffer_full_rands[274]  = 1'b1;
    buffer_full_rands[275]  = 1'b0;
    buffer_full_rands[276]  = 1'b1;
    buffer_full_rands[277]  = 1'b1;
    buffer_full_rands[278]  = 1'b0;
    buffer_full_rands[279]  = 1'b0;
    buffer_full_rands[280]  = 1'b0;
    buffer_full_rands[281]  = 1'b0;
    buffer_full_rands[282]  = 1'b1;
    buffer_full_rands[283]  = 1'b0;
    buffer_full_rands[284]  = 1'b1;
    buffer_full_rands[285]  = 1'b0;
    buffer_full_rands[286]  = 1'b0;
    buffer_full_rands[287]  = 1'b0;
    buffer_full_rands[288]  = 1'b1;
    buffer_full_rands[289]  = 1'b1;
    buffer_full_rands[290]  = 1'b0;
    buffer_full_rands[291]  = 1'b0;
    buffer_full_rands[292]  = 1'b1;
    buffer_full_rands[293]  = 1'b0;
    buffer_full_rands[294]  = 1'b1;
    buffer_full_rands[295]  = 1'b1;
    buffer_full_rands[296]  = 1'b1;
    buffer_full_rands[297]  = 1'b0;
    buffer_full_rands[298]  = 1'b1;
    buffer_full_rands[299]  = 1'b1;
    buffer_full_rands[300]  = 1'b1;
    buffer_full_rands[301]  = 1'b1;
    buffer_full_rands[302]  = 1'b0;
    buffer_full_rands[303]  = 1'b1;
    buffer_full_rands[304]  = 1'b0;
    buffer_full_rands[305]  = 1'b0;
    buffer_full_rands[306]  = 1'b1;
    buffer_full_rands[307]  = 1'b0;
    buffer_full_rands[308]  = 1'b0;
    buffer_full_rands[309]  = 1'b1;
    buffer_full_rands[310]  = 1'b0;
    buffer_full_rands[311]  = 1'b1;
    buffer_full_rands[312]  = 1'b1;
    buffer_full_rands[313]  = 1'b1;
    buffer_full_rands[314]  = 1'b1;
    buffer_full_rands[315]  = 1'b0;
    buffer_full_rands[316]  = 1'b0;
    buffer_full_rands[317]  = 1'b0;
    buffer_full_rands[318]  = 1'b0;
    buffer_full_rands[319]  = 1'b1;
    buffer_full_rands[320]  = 1'b1;
    buffer_full_rands[321]  = 1'b1;
    buffer_full_rands[322]  = 1'b0;
    buffer_full_rands[323]  = 1'b1;
    buffer_full_rands[324]  = 1'b1;
    buffer_full_rands[325]  = 1'b1;
    buffer_full_rands[326]  = 1'b0;
    buffer_full_rands[327]  = 1'b1;
    buffer_full_rands[328]  = 1'b1;
    buffer_full_rands[329]  = 1'b1;
    buffer_full_rands[330]  = 1'b1;
    buffer_full_rands[331]  = 1'b1;
    buffer_full_rands[332]  = 1'b1;
    buffer_full_rands[333]  = 1'b1;
    buffer_full_rands[334]  = 1'b0;
    buffer_full_rands[335]  = 1'b1;
    buffer_full_rands[336]  = 1'b0;
    buffer_full_rands[337]  = 1'b1;
    buffer_full_rands[338]  = 1'b0;
    buffer_full_rands[339]  = 1'b0;
    buffer_full_rands[340]  = 1'b0;
    buffer_full_rands[341]  = 1'b1;
    buffer_full_rands[342]  = 1'b0;
    buffer_full_rands[343]  = 1'b1;
    buffer_full_rands[344]  = 1'b0;
    buffer_full_rands[345]  = 1'b0;
    buffer_full_rands[346]  = 1'b1;
    buffer_full_rands[347]  = 1'b0;
    buffer_full_rands[348]  = 1'b1;
    buffer_full_rands[349]  = 1'b0;
    buffer_full_rands[350]  = 1'b1;
    buffer_full_rands[351]  = 1'b0;
    buffer_full_rands[352]  = 1'b0;
    buffer_full_rands[353]  = 1'b0;
    buffer_full_rands[354]  = 1'b0;
    buffer_full_rands[355]  = 1'b0;
    buffer_full_rands[356]  = 1'b0;
    buffer_full_rands[357]  = 1'b1;
    buffer_full_rands[358]  = 1'b0;
    buffer_full_rands[359]  = 1'b1;
    buffer_full_rands[360]  = 1'b1;
    buffer_full_rands[361]  = 1'b1;
    buffer_full_rands[362]  = 1'b0;
    buffer_full_rands[363]  = 1'b1;
    buffer_full_rands[364]  = 1'b0;
    buffer_full_rands[365]  = 1'b1;
    buffer_full_rands[366]  = 1'b1;
    buffer_full_rands[367]  = 1'b1;
    buffer_full_rands[368]  = 1'b0;
    buffer_full_rands[369]  = 1'b1;
    buffer_full_rands[370]  = 1'b1;
    buffer_full_rands[371]  = 1'b1;
    buffer_full_rands[372]  = 1'b0;
    buffer_full_rands[373]  = 1'b0;
    buffer_full_rands[374]  = 1'b0;
    buffer_full_rands[375]  = 1'b0;
    buffer_full_rands[376]  = 1'b0;
    buffer_full_rands[377]  = 1'b0;
    buffer_full_rands[378]  = 1'b1;
    buffer_full_rands[379]  = 1'b1;
    buffer_full_rands[380]  = 1'b0;
    buffer_full_rands[381]  = 1'b0;
    buffer_full_rands[382]  = 1'b0;
    buffer_full_rands[383]  = 1'b0;
    buffer_full_rands[384]  = 1'b0;
    buffer_full_rands[385]  = 1'b1;
    buffer_full_rands[386]  = 1'b1;
    buffer_full_rands[387]  = 1'b0;
    buffer_full_rands[388]  = 1'b0;
    buffer_full_rands[389]  = 1'b1;
    buffer_full_rands[390]  = 1'b0;
    buffer_full_rands[391]  = 1'b1;
    buffer_full_rands[392]  = 1'b0;
    buffer_full_rands[393]  = 1'b1;
    buffer_full_rands[394]  = 1'b1;
    buffer_full_rands[395]  = 1'b1;
    buffer_full_rands[396]  = 1'b1;
    buffer_full_rands[397]  = 1'b1;
    buffer_full_rands[398]  = 1'b0;
    buffer_full_rands[399]  = 1'b1;
    buffer_full_rands[400]  = 1'b1;
    buffer_full_rands[401]  = 1'b1;
    buffer_full_rands[402]  = 1'b1;
    buffer_full_rands[403]  = 1'b1;
    buffer_full_rands[404]  = 1'b1;
    buffer_full_rands[405]  = 1'b1;
    buffer_full_rands[406]  = 1'b1;
    buffer_full_rands[407]  = 1'b0;
    buffer_full_rands[408]  = 1'b0;
    buffer_full_rands[409]  = 1'b0;
    buffer_full_rands[410]  = 1'b1;
    buffer_full_rands[411]  = 1'b0;
    buffer_full_rands[412]  = 1'b0;
    buffer_full_rands[413]  = 1'b0;
    buffer_full_rands[414]  = 1'b1;
    buffer_full_rands[415]  = 1'b1;
    buffer_full_rands[416]  = 1'b1;
    buffer_full_rands[417]  = 1'b0;
    buffer_full_rands[418]  = 1'b1;
    buffer_full_rands[419]  = 1'b1;
    buffer_full_rands[420]  = 1'b1;
    buffer_full_rands[421]  = 1'b0;
    buffer_full_rands[422]  = 1'b0;
    buffer_full_rands[423]  = 1'b1;
    buffer_full_rands[424]  = 1'b1;
    buffer_full_rands[425]  = 1'b0;
    buffer_full_rands[426]  = 1'b0;
    buffer_full_rands[427]  = 1'b0;
    buffer_full_rands[428]  = 1'b1;
    buffer_full_rands[429]  = 1'b0;
    buffer_full_rands[430]  = 1'b1;
    buffer_full_rands[431]  = 1'b1;
    buffer_full_rands[432]  = 1'b0;
    buffer_full_rands[433]  = 1'b1;
    buffer_full_rands[434]  = 1'b0;
    buffer_full_rands[435]  = 1'b1;
    buffer_full_rands[436]  = 1'b1;
    buffer_full_rands[437]  = 1'b0;
    buffer_full_rands[438]  = 1'b0;
    buffer_full_rands[439]  = 1'b1;
    buffer_full_rands[440]  = 1'b0;
    buffer_full_rands[441]  = 1'b1;
    buffer_full_rands[442]  = 1'b1;
    buffer_full_rands[443]  = 1'b0;
    buffer_full_rands[444]  = 1'b0;
    buffer_full_rands[445]  = 1'b0;
    buffer_full_rands[446]  = 1'b0;
    buffer_full_rands[447]  = 1'b1;
    buffer_full_rands[448]  = 1'b0;
    buffer_full_rands[449]  = 1'b1;
    buffer_full_rands[450]  = 1'b0;
    buffer_full_rands[451]  = 1'b0;
    buffer_full_rands[452]  = 1'b1;
    buffer_full_rands[453]  = 1'b0;
    buffer_full_rands[454]  = 1'b0;
    buffer_full_rands[455]  = 1'b1;
    buffer_full_rands[456]  = 1'b0;
    buffer_full_rands[457]  = 1'b0;
    buffer_full_rands[458]  = 1'b0;
    buffer_full_rands[459]  = 1'b0;
    buffer_full_rands[460]  = 1'b0;
    buffer_full_rands[461]  = 1'b0;
    buffer_full_rands[462]  = 1'b1;
    buffer_full_rands[463]  = 1'b1;
    buffer_full_rands[464]  = 1'b0;
    buffer_full_rands[465]  = 1'b1;
    buffer_full_rands[466]  = 1'b1;
    buffer_full_rands[467]  = 1'b0;
    buffer_full_rands[468]  = 1'b0;
    buffer_full_rands[469]  = 1'b0;
    buffer_full_rands[470]  = 1'b0;
    buffer_full_rands[471]  = 1'b0;
    buffer_full_rands[472]  = 1'b0;
    buffer_full_rands[473]  = 1'b1;
    buffer_full_rands[474]  = 1'b0;
    buffer_full_rands[475]  = 1'b1;
    buffer_full_rands[476]  = 1'b0;
    buffer_full_rands[477]  = 1'b0;
    buffer_full_rands[478]  = 1'b1;
    buffer_full_rands[479]  = 1'b1;
    buffer_full_rands[480]  = 1'b1;
    buffer_full_rands[481]  = 1'b0;
    buffer_full_rands[482]  = 1'b0;
    buffer_full_rands[483]  = 1'b0;
    buffer_full_rands[484]  = 1'b1;
    buffer_full_rands[485]  = 1'b0;
    buffer_full_rands[486]  = 1'b1;
    buffer_full_rands[487]  = 1'b1;
    buffer_full_rands[488]  = 1'b0;
    buffer_full_rands[489]  = 1'b1;
    buffer_full_rands[490]  = 1'b0;
    buffer_full_rands[491]  = 1'b0;
    buffer_full_rands[492]  = 1'b0;
    buffer_full_rands[493]  = 1'b1;
    buffer_full_rands[494]  = 1'b1;
    buffer_full_rands[495]  = 1'b1;
    buffer_full_rands[496]  = 1'b1;
    buffer_full_rands[497]  = 1'b0;
    buffer_full_rands[498]  = 1'b1;
    buffer_full_rands[499]  = 1'b0;
    buffer_full_rands[500]  = 1'b0;
    buffer_full_rands[501]  = 1'b1;
    buffer_full_rands[502]  = 1'b0;
    buffer_full_rands[503]  = 1'b0;
    buffer_full_rands[504]  = 1'b1;
    buffer_full_rands[505]  = 1'b0;
    buffer_full_rands[506]  = 1'b0;
    buffer_full_rands[507]  = 1'b0;
    buffer_full_rands[508]  = 1'b0;
    buffer_full_rands[509]  = 1'b0;
    buffer_full_rands[510]  = 1'b1;
    buffer_full_rands[511]  = 1'b0;
    buffer_full_rands[512]  = 1'b0;
    buffer_full_rands[513]  = 1'b1;
    buffer_full_rands[514]  = 1'b1;
    buffer_full_rands[515]  = 1'b1;
    buffer_full_rands[516]  = 1'b1;
    buffer_full_rands[517]  = 1'b0;
    buffer_full_rands[518]  = 1'b0;
    buffer_full_rands[519]  = 1'b1;
    buffer_full_rands[520]  = 1'b1;
    buffer_full_rands[521]  = 1'b1;
    buffer_full_rands[522]  = 1'b0;
    buffer_full_rands[523]  = 1'b1;
    buffer_full_rands[524]  = 1'b1;
    buffer_full_rands[525]  = 1'b0;
    buffer_full_rands[526]  = 1'b1;
    buffer_full_rands[527]  = 1'b0;
    buffer_full_rands[528]  = 1'b1;
    buffer_full_rands[529]  = 1'b1;
    buffer_full_rands[530]  = 1'b1;
    buffer_full_rands[531]  = 1'b0;
    buffer_full_rands[532]  = 1'b0;
    buffer_full_rands[533]  = 1'b0;
    buffer_full_rands[534]  = 1'b0;
    buffer_full_rands[535]  = 1'b0;
    buffer_full_rands[536]  = 1'b1;
    buffer_full_rands[537]  = 1'b0;
    buffer_full_rands[538]  = 1'b0;
    buffer_full_rands[539]  = 1'b0;
    buffer_full_rands[540]  = 1'b0;
    buffer_full_rands[541]  = 1'b0;
    buffer_full_rands[542]  = 1'b1;
    buffer_full_rands[543]  = 1'b1;
    buffer_full_rands[544]  = 1'b0;
    buffer_full_rands[545]  = 1'b1;
    buffer_full_rands[546]  = 1'b1;
    buffer_full_rands[547]  = 1'b1;
    buffer_full_rands[548]  = 1'b0;
    buffer_full_rands[549]  = 1'b0;
    buffer_full_rands[550]  = 1'b0;
    buffer_full_rands[551]  = 1'b1;
    buffer_full_rands[552]  = 1'b0;
    buffer_full_rands[553]  = 1'b0;
    buffer_full_rands[554]  = 1'b0;
    buffer_full_rands[555]  = 1'b1;
    buffer_full_rands[556]  = 1'b1;
    buffer_full_rands[557]  = 1'b1;
    buffer_full_rands[558]  = 1'b1;
    buffer_full_rands[559]  = 1'b1;
    buffer_full_rands[560]  = 1'b1;
    buffer_full_rands[561]  = 1'b1;
    buffer_full_rands[562]  = 1'b0;
    buffer_full_rands[563]  = 1'b1;
    buffer_full_rands[564]  = 1'b0;
    buffer_full_rands[565]  = 1'b0;
    buffer_full_rands[566]  = 1'b0;
    buffer_full_rands[567]  = 1'b1;
    buffer_full_rands[568]  = 1'b0;
    buffer_full_rands[569]  = 1'b0;
    buffer_full_rands[570]  = 1'b1;
    buffer_full_rands[571]  = 1'b1;
    buffer_full_rands[572]  = 1'b0;
    buffer_full_rands[573]  = 1'b0;
    buffer_full_rands[574]  = 1'b0;
    buffer_full_rands[575]  = 1'b1;
    buffer_full_rands[576]  = 1'b1;
    buffer_full_rands[577]  = 1'b1;
    buffer_full_rands[578]  = 1'b0;
    buffer_full_rands[579]  = 1'b0;
    buffer_full_rands[580]  = 1'b0;
    buffer_full_rands[581]  = 1'b1;
    buffer_full_rands[582]  = 1'b0;
    buffer_full_rands[583]  = 1'b1;
    buffer_full_rands[584]  = 1'b1;
    buffer_full_rands[585]  = 1'b0;
    buffer_full_rands[586]  = 1'b0;
    buffer_full_rands[587]  = 1'b0;
    buffer_full_rands[588]  = 1'b0;
    buffer_full_rands[589]  = 1'b1;
    buffer_full_rands[590]  = 1'b0;
    buffer_full_rands[591]  = 1'b1;
    buffer_full_rands[592]  = 1'b0;
    buffer_full_rands[593]  = 1'b1;
    buffer_full_rands[594]  = 1'b1;
    buffer_full_rands[595]  = 1'b1;
    buffer_full_rands[596]  = 1'b1;
    buffer_full_rands[597]  = 1'b0;
    buffer_full_rands[598]  = 1'b0;
    buffer_full_rands[599]  = 1'b0;
    buffer_full_rands[600]  = 1'b1;
    buffer_full_rands[601]  = 1'b1;
    buffer_full_rands[602]  = 1'b1;
    buffer_full_rands[603]  = 1'b0;
    buffer_full_rands[604]  = 1'b0;
    buffer_full_rands[605]  = 1'b0;
    buffer_full_rands[606]  = 1'b0;
    buffer_full_rands[607]  = 1'b0;
    buffer_full_rands[608]  = 1'b1;
    buffer_full_rands[609]  = 1'b0;
    buffer_full_rands[610]  = 1'b1;
    buffer_full_rands[611]  = 1'b1;
    buffer_full_rands[612]  = 1'b0;
    buffer_full_rands[613]  = 1'b1;
    buffer_full_rands[614]  = 1'b1;
    buffer_full_rands[615]  = 1'b1;
    buffer_full_rands[616]  = 1'b1;
    buffer_full_rands[617]  = 1'b1;
    buffer_full_rands[618]  = 1'b1;
    buffer_full_rands[619]  = 1'b1;
    buffer_full_rands[620]  = 1'b0;
    buffer_full_rands[621]  = 1'b1;
    buffer_full_rands[622]  = 1'b1;
    buffer_full_rands[623]  = 1'b0;
    buffer_full_rands[624]  = 1'b0;
    buffer_full_rands[625]  = 1'b0;
    buffer_full_rands[626]  = 1'b0;
    buffer_full_rands[627]  = 1'b0;
    buffer_full_rands[628]  = 1'b0;
    buffer_full_rands[629]  = 1'b0;
    buffer_full_rands[630]  = 1'b1;
    buffer_full_rands[631]  = 1'b1;
    buffer_full_rands[632]  = 1'b0;
    buffer_full_rands[633]  = 1'b0;
    buffer_full_rands[634]  = 1'b0;
    buffer_full_rands[635]  = 1'b0;
    buffer_full_rands[636]  = 1'b1;
    buffer_full_rands[637]  = 1'b1;
    buffer_full_rands[638]  = 1'b0;
    buffer_full_rands[639]  = 1'b0;
    buffer_full_rands[640]  = 1'b1;
    buffer_full_rands[641]  = 1'b0;
    buffer_full_rands[642]  = 1'b0;
    buffer_full_rands[643]  = 1'b0;
    buffer_full_rands[644]  = 1'b1;
    buffer_full_rands[645]  = 1'b0;
    buffer_full_rands[646]  = 1'b0;
    buffer_full_rands[647]  = 1'b1;
    buffer_full_rands[648]  = 1'b0;
    buffer_full_rands[649]  = 1'b0;
    buffer_full_rands[650]  = 1'b1;
    buffer_full_rands[651]  = 1'b1;
    buffer_full_rands[652]  = 1'b1;
    buffer_full_rands[653]  = 1'b0;
    buffer_full_rands[654]  = 1'b1;
    buffer_full_rands[655]  = 1'b1;
    buffer_full_rands[656]  = 1'b0;
    buffer_full_rands[657]  = 1'b0;
    buffer_full_rands[658]  = 1'b1;
    buffer_full_rands[659]  = 1'b1;
    buffer_full_rands[660]  = 1'b1;
    buffer_full_rands[661]  = 1'b1;
    buffer_full_rands[662]  = 1'b1;
    buffer_full_rands[663]  = 1'b0;
    buffer_full_rands[664]  = 1'b1;
    buffer_full_rands[665]  = 1'b1;
    buffer_full_rands[666]  = 1'b0;
    buffer_full_rands[667]  = 1'b1;
    buffer_full_rands[668]  = 1'b0;
    buffer_full_rands[669]  = 1'b0;
    buffer_full_rands[670]  = 1'b1;
    buffer_full_rands[671]  = 1'b1;
    buffer_full_rands[672]  = 1'b0;
    buffer_full_rands[673]  = 1'b0;
    buffer_full_rands[674]  = 1'b0;
    buffer_full_rands[675]  = 1'b0;
    buffer_full_rands[676]  = 1'b0;
    buffer_full_rands[677]  = 1'b1;
    buffer_full_rands[678]  = 1'b1;
    buffer_full_rands[679]  = 1'b0;
    buffer_full_rands[680]  = 1'b1;
    buffer_full_rands[681]  = 1'b1;
    buffer_full_rands[682]  = 1'b1;
    buffer_full_rands[683]  = 1'b1;
    buffer_full_rands[684]  = 1'b1;
    buffer_full_rands[685]  = 1'b1;
    buffer_full_rands[686]  = 1'b1;
    buffer_full_rands[687]  = 1'b0;
    buffer_full_rands[688]  = 1'b0;
    buffer_full_rands[689]  = 1'b1;
    buffer_full_rands[690]  = 1'b1;
    buffer_full_rands[691]  = 1'b0;
    buffer_full_rands[692]  = 1'b0;
    buffer_full_rands[693]  = 1'b0;
    buffer_full_rands[694]  = 1'b1;
    buffer_full_rands[695]  = 1'b0;
    buffer_full_rands[696]  = 1'b0;
    buffer_full_rands[697]  = 1'b1;
    buffer_full_rands[698]  = 1'b1;
    buffer_full_rands[699]  = 1'b0;
    buffer_full_rands[700]  = 1'b0;
    buffer_full_rands[701]  = 1'b0;
    buffer_full_rands[702]  = 1'b0;
    buffer_full_rands[703]  = 1'b0;
    buffer_full_rands[704]  = 1'b0;
    buffer_full_rands[705]  = 1'b0;
    buffer_full_rands[706]  = 1'b1;
    buffer_full_rands[707]  = 1'b1;
    buffer_full_rands[708]  = 1'b1;
    buffer_full_rands[709]  = 1'b1;
    buffer_full_rands[710]  = 1'b0;
    buffer_full_rands[711]  = 1'b1;
    buffer_full_rands[712]  = 1'b0;
    buffer_full_rands[713]  = 1'b0;
    buffer_full_rands[714]  = 1'b0;
    buffer_full_rands[715]  = 1'b0;
    buffer_full_rands[716]  = 1'b1;
    buffer_full_rands[717]  = 1'b0;
    buffer_full_rands[718]  = 1'b0;
    buffer_full_rands[719]  = 1'b1;
    buffer_full_rands[720]  = 1'b1;
    buffer_full_rands[721]  = 1'b0;
    buffer_full_rands[722]  = 1'b1;
    buffer_full_rands[723]  = 1'b0;
    buffer_full_rands[724]  = 1'b0;
    buffer_full_rands[725]  = 1'b0;
    buffer_full_rands[726]  = 1'b1;
    buffer_full_rands[727]  = 1'b1;
    buffer_full_rands[728]  = 1'b1;
    buffer_full_rands[729]  = 1'b0;
    buffer_full_rands[730]  = 1'b1;
    buffer_full_rands[731]  = 1'b1;
    buffer_full_rands[732]  = 1'b0;
    buffer_full_rands[733]  = 1'b1;
    buffer_full_rands[734]  = 1'b0;
    buffer_full_rands[735]  = 1'b1;
    buffer_full_rands[736]  = 1'b1;
    buffer_full_rands[737]  = 1'b0;
    buffer_full_rands[738]  = 1'b1;
    buffer_full_rands[739]  = 1'b1;
    buffer_full_rands[740]  = 1'b0;
    buffer_full_rands[741]  = 1'b1;
    buffer_full_rands[742]  = 1'b0;
    buffer_full_rands[743]  = 1'b0;
    buffer_full_rands[744]  = 1'b0;
    buffer_full_rands[745]  = 1'b0;
    buffer_full_rands[746]  = 1'b1;
    buffer_full_rands[747]  = 1'b0;
    buffer_full_rands[748]  = 1'b0;
    buffer_full_rands[749]  = 1'b1;
    buffer_full_rands[750]  = 1'b1;
    buffer_full_rands[751]  = 1'b0;
    buffer_full_rands[752]  = 1'b0;
    buffer_full_rands[753]  = 1'b0;
    buffer_full_rands[754]  = 1'b0;
    buffer_full_rands[755]  = 1'b1;
    buffer_full_rands[756]  = 1'b0;
    buffer_full_rands[757]  = 1'b0;
    buffer_full_rands[758]  = 1'b1;
    buffer_full_rands[759]  = 1'b1;
    buffer_full_rands[760]  = 1'b0;
    buffer_full_rands[761]  = 1'b1;
    buffer_full_rands[762]  = 1'b1;
    buffer_full_rands[763]  = 1'b1;
    buffer_full_rands[764]  = 1'b1;
    buffer_full_rands[765]  = 1'b1;
    buffer_full_rands[766]  = 1'b0;
    buffer_full_rands[767]  = 1'b0;
    buffer_full_rands[768]  = 1'b1;
    buffer_full_rands[769]  = 1'b0;
    buffer_full_rands[770]  = 1'b1;
    buffer_full_rands[771]  = 1'b0;
    buffer_full_rands[772]  = 1'b0;
    buffer_full_rands[773]  = 1'b1;
    buffer_full_rands[774]  = 1'b1;
    buffer_full_rands[775]  = 1'b1;
    buffer_full_rands[776]  = 1'b0;
    buffer_full_rands[777]  = 1'b1;
    buffer_full_rands[778]  = 1'b1;
    buffer_full_rands[779]  = 1'b0;
    buffer_full_rands[780]  = 1'b1;
    buffer_full_rands[781]  = 1'b1;
    buffer_full_rands[782]  = 1'b1;
    buffer_full_rands[783]  = 1'b0;
    buffer_full_rands[784]  = 1'b0;
    buffer_full_rands[785]  = 1'b1;
    buffer_full_rands[786]  = 1'b0;
    buffer_full_rands[787]  = 1'b0;
    buffer_full_rands[788]  = 1'b1;
    buffer_full_rands[789]  = 1'b0;
    buffer_full_rands[790]  = 1'b1;
    buffer_full_rands[791]  = 1'b0;
    buffer_full_rands[792]  = 1'b1;
    buffer_full_rands[793]  = 1'b1;
    buffer_full_rands[794]  = 1'b0;
    buffer_full_rands[795]  = 1'b1;
    buffer_full_rands[796]  = 1'b0;
    buffer_full_rands[797]  = 1'b1;
    buffer_full_rands[798]  = 1'b1;
    buffer_full_rands[799]  = 1'b0;
    buffer_full_rands[800]  = 1'b1;
    buffer_full_rands[801]  = 1'b1;
    buffer_full_rands[802]  = 1'b1;
    buffer_full_rands[803]  = 1'b1;
    buffer_full_rands[804]  = 1'b1;
    buffer_full_rands[805]  = 1'b1;
    buffer_full_rands[806]  = 1'b0;
    buffer_full_rands[807]  = 1'b1;
    buffer_full_rands[808]  = 1'b1;
    buffer_full_rands[809]  = 1'b0;
    buffer_full_rands[810]  = 1'b0;
    buffer_full_rands[811]  = 1'b1;
    buffer_full_rands[812]  = 1'b0;
    buffer_full_rands[813]  = 1'b0;
    buffer_full_rands[814]  = 1'b1;
    buffer_full_rands[815]  = 1'b0;
    buffer_full_rands[816]  = 1'b1;
    buffer_full_rands[817]  = 1'b1;
    buffer_full_rands[818]  = 1'b0;
    buffer_full_rands[819]  = 1'b1;
    buffer_full_rands[820]  = 1'b1;
    buffer_full_rands[821]  = 1'b1;
    buffer_full_rands[822]  = 1'b1;
    buffer_full_rands[823]  = 1'b1;
    buffer_full_rands[824]  = 1'b0;
    buffer_full_rands[825]  = 1'b0;
    buffer_full_rands[826]  = 1'b1;
    buffer_full_rands[827]  = 1'b0;
    buffer_full_rands[828]  = 1'b1;
    buffer_full_rands[829]  = 1'b0;
    buffer_full_rands[830]  = 1'b0;
    buffer_full_rands[831]  = 1'b1;
    buffer_full_rands[832]  = 1'b0;
    buffer_full_rands[833]  = 1'b0;
    buffer_full_rands[834]  = 1'b1;
    buffer_full_rands[835]  = 1'b0;
    buffer_full_rands[836]  = 1'b0;
    buffer_full_rands[837]  = 1'b1;
    buffer_full_rands[838]  = 1'b1;
    buffer_full_rands[839]  = 1'b1;
    buffer_full_rands[840]  = 1'b0;
    buffer_full_rands[841]  = 1'b1;
    buffer_full_rands[842]  = 1'b0;
    buffer_full_rands[843]  = 1'b0;
    buffer_full_rands[844]  = 1'b1;
    buffer_full_rands[845]  = 1'b0;
    buffer_full_rands[846]  = 1'b1;
    buffer_full_rands[847]  = 1'b1;
    buffer_full_rands[848]  = 1'b0;
    buffer_full_rands[849]  = 1'b0;
    buffer_full_rands[850]  = 1'b1;
    buffer_full_rands[851]  = 1'b0;
    buffer_full_rands[852]  = 1'b1;
    buffer_full_rands[853]  = 1'b1;
    buffer_full_rands[854]  = 1'b1;
    buffer_full_rands[855]  = 1'b0;
    buffer_full_rands[856]  = 1'b1;
    buffer_full_rands[857]  = 1'b0;
    buffer_full_rands[858]  = 1'b0;
    buffer_full_rands[859]  = 1'b0;
    buffer_full_rands[860]  = 1'b1;
    buffer_full_rands[861]  = 1'b0;
    buffer_full_rands[862]  = 1'b1;
    buffer_full_rands[863]  = 1'b0;
    buffer_full_rands[864]  = 1'b0;
    buffer_full_rands[865]  = 1'b1;
    buffer_full_rands[866]  = 1'b0;
    buffer_full_rands[867]  = 1'b0;
    buffer_full_rands[868]  = 1'b1;
    buffer_full_rands[869]  = 1'b1;
    buffer_full_rands[870]  = 1'b1;
    buffer_full_rands[871]  = 1'b0;
    buffer_full_rands[872]  = 1'b0;
    buffer_full_rands[873]  = 1'b1;
    buffer_full_rands[874]  = 1'b1;
    buffer_full_rands[875]  = 1'b1;
    buffer_full_rands[876]  = 1'b0;
    buffer_full_rands[877]  = 1'b0;
    buffer_full_rands[878]  = 1'b1;
    buffer_full_rands[879]  = 1'b1;
    buffer_full_rands[880]  = 1'b1;
    buffer_full_rands[881]  = 1'b1;
    buffer_full_rands[882]  = 1'b0;
    buffer_full_rands[883]  = 1'b1;
    buffer_full_rands[884]  = 1'b1;
    buffer_full_rands[885]  = 1'b1;
    buffer_full_rands[886]  = 1'b1;
    buffer_full_rands[887]  = 1'b1;
    buffer_full_rands[888]  = 1'b1;
    buffer_full_rands[889]  = 1'b0;
    buffer_full_rands[890]  = 1'b1;
    buffer_full_rands[891]  = 1'b0;
    buffer_full_rands[892]  = 1'b1;
    buffer_full_rands[893]  = 1'b0;
    buffer_full_rands[894]  = 1'b1;
    buffer_full_rands[895]  = 1'b0;
    buffer_full_rands[896]  = 1'b1;
    buffer_full_rands[897]  = 1'b0;
    buffer_full_rands[898]  = 1'b0;
    buffer_full_rands[899]  = 1'b1;
    buffer_full_rands[900]  = 1'b1;
    buffer_full_rands[901]  = 1'b0;
    buffer_full_rands[902]  = 1'b0;
    buffer_full_rands[903]  = 1'b1;
    buffer_full_rands[904]  = 1'b0;
    buffer_full_rands[905]  = 1'b1;
    buffer_full_rands[906]  = 1'b0;
    buffer_full_rands[907]  = 1'b1;
    buffer_full_rands[908]  = 1'b0;
    buffer_full_rands[909]  = 1'b0;
    buffer_full_rands[910]  = 1'b1;
    buffer_full_rands[911]  = 1'b0;
    buffer_full_rands[912]  = 1'b0;
    buffer_full_rands[913]  = 1'b1;
    buffer_full_rands[914]  = 1'b0;
    buffer_full_rands[915]  = 1'b0;
    buffer_full_rands[916]  = 1'b1;
    buffer_full_rands[917]  = 1'b0;
    buffer_full_rands[918]  = 1'b0;
    buffer_full_rands[919]  = 1'b1;
    buffer_full_rands[920]  = 1'b1;
    buffer_full_rands[921]  = 1'b1;
    buffer_full_rands[922]  = 1'b0;
    buffer_full_rands[923]  = 1'b0;
    buffer_full_rands[924]  = 1'b0;
    buffer_full_rands[925]  = 1'b0;
    buffer_full_rands[926]  = 1'b1;
    buffer_full_rands[927]  = 1'b0;
    buffer_full_rands[928]  = 1'b1;
    buffer_full_rands[929]  = 1'b0;
    buffer_full_rands[930]  = 1'b1;
    buffer_full_rands[931]  = 1'b0;
    buffer_full_rands[932]  = 1'b1;
    buffer_full_rands[933]  = 1'b0;
    buffer_full_rands[934]  = 1'b0;
    buffer_full_rands[935]  = 1'b0;
    buffer_full_rands[936]  = 1'b1;
    buffer_full_rands[937]  = 1'b1;
    buffer_full_rands[938]  = 1'b0;
    buffer_full_rands[939]  = 1'b1;
    buffer_full_rands[940]  = 1'b1;
    buffer_full_rands[941]  = 1'b1;
    buffer_full_rands[942]  = 1'b1;
    buffer_full_rands[943]  = 1'b0;
    buffer_full_rands[944]  = 1'b1;
    buffer_full_rands[945]  = 1'b1;
    buffer_full_rands[946]  = 1'b1;
    buffer_full_rands[947]  = 1'b1;
    buffer_full_rands[948]  = 1'b1;
    buffer_full_rands[949]  = 1'b1;
    buffer_full_rands[950]  = 1'b1;
    buffer_full_rands[951]  = 1'b1;
    buffer_full_rands[952]  = 1'b0;
    buffer_full_rands[953]  = 1'b0;
    buffer_full_rands[954]  = 1'b1;
    buffer_full_rands[955]  = 1'b0;
    buffer_full_rands[956]  = 1'b0;
    buffer_full_rands[957]  = 1'b0;
    buffer_full_rands[958]  = 1'b0;
    buffer_full_rands[959]  = 1'b1;
    buffer_full_rands[960]  = 1'b0;
    buffer_full_rands[961]  = 1'b0;
    buffer_full_rands[962]  = 1'b1;
    buffer_full_rands[963]  = 1'b0;
    buffer_full_rands[964]  = 1'b0;
    buffer_full_rands[965]  = 1'b1;
    buffer_full_rands[966]  = 1'b1;
    buffer_full_rands[967]  = 1'b0;
    buffer_full_rands[968]  = 1'b1;
    buffer_full_rands[969]  = 1'b0;
    buffer_full_rands[970]  = 1'b1;
    buffer_full_rands[971]  = 1'b0;
    buffer_full_rands[972]  = 1'b1;
    buffer_full_rands[973]  = 1'b0;
    buffer_full_rands[974]  = 1'b1;
    buffer_full_rands[975]  = 1'b0;
    buffer_full_rands[976]  = 1'b1;
    buffer_full_rands[977]  = 1'b1;
    buffer_full_rands[978]  = 1'b0;
    buffer_full_rands[979]  = 1'b0;
    buffer_full_rands[980]  = 1'b0;
    buffer_full_rands[981]  = 1'b0;
    buffer_full_rands[982]  = 1'b0;
    buffer_full_rands[983]  = 1'b0;
    buffer_full_rands[984]  = 1'b1;
    buffer_full_rands[985]  = 1'b1;
    buffer_full_rands[986]  = 1'b1;
    buffer_full_rands[987]  = 1'b1;
    buffer_full_rands[988]  = 1'b1;
    buffer_full_rands[989]  = 1'b0;
    buffer_full_rands[990]  = 1'b1;
    buffer_full_rands[991]  = 1'b0;
    buffer_full_rands[992]  = 1'b0;
    buffer_full_rands[993]  = 1'b1;
    buffer_full_rands[994]  = 1'b1;
    buffer_full_rands[995]  = 1'b0;
    buffer_full_rands[996]  = 1'b0;
    buffer_full_rands[997]  = 1'b1;
    buffer_full_rands[998]  = 1'b1;
    buffer_full_rands[999]  = 1'b1;
    //buffer_full_rands[1000] = 1'b0;

    stream_full_rands[0]    = 1'b0;
    stream_full_rands[1]    = 1'b0;
    stream_full_rands[2]    = 1'b0;
    stream_full_rands[3]    = 1'b0;
    stream_full_rands[4]    = 1'b0;
    stream_full_rands[5]    = 1'b1;
    stream_full_rands[6]    = 1'b0;
    stream_full_rands[7]    = 1'b0;
    stream_full_rands[8]    = 1'b1;
    stream_full_rands[9]    = 1'b0;
    stream_full_rands[10]   = 1'b0;
    stream_full_rands[11]   = 1'b1;
    stream_full_rands[12]   = 1'b0;
    stream_full_rands[13]   = 1'b1;
    stream_full_rands[14]   = 1'b1;
    stream_full_rands[15]   = 1'b0;
    stream_full_rands[16]   = 1'b0;
    stream_full_rands[17]   = 1'b1;
    stream_full_rands[18]   = 1'b0;
    stream_full_rands[19]   = 1'b1;
    stream_full_rands[20]   = 1'b0;
    stream_full_rands[21]   = 1'b1;
    stream_full_rands[22]   = 1'b0;
    stream_full_rands[23]   = 1'b0;
    stream_full_rands[24]   = 1'b0;
    stream_full_rands[25]   = 1'b1;
    stream_full_rands[26]   = 1'b0;
    stream_full_rands[27]   = 1'b0;
    stream_full_rands[28]   = 1'b1;
    stream_full_rands[29]   = 1'b1;
    stream_full_rands[30]   = 1'b1;
    stream_full_rands[31]   = 1'b1;
    stream_full_rands[32]   = 1'b1;
    stream_full_rands[33]   = 1'b1;
    stream_full_rands[34]   = 1'b1;
    stream_full_rands[35]   = 1'b1;
    stream_full_rands[36]   = 1'b0;
    stream_full_rands[37]   = 1'b1;
    stream_full_rands[38]   = 1'b0;
    stream_full_rands[39]   = 1'b1;
    stream_full_rands[40]   = 1'b1;
    stream_full_rands[41]   = 1'b1;
    stream_full_rands[42]   = 1'b1;
    stream_full_rands[43]   = 1'b1;
    stream_full_rands[44]   = 1'b0;
    stream_full_rands[45]   = 1'b1;
    stream_full_rands[46]   = 1'b0;
    stream_full_rands[47]   = 1'b0;
    stream_full_rands[48]   = 1'b0;
    stream_full_rands[49]   = 1'b1;
    stream_full_rands[50]   = 1'b0;
    stream_full_rands[51]   = 1'b0;
    stream_full_rands[52]   = 1'b1;
    stream_full_rands[53]   = 1'b0;
    stream_full_rands[54]   = 1'b1;
    stream_full_rands[55]   = 1'b0;
    stream_full_rands[56]   = 1'b0;
    stream_full_rands[57]   = 1'b1;
    stream_full_rands[58]   = 1'b0;
    stream_full_rands[59]   = 1'b0;
    stream_full_rands[60]   = 1'b1;
    stream_full_rands[61]   = 1'b1;
    stream_full_rands[62]   = 1'b1;
    stream_full_rands[63]   = 1'b1;
    stream_full_rands[64]   = 1'b1;
    stream_full_rands[65]   = 1'b0;
    stream_full_rands[66]   = 1'b1;
    stream_full_rands[67]   = 1'b0;
    stream_full_rands[68]   = 1'b1;
    stream_full_rands[69]   = 1'b1;
    stream_full_rands[70]   = 1'b1;
    stream_full_rands[71]   = 1'b1;
    stream_full_rands[72]   = 1'b0;
    stream_full_rands[73]   = 1'b0;
    stream_full_rands[74]   = 1'b0;
    stream_full_rands[75]   = 1'b1;
    stream_full_rands[76]   = 1'b0;
    stream_full_rands[77]   = 1'b1;
    stream_full_rands[78]   = 1'b0;
    stream_full_rands[79]   = 1'b0;
    stream_full_rands[80]   = 1'b0;
    stream_full_rands[81]   = 1'b0;
    stream_full_rands[82]   = 1'b0;
    stream_full_rands[83]   = 1'b1;
    stream_full_rands[84]   = 1'b1;
    stream_full_rands[85]   = 1'b1;
    stream_full_rands[86]   = 1'b0;
    stream_full_rands[87]   = 1'b0;
    stream_full_rands[88]   = 1'b0;
    stream_full_rands[89]   = 1'b1;
    stream_full_rands[90]   = 1'b1;
    stream_full_rands[91]   = 1'b1;
    stream_full_rands[92]   = 1'b0;
    stream_full_rands[93]   = 1'b1;
    stream_full_rands[94]   = 1'b1;
    stream_full_rands[95]   = 1'b1;
    stream_full_rands[96]   = 1'b0;
    stream_full_rands[97]   = 1'b1;
    stream_full_rands[98]   = 1'b0;
    stream_full_rands[99]   = 1'b0;
    stream_full_rands[100]  = 1'b1;
    stream_full_rands[101]  = 1'b0;
    stream_full_rands[102]  = 1'b0;
    stream_full_rands[103]  = 1'b1;
    stream_full_rands[104]  = 1'b1;
    stream_full_rands[105]  = 1'b0;
    stream_full_rands[106]  = 1'b0;
    stream_full_rands[107]  = 1'b0;
    stream_full_rands[108]  = 1'b1;
    stream_full_rands[109]  = 1'b0;
    stream_full_rands[110]  = 1'b1;
    stream_full_rands[111]  = 1'b0;
    stream_full_rands[112]  = 1'b1;
    stream_full_rands[113]  = 1'b1;
    stream_full_rands[114]  = 1'b0;
    stream_full_rands[115]  = 1'b1;
    stream_full_rands[116]  = 1'b0;
    stream_full_rands[117]  = 1'b1;
    stream_full_rands[118]  = 1'b1;
    stream_full_rands[119]  = 1'b1;
    stream_full_rands[120]  = 1'b0;
    stream_full_rands[121]  = 1'b0;
    stream_full_rands[122]  = 1'b0;
    stream_full_rands[123]  = 1'b1;
    stream_full_rands[124]  = 1'b0;
    stream_full_rands[125]  = 1'b0;
    stream_full_rands[126]  = 1'b0;
    stream_full_rands[127]  = 1'b0;
    stream_full_rands[128]  = 1'b0;
    stream_full_rands[129]  = 1'b0;
    stream_full_rands[130]  = 1'b1;
    stream_full_rands[131]  = 1'b1;
    stream_full_rands[132]  = 1'b0;
    stream_full_rands[133]  = 1'b0;
    stream_full_rands[134]  = 1'b0;
    stream_full_rands[135]  = 1'b1;
    stream_full_rands[136]  = 1'b1;
    stream_full_rands[137]  = 1'b1;
    stream_full_rands[138]  = 1'b0;
    stream_full_rands[139]  = 1'b0;
    stream_full_rands[140]  = 1'b0;
    stream_full_rands[141]  = 1'b1;
    stream_full_rands[142]  = 1'b1;
    stream_full_rands[143]  = 1'b1;
    stream_full_rands[144]  = 1'b1;
    stream_full_rands[145]  = 1'b1;
    stream_full_rands[146]  = 1'b0;
    stream_full_rands[147]  = 1'b1;
    stream_full_rands[148]  = 1'b0;
    stream_full_rands[149]  = 1'b1;
    stream_full_rands[150]  = 1'b1;
    stream_full_rands[151]  = 1'b1;
    stream_full_rands[152]  = 1'b0;
    stream_full_rands[153]  = 1'b0;
    stream_full_rands[154]  = 1'b1;
    stream_full_rands[155]  = 1'b1;
    stream_full_rands[156]  = 1'b1;
    stream_full_rands[157]  = 1'b1;
    stream_full_rands[158]  = 1'b0;
    stream_full_rands[159]  = 1'b1;
    stream_full_rands[160]  = 1'b1;
    stream_full_rands[161]  = 1'b1;
    stream_full_rands[162]  = 1'b0;
    stream_full_rands[163]  = 1'b1;
    stream_full_rands[164]  = 1'b1;
    stream_full_rands[165]  = 1'b1;
    stream_full_rands[166]  = 1'b0;
    stream_full_rands[167]  = 1'b1;
    stream_full_rands[168]  = 1'b0;
    stream_full_rands[169]  = 1'b1;
    stream_full_rands[170]  = 1'b1;
    stream_full_rands[171]  = 1'b0;
    stream_full_rands[172]  = 1'b1;
    stream_full_rands[173]  = 1'b0;
    stream_full_rands[174]  = 1'b1;
    stream_full_rands[175]  = 1'b0;
    stream_full_rands[176]  = 1'b0;
    stream_full_rands[177]  = 1'b0;
    stream_full_rands[178]  = 1'b0;
    stream_full_rands[179]  = 1'b1;
    stream_full_rands[180]  = 1'b0;
    stream_full_rands[181]  = 1'b0;
    stream_full_rands[182]  = 1'b0;
    stream_full_rands[183]  = 1'b0;
    stream_full_rands[184]  = 1'b0;
    stream_full_rands[185]  = 1'b0;
    stream_full_rands[186]  = 1'b0;
    stream_full_rands[187]  = 1'b1;
    stream_full_rands[188]  = 1'b1;
    stream_full_rands[189]  = 1'b1;
    stream_full_rands[190]  = 1'b1;
    stream_full_rands[191]  = 1'b1;
    stream_full_rands[192]  = 1'b1;
    stream_full_rands[193]  = 1'b0;
    stream_full_rands[194]  = 1'b0;
    stream_full_rands[195]  = 1'b0;
    stream_full_rands[196]  = 1'b1;
    stream_full_rands[197]  = 1'b1;
    stream_full_rands[198]  = 1'b0;
    stream_full_rands[199]  = 1'b1;
    stream_full_rands[200]  = 1'b1;
    stream_full_rands[201]  = 1'b0;
    stream_full_rands[202]  = 1'b1;
    stream_full_rands[203]  = 1'b0;
    stream_full_rands[204]  = 1'b0;
    stream_full_rands[205]  = 1'b0;
    stream_full_rands[206]  = 1'b0;
    stream_full_rands[207]  = 1'b1;
    stream_full_rands[208]  = 1'b1;
    stream_full_rands[209]  = 1'b0;
    stream_full_rands[210]  = 1'b1;
    stream_full_rands[211]  = 1'b1;
    stream_full_rands[212]  = 1'b1;
    stream_full_rands[213]  = 1'b0;
    stream_full_rands[214]  = 1'b1;
    stream_full_rands[215]  = 1'b1;
    stream_full_rands[216]  = 1'b1;
    stream_full_rands[217]  = 1'b1;
    stream_full_rands[218]  = 1'b1;
    stream_full_rands[219]  = 1'b1;
    stream_full_rands[220]  = 1'b0;
    stream_full_rands[221]  = 1'b1;
    stream_full_rands[222]  = 1'b1;
    stream_full_rands[223]  = 1'b0;
    stream_full_rands[224]  = 1'b0;
    stream_full_rands[225]  = 1'b1;
    stream_full_rands[226]  = 1'b0;
    stream_full_rands[227]  = 1'b0;
    stream_full_rands[228]  = 1'b0;
    stream_full_rands[229]  = 1'b1;
    stream_full_rands[230]  = 1'b0;
    stream_full_rands[231]  = 1'b1;
    stream_full_rands[232]  = 1'b1;
    stream_full_rands[233]  = 1'b0;
    stream_full_rands[234]  = 1'b0;
    stream_full_rands[235]  = 1'b0;
    stream_full_rands[236]  = 1'b1;
    stream_full_rands[237]  = 1'b1;
    stream_full_rands[238]  = 1'b1;
    stream_full_rands[239]  = 1'b0;
    stream_full_rands[240]  = 1'b1;
    stream_full_rands[241]  = 1'b0;
    stream_full_rands[242]  = 1'b0;
    stream_full_rands[243]  = 1'b0;
    stream_full_rands[244]  = 1'b0;
    stream_full_rands[245]  = 1'b0;
    stream_full_rands[246]  = 1'b1;
    stream_full_rands[247]  = 1'b0;
    stream_full_rands[248]  = 1'b0;
    stream_full_rands[249]  = 1'b1;
    stream_full_rands[250]  = 1'b0;
    stream_full_rands[251]  = 1'b0;
    stream_full_rands[252]  = 1'b1;
    stream_full_rands[253]  = 1'b1;
    stream_full_rands[254]  = 1'b0;
    stream_full_rands[255]  = 1'b1;
    stream_full_rands[256]  = 1'b0;
    stream_full_rands[257]  = 1'b1;
    stream_full_rands[258]  = 1'b0;
    stream_full_rands[259]  = 1'b0;
    stream_full_rands[260]  = 1'b1;
    stream_full_rands[261]  = 1'b1;
    stream_full_rands[262]  = 1'b1;
    stream_full_rands[263]  = 1'b1;
    stream_full_rands[264]  = 1'b1;
    stream_full_rands[265]  = 1'b0;
    stream_full_rands[266]  = 1'b0;
    stream_full_rands[267]  = 1'b0;
    stream_full_rands[268]  = 1'b0;
    stream_full_rands[269]  = 1'b1;
    stream_full_rands[270]  = 1'b1;
    stream_full_rands[271]  = 1'b1;
    stream_full_rands[272]  = 1'b0;
    stream_full_rands[273]  = 1'b0;
    stream_full_rands[274]  = 1'b1;
    stream_full_rands[275]  = 1'b0;
    stream_full_rands[276]  = 1'b1;
    stream_full_rands[277]  = 1'b1;
    stream_full_rands[278]  = 1'b0;
    stream_full_rands[279]  = 1'b0;
    stream_full_rands[280]  = 1'b1;
    stream_full_rands[281]  = 1'b0;
    stream_full_rands[282]  = 1'b1;
    stream_full_rands[283]  = 1'b0;
    stream_full_rands[284]  = 1'b0;
    stream_full_rands[285]  = 1'b0;
    stream_full_rands[286]  = 1'b0;
    stream_full_rands[287]  = 1'b0;
    stream_full_rands[288]  = 1'b0;
    stream_full_rands[289]  = 1'b0;
    stream_full_rands[290]  = 1'b1;
    stream_full_rands[291]  = 1'b0;
    stream_full_rands[292]  = 1'b1;
    stream_full_rands[293]  = 1'b0;
    stream_full_rands[294]  = 1'b0;
    stream_full_rands[295]  = 1'b1;
    stream_full_rands[296]  = 1'b0;
    stream_full_rands[297]  = 1'b1;
    stream_full_rands[298]  = 1'b0;
    stream_full_rands[299]  = 1'b0;
    stream_full_rands[300]  = 1'b1;
    stream_full_rands[301]  = 1'b0;
    stream_full_rands[302]  = 1'b1;
    stream_full_rands[303]  = 1'b1;
    stream_full_rands[304]  = 1'b1;
    stream_full_rands[305]  = 1'b1;
    stream_full_rands[306]  = 1'b1;
    stream_full_rands[307]  = 1'b1;
    stream_full_rands[308]  = 1'b0;
    stream_full_rands[309]  = 1'b1;
    stream_full_rands[310]  = 1'b1;
    stream_full_rands[311]  = 1'b0;
    stream_full_rands[312]  = 1'b0;
    stream_full_rands[313]  = 1'b1;
    stream_full_rands[314]  = 1'b0;
    stream_full_rands[315]  = 1'b1;
    stream_full_rands[316]  = 1'b1;
    stream_full_rands[317]  = 1'b1;
    stream_full_rands[318]  = 1'b0;
    stream_full_rands[319]  = 1'b0;
    stream_full_rands[320]  = 1'b0;
    stream_full_rands[321]  = 1'b0;
    stream_full_rands[322]  = 1'b0;
    stream_full_rands[323]  = 1'b1;
    stream_full_rands[324]  = 1'b1;
    stream_full_rands[325]  = 1'b0;
    stream_full_rands[326]  = 1'b1;
    stream_full_rands[327]  = 1'b0;
    stream_full_rands[328]  = 1'b0;
    stream_full_rands[329]  = 1'b0;
    stream_full_rands[330]  = 1'b0;
    stream_full_rands[331]  = 1'b1;
    stream_full_rands[332]  = 1'b1;
    stream_full_rands[333]  = 1'b0;
    stream_full_rands[334]  = 1'b1;
    stream_full_rands[335]  = 1'b0;
    stream_full_rands[336]  = 1'b0;
    stream_full_rands[337]  = 1'b1;
    stream_full_rands[338]  = 1'b0;
    stream_full_rands[339]  = 1'b0;
    stream_full_rands[340]  = 1'b0;
    stream_full_rands[341]  = 1'b1;
    stream_full_rands[342]  = 1'b1;
    stream_full_rands[343]  = 1'b1;
    stream_full_rands[344]  = 1'b0;
    stream_full_rands[345]  = 1'b1;
    stream_full_rands[346]  = 1'b0;
    stream_full_rands[347]  = 1'b1;
    stream_full_rands[348]  = 1'b0;
    stream_full_rands[349]  = 1'b1;
    stream_full_rands[350]  = 1'b0;
    stream_full_rands[351]  = 1'b1;
    stream_full_rands[352]  = 1'b0;
    stream_full_rands[353]  = 1'b0;
    stream_full_rands[354]  = 1'b0;
    stream_full_rands[355]  = 1'b0;
    stream_full_rands[356]  = 1'b1;
    stream_full_rands[357]  = 1'b1;
    stream_full_rands[358]  = 1'b1;
    stream_full_rands[359]  = 1'b0;
    stream_full_rands[360]  = 1'b1;
    stream_full_rands[361]  = 1'b1;
    stream_full_rands[362]  = 1'b0;
    stream_full_rands[363]  = 1'b1;
    stream_full_rands[364]  = 1'b0;
    stream_full_rands[365]  = 1'b0;
    stream_full_rands[366]  = 1'b1;
    stream_full_rands[367]  = 1'b0;
    stream_full_rands[368]  = 1'b0;
    stream_full_rands[369]  = 1'b0;
    stream_full_rands[370]  = 1'b1;
    stream_full_rands[371]  = 1'b1;
    stream_full_rands[372]  = 1'b0;
    stream_full_rands[373]  = 1'b1;
    stream_full_rands[374]  = 1'b1;
    stream_full_rands[375]  = 1'b1;
    stream_full_rands[376]  = 1'b0;
    stream_full_rands[377]  = 1'b1;
    stream_full_rands[378]  = 1'b0;
    stream_full_rands[379]  = 1'b1;
    stream_full_rands[380]  = 1'b1;
    stream_full_rands[381]  = 1'b0;
    stream_full_rands[382]  = 1'b0;
    stream_full_rands[383]  = 1'b0;
    stream_full_rands[384]  = 1'b0;
    stream_full_rands[385]  = 1'b1;
    stream_full_rands[386]  = 1'b0;
    stream_full_rands[387]  = 1'b1;
    stream_full_rands[388]  = 1'b1;
    stream_full_rands[389]  = 1'b1;
    stream_full_rands[390]  = 1'b0;
    stream_full_rands[391]  = 1'b0;
    stream_full_rands[392]  = 1'b0;
    stream_full_rands[393]  = 1'b1;
    stream_full_rands[394]  = 1'b1;
    stream_full_rands[395]  = 1'b0;
    stream_full_rands[396]  = 1'b0;
    stream_full_rands[397]  = 1'b0;
    stream_full_rands[398]  = 1'b1;
    stream_full_rands[399]  = 1'b1;
    stream_full_rands[400]  = 1'b1;
    stream_full_rands[401]  = 1'b0;
    stream_full_rands[402]  = 1'b0;
    stream_full_rands[403]  = 1'b0;
    stream_full_rands[404]  = 1'b1;
    stream_full_rands[405]  = 1'b1;
    stream_full_rands[406]  = 1'b0;
    stream_full_rands[407]  = 1'b1;
    stream_full_rands[408]  = 1'b1;
    stream_full_rands[409]  = 1'b1;
    stream_full_rands[410]  = 1'b1;
    stream_full_rands[411]  = 1'b0;
    stream_full_rands[412]  = 1'b1;
    stream_full_rands[413]  = 1'b0;
    stream_full_rands[414]  = 1'b1;
    stream_full_rands[415]  = 1'b1;
    stream_full_rands[416]  = 1'b0;
    stream_full_rands[417]  = 1'b1;
    stream_full_rands[418]  = 1'b0;
    stream_full_rands[419]  = 1'b0;
    stream_full_rands[420]  = 1'b1;
    stream_full_rands[421]  = 1'b0;
    stream_full_rands[422]  = 1'b0;
    stream_full_rands[423]  = 1'b0;
    stream_full_rands[424]  = 1'b1;
    stream_full_rands[425]  = 1'b0;
    stream_full_rands[426]  = 1'b0;
    stream_full_rands[427]  = 1'b1;
    stream_full_rands[428]  = 1'b0;
    stream_full_rands[429]  = 1'b0;
    stream_full_rands[430]  = 1'b1;
    stream_full_rands[431]  = 1'b0;
    stream_full_rands[432]  = 1'b1;
    stream_full_rands[433]  = 1'b1;
    stream_full_rands[434]  = 1'b0;
    stream_full_rands[435]  = 1'b1;
    stream_full_rands[436]  = 1'b0;
    stream_full_rands[437]  = 1'b0;
    stream_full_rands[438]  = 1'b1;
    stream_full_rands[439]  = 1'b1;
    stream_full_rands[440]  = 1'b1;
    stream_full_rands[441]  = 1'b0;
    stream_full_rands[442]  = 1'b1;
    stream_full_rands[443]  = 1'b1;
    stream_full_rands[444]  = 1'b0;
    stream_full_rands[445]  = 1'b0;
    stream_full_rands[446]  = 1'b1;
    stream_full_rands[447]  = 1'b0;
    stream_full_rands[448]  = 1'b1;
    stream_full_rands[449]  = 1'b1;
    stream_full_rands[450]  = 1'b0;
    stream_full_rands[451]  = 1'b1;
    stream_full_rands[452]  = 1'b1;
    stream_full_rands[453]  = 1'b1;
    stream_full_rands[454]  = 1'b1;
    stream_full_rands[455]  = 1'b1;
    stream_full_rands[456]  = 1'b1;
    stream_full_rands[457]  = 1'b0;
    stream_full_rands[458]  = 1'b0;
    stream_full_rands[459]  = 1'b0;
    stream_full_rands[460]  = 1'b1;
    stream_full_rands[461]  = 1'b0;
    stream_full_rands[462]  = 1'b1;
    stream_full_rands[463]  = 1'b1;
    stream_full_rands[464]  = 1'b1;
    stream_full_rands[465]  = 1'b0;
    stream_full_rands[466]  = 1'b1;
    stream_full_rands[467]  = 1'b1;
    stream_full_rands[468]  = 1'b1;
    stream_full_rands[469]  = 1'b0;
    stream_full_rands[470]  = 1'b0;
    stream_full_rands[471]  = 1'b1;
    stream_full_rands[472]  = 1'b1;
    stream_full_rands[473]  = 1'b0;
    stream_full_rands[474]  = 1'b1;
    stream_full_rands[475]  = 1'b1;
    stream_full_rands[476]  = 1'b0;
    stream_full_rands[477]  = 1'b1;
    stream_full_rands[478]  = 1'b1;
    stream_full_rands[479]  = 1'b0;
    stream_full_rands[480]  = 1'b0;
    stream_full_rands[481]  = 1'b0;
    stream_full_rands[482]  = 1'b1;
    stream_full_rands[483]  = 1'b0;
    stream_full_rands[484]  = 1'b1;
    stream_full_rands[485]  = 1'b0;
    stream_full_rands[486]  = 1'b1;
    stream_full_rands[487]  = 1'b0;
    stream_full_rands[488]  = 1'b1;
    stream_full_rands[489]  = 1'b1;
    stream_full_rands[490]  = 1'b0;
    stream_full_rands[491]  = 1'b1;
    stream_full_rands[492]  = 1'b0;
    stream_full_rands[493]  = 1'b0;
    stream_full_rands[494]  = 1'b0;
    stream_full_rands[495]  = 1'b1;
    stream_full_rands[496]  = 1'b1;
    stream_full_rands[497]  = 1'b0;
    stream_full_rands[498]  = 1'b0;
    stream_full_rands[499]  = 1'b0;
    stream_full_rands[500]  = 1'b0;
    stream_full_rands[501]  = 1'b0;
    stream_full_rands[502]  = 1'b0;
    stream_full_rands[503]  = 1'b0;
    stream_full_rands[504]  = 1'b1;
    stream_full_rands[505]  = 1'b0;
    stream_full_rands[506]  = 1'b1;
    stream_full_rands[507]  = 1'b1;
    stream_full_rands[508]  = 1'b0;
    stream_full_rands[509]  = 1'b1;
    stream_full_rands[510]  = 1'b0;
    stream_full_rands[511]  = 1'b1;
    stream_full_rands[512]  = 1'b1;
    stream_full_rands[513]  = 1'b0;
    stream_full_rands[514]  = 1'b0;
    stream_full_rands[515]  = 1'b1;
    stream_full_rands[516]  = 1'b0;
    stream_full_rands[517]  = 1'b1;
    stream_full_rands[518]  = 1'b1;
    stream_full_rands[519]  = 1'b1;
    stream_full_rands[520]  = 1'b0;
    stream_full_rands[521]  = 1'b0;
    stream_full_rands[522]  = 1'b0;
    stream_full_rands[523]  = 1'b1;
    stream_full_rands[524]  = 1'b1;
    stream_full_rands[525]  = 1'b0;
    stream_full_rands[526]  = 1'b1;
    stream_full_rands[527]  = 1'b1;
    stream_full_rands[528]  = 1'b1;
    stream_full_rands[529]  = 1'b0;
    stream_full_rands[530]  = 1'b0;
    stream_full_rands[531]  = 1'b0;
    stream_full_rands[532]  = 1'b1;
    stream_full_rands[533]  = 1'b0;
    stream_full_rands[534]  = 1'b0;
    stream_full_rands[535]  = 1'b0;
    stream_full_rands[536]  = 1'b0;
    stream_full_rands[537]  = 1'b1;
    stream_full_rands[538]  = 1'b0;
    stream_full_rands[539]  = 1'b0;
    stream_full_rands[540]  = 1'b0;
    stream_full_rands[541]  = 1'b0;
    stream_full_rands[542]  = 1'b1;
    stream_full_rands[543]  = 1'b0;
    stream_full_rands[544]  = 1'b1;
    stream_full_rands[545]  = 1'b1;
    stream_full_rands[546]  = 1'b0;
    stream_full_rands[547]  = 1'b1;
    stream_full_rands[548]  = 1'b0;
    stream_full_rands[549]  = 1'b0;
    stream_full_rands[550]  = 1'b0;
    stream_full_rands[551]  = 1'b1;
    stream_full_rands[552]  = 1'b0;
    stream_full_rands[553]  = 1'b0;
    stream_full_rands[554]  = 1'b0;
    stream_full_rands[555]  = 1'b1;
    stream_full_rands[556]  = 1'b0;
    stream_full_rands[557]  = 1'b1;
    stream_full_rands[558]  = 1'b0;
    stream_full_rands[559]  = 1'b1;
    stream_full_rands[560]  = 1'b1;
    stream_full_rands[561]  = 1'b0;
    stream_full_rands[562]  = 1'b0;
    stream_full_rands[563]  = 1'b0;
    stream_full_rands[564]  = 1'b1;
    stream_full_rands[565]  = 1'b1;
    stream_full_rands[566]  = 1'b0;
    stream_full_rands[567]  = 1'b0;
    stream_full_rands[568]  = 1'b0;
    stream_full_rands[569]  = 1'b1;
    stream_full_rands[570]  = 1'b0;
    stream_full_rands[571]  = 1'b1;
    stream_full_rands[572]  = 1'b1;
    stream_full_rands[573]  = 1'b1;
    stream_full_rands[574]  = 1'b0;
    stream_full_rands[575]  = 1'b1;
    stream_full_rands[576]  = 1'b1;
    stream_full_rands[577]  = 1'b0;
    stream_full_rands[578]  = 1'b0;
    stream_full_rands[579]  = 1'b1;
    stream_full_rands[580]  = 1'b0;
    stream_full_rands[581]  = 1'b1;
    stream_full_rands[582]  = 1'b1;
    stream_full_rands[583]  = 1'b0;
    stream_full_rands[584]  = 1'b1;
    stream_full_rands[585]  = 1'b1;
    stream_full_rands[586]  = 1'b1;
    stream_full_rands[587]  = 1'b0;
    stream_full_rands[588]  = 1'b1;
    stream_full_rands[589]  = 1'b0;
    stream_full_rands[590]  = 1'b1;
    stream_full_rands[591]  = 1'b1;
    stream_full_rands[592]  = 1'b0;
    stream_full_rands[593]  = 1'b0;
    stream_full_rands[594]  = 1'b1;
    stream_full_rands[595]  = 1'b1;
    stream_full_rands[596]  = 1'b0;
    stream_full_rands[597]  = 1'b0;
    stream_full_rands[598]  = 1'b1;
    stream_full_rands[599]  = 1'b1;
    stream_full_rands[600]  = 1'b1;
    stream_full_rands[601]  = 1'b0;
    stream_full_rands[602]  = 1'b1;
    stream_full_rands[603]  = 1'b0;
    stream_full_rands[604]  = 1'b0;
    stream_full_rands[605]  = 1'b1;
    stream_full_rands[606]  = 1'b0;
    stream_full_rands[607]  = 1'b0;
    stream_full_rands[608]  = 1'b1;
    stream_full_rands[609]  = 1'b1;
    stream_full_rands[610]  = 1'b0;
    stream_full_rands[611]  = 1'b1;
    stream_full_rands[612]  = 1'b0;
    stream_full_rands[613]  = 1'b0;
    stream_full_rands[614]  = 1'b0;
    stream_full_rands[615]  = 1'b1;
    stream_full_rands[616]  = 1'b0;
    stream_full_rands[617]  = 1'b0;
    stream_full_rands[618]  = 1'b1;
    stream_full_rands[619]  = 1'b1;
    stream_full_rands[620]  = 1'b1;
    stream_full_rands[621]  = 1'b1;
    stream_full_rands[622]  = 1'b0;
    stream_full_rands[623]  = 1'b1;
    stream_full_rands[624]  = 1'b1;
    stream_full_rands[625]  = 1'b0;
    stream_full_rands[626]  = 1'b1;
    stream_full_rands[627]  = 1'b0;
    stream_full_rands[628]  = 1'b0;
    stream_full_rands[629]  = 1'b1;
    stream_full_rands[630]  = 1'b1;
    stream_full_rands[631]  = 1'b0;
    stream_full_rands[632]  = 1'b1;
    stream_full_rands[633]  = 1'b0;
    stream_full_rands[634]  = 1'b1;
    stream_full_rands[635]  = 1'b0;
    stream_full_rands[636]  = 1'b0;
    stream_full_rands[637]  = 1'b0;
    stream_full_rands[638]  = 1'b0;
    stream_full_rands[639]  = 1'b1;
    stream_full_rands[640]  = 1'b1;
    stream_full_rands[641]  = 1'b0;
    stream_full_rands[642]  = 1'b0;
    stream_full_rands[643]  = 1'b0;
    stream_full_rands[644]  = 1'b1;
    stream_full_rands[645]  = 1'b0;
    stream_full_rands[646]  = 1'b1;
    stream_full_rands[647]  = 1'b0;
    stream_full_rands[648]  = 1'b1;
    stream_full_rands[649]  = 1'b0;
    stream_full_rands[650]  = 1'b1;
    stream_full_rands[651]  = 1'b1;
    stream_full_rands[652]  = 1'b1;
    stream_full_rands[653]  = 1'b1;
    stream_full_rands[654]  = 1'b0;
    stream_full_rands[655]  = 1'b0;
    stream_full_rands[656]  = 1'b1;
    stream_full_rands[657]  = 1'b1;
    stream_full_rands[658]  = 1'b1;
    stream_full_rands[659]  = 1'b1;
    stream_full_rands[660]  = 1'b1;
    stream_full_rands[661]  = 1'b0;
    stream_full_rands[662]  = 1'b1;
    stream_full_rands[663]  = 1'b0;
    stream_full_rands[664]  = 1'b1;
    stream_full_rands[665]  = 1'b1;
    stream_full_rands[666]  = 1'b0;
    stream_full_rands[667]  = 1'b0;
    stream_full_rands[668]  = 1'b1;
    stream_full_rands[669]  = 1'b0;
    stream_full_rands[670]  = 1'b0;
    stream_full_rands[671]  = 1'b1;
    stream_full_rands[672]  = 1'b1;
    stream_full_rands[673]  = 1'b1;
    stream_full_rands[674]  = 1'b1;
    stream_full_rands[675]  = 1'b1;
    stream_full_rands[676]  = 1'b0;
    stream_full_rands[677]  = 1'b1;
    stream_full_rands[678]  = 1'b1;
    stream_full_rands[679]  = 1'b1;
    stream_full_rands[680]  = 1'b0;
    stream_full_rands[681]  = 1'b0;
    stream_full_rands[682]  = 1'b0;
    stream_full_rands[683]  = 1'b0;
    stream_full_rands[684]  = 1'b1;
    stream_full_rands[685]  = 1'b0;
    stream_full_rands[686]  = 1'b0;
    stream_full_rands[687]  = 1'b1;
    stream_full_rands[688]  = 1'b0;
    stream_full_rands[689]  = 1'b0;
    stream_full_rands[690]  = 1'b1;
    stream_full_rands[691]  = 1'b0;
    stream_full_rands[692]  = 1'b1;
    stream_full_rands[693]  = 1'b1;
    stream_full_rands[694]  = 1'b0;
    stream_full_rands[695]  = 1'b1;
    stream_full_rands[696]  = 1'b0;
    stream_full_rands[697]  = 1'b1;
    stream_full_rands[698]  = 1'b1;
    stream_full_rands[699]  = 1'b0;
    stream_full_rands[700]  = 1'b0;
    stream_full_rands[701]  = 1'b1;
    stream_full_rands[702]  = 1'b0;
    stream_full_rands[703]  = 1'b0;
    stream_full_rands[704]  = 1'b1;
    stream_full_rands[705]  = 1'b1;
    stream_full_rands[706]  = 1'b0;
    stream_full_rands[707]  = 1'b0;
    stream_full_rands[708]  = 1'b0;
    stream_full_rands[709]  = 1'b1;
    stream_full_rands[710]  = 1'b1;
    stream_full_rands[711]  = 1'b0;
    stream_full_rands[712]  = 1'b1;
    stream_full_rands[713]  = 1'b0;
    stream_full_rands[714]  = 1'b1;
    stream_full_rands[715]  = 1'b0;
    stream_full_rands[716]  = 1'b0;
    stream_full_rands[717]  = 1'b1;
    stream_full_rands[718]  = 1'b0;
    stream_full_rands[719]  = 1'b1;
    stream_full_rands[720]  = 1'b1;
    stream_full_rands[721]  = 1'b1;
    stream_full_rands[722]  = 1'b0;
    stream_full_rands[723]  = 1'b0;
    stream_full_rands[724]  = 1'b0;
    stream_full_rands[725]  = 1'b0;
    stream_full_rands[726]  = 1'b1;
    stream_full_rands[727]  = 1'b0;
    stream_full_rands[728]  = 1'b1;
    stream_full_rands[729]  = 1'b1;
    stream_full_rands[730]  = 1'b1;
    stream_full_rands[731]  = 1'b1;
    stream_full_rands[732]  = 1'b0;
    stream_full_rands[733]  = 1'b0;
    stream_full_rands[734]  = 1'b0;
    stream_full_rands[735]  = 1'b1;
    stream_full_rands[736]  = 1'b0;
    stream_full_rands[737]  = 1'b1;
    stream_full_rands[738]  = 1'b1;
    stream_full_rands[739]  = 1'b1;
    stream_full_rands[740]  = 1'b0;
    stream_full_rands[741]  = 1'b0;
    stream_full_rands[742]  = 1'b0;
    stream_full_rands[743]  = 1'b1;
    stream_full_rands[744]  = 1'b0;
    stream_full_rands[745]  = 1'b0;
    stream_full_rands[746]  = 1'b0;
    stream_full_rands[747]  = 1'b0;
    stream_full_rands[748]  = 1'b1;
    stream_full_rands[749]  = 1'b0;
    stream_full_rands[750]  = 1'b0;
    stream_full_rands[751]  = 1'b0;
    stream_full_rands[752]  = 1'b1;
    stream_full_rands[753]  = 1'b0;
    stream_full_rands[754]  = 1'b1;
    stream_full_rands[755]  = 1'b0;
    stream_full_rands[756]  = 1'b1;
    stream_full_rands[757]  = 1'b1;
    stream_full_rands[758]  = 1'b1;
    stream_full_rands[759]  = 1'b1;
    stream_full_rands[760]  = 1'b0;
    stream_full_rands[761]  = 1'b1;
    stream_full_rands[762]  = 1'b1;
    stream_full_rands[763]  = 1'b0;
    stream_full_rands[764]  = 1'b0;
    stream_full_rands[765]  = 1'b1;
    stream_full_rands[766]  = 1'b1;
    stream_full_rands[767]  = 1'b0;
    stream_full_rands[768]  = 1'b0;
    stream_full_rands[769]  = 1'b1;
    stream_full_rands[770]  = 1'b0;
    stream_full_rands[771]  = 1'b1;
    stream_full_rands[772]  = 1'b0;
    stream_full_rands[773]  = 1'b1;
    stream_full_rands[774]  = 1'b1;
    stream_full_rands[775]  = 1'b1;
    stream_full_rands[776]  = 1'b1;
    stream_full_rands[777]  = 1'b0;
    stream_full_rands[778]  = 1'b0;
    stream_full_rands[779]  = 1'b0;
    stream_full_rands[780]  = 1'b1;
    stream_full_rands[781]  = 1'b1;
    stream_full_rands[782]  = 1'b0;
    stream_full_rands[783]  = 1'b0;
    stream_full_rands[784]  = 1'b0;
    stream_full_rands[785]  = 1'b0;
    stream_full_rands[786]  = 1'b0;
    stream_full_rands[787]  = 1'b1;
    stream_full_rands[788]  = 1'b0;
    stream_full_rands[789]  = 1'b1;
    stream_full_rands[790]  = 1'b1;
    stream_full_rands[791]  = 1'b0;
    stream_full_rands[792]  = 1'b0;
    stream_full_rands[793]  = 1'b0;
    stream_full_rands[794]  = 1'b1;
    stream_full_rands[795]  = 1'b1;
    stream_full_rands[796]  = 1'b1;
    stream_full_rands[797]  = 1'b1;
    stream_full_rands[798]  = 1'b0;
    stream_full_rands[799]  = 1'b1;
    stream_full_rands[800]  = 1'b1;
    stream_full_rands[801]  = 1'b0;
    stream_full_rands[802]  = 1'b1;
    stream_full_rands[803]  = 1'b0;
    stream_full_rands[804]  = 1'b0;
    stream_full_rands[805]  = 1'b1;
    stream_full_rands[806]  = 1'b1;
    stream_full_rands[807]  = 1'b1;
    stream_full_rands[808]  = 1'b1;
    stream_full_rands[809]  = 1'b1;
    stream_full_rands[810]  = 1'b1;
    stream_full_rands[811]  = 1'b1;
    stream_full_rands[812]  = 1'b1;
    stream_full_rands[813]  = 1'b1;
    stream_full_rands[814]  = 1'b0;
    stream_full_rands[815]  = 1'b0;
    stream_full_rands[816]  = 1'b0;
    stream_full_rands[817]  = 1'b1;
    stream_full_rands[818]  = 1'b1;
    stream_full_rands[819]  = 1'b1;
    stream_full_rands[820]  = 1'b1;
    stream_full_rands[821]  = 1'b0;
    stream_full_rands[822]  = 1'b1;
    stream_full_rands[823]  = 1'b1;
    stream_full_rands[824]  = 1'b1;
    stream_full_rands[825]  = 1'b1;
    stream_full_rands[826]  = 1'b0;
    stream_full_rands[827]  = 1'b0;
    stream_full_rands[828]  = 1'b1;
    stream_full_rands[829]  = 1'b0;
    stream_full_rands[830]  = 1'b0;
    stream_full_rands[831]  = 1'b1;
    stream_full_rands[832]  = 1'b0;
    stream_full_rands[833]  = 1'b0;
    stream_full_rands[834]  = 1'b0;
    stream_full_rands[835]  = 1'b0;
    stream_full_rands[836]  = 1'b1;
    stream_full_rands[837]  = 1'b1;
    stream_full_rands[838]  = 1'b0;
    stream_full_rands[839]  = 1'b0;
    stream_full_rands[840]  = 1'b0;
    stream_full_rands[841]  = 1'b1;
    stream_full_rands[842]  = 1'b1;
    stream_full_rands[843]  = 1'b1;
    stream_full_rands[844]  = 1'b1;
    stream_full_rands[845]  = 1'b0;
    stream_full_rands[846]  = 1'b0;
    stream_full_rands[847]  = 1'b0;
    stream_full_rands[848]  = 1'b0;
    stream_full_rands[849]  = 1'b0;
    stream_full_rands[850]  = 1'b1;
    stream_full_rands[851]  = 1'b1;
    stream_full_rands[852]  = 1'b0;
    stream_full_rands[853]  = 1'b1;
    stream_full_rands[854]  = 1'b0;
    stream_full_rands[855]  = 1'b0;
    stream_full_rands[856]  = 1'b0;
    stream_full_rands[857]  = 1'b1;
    stream_full_rands[858]  = 1'b1;
    stream_full_rands[859]  = 1'b0;
    stream_full_rands[860]  = 1'b0;
    stream_full_rands[861]  = 1'b0;
    stream_full_rands[862]  = 1'b1;
    stream_full_rands[863]  = 1'b1;
    stream_full_rands[864]  = 1'b0;
    stream_full_rands[865]  = 1'b0;
    stream_full_rands[866]  = 1'b1;
    stream_full_rands[867]  = 1'b0;
    stream_full_rands[868]  = 1'b1;
    stream_full_rands[869]  = 1'b0;
    stream_full_rands[870]  = 1'b1;
    stream_full_rands[871]  = 1'b0;
    stream_full_rands[872]  = 1'b1;
    stream_full_rands[873]  = 1'b0;
    stream_full_rands[874]  = 1'b1;
    stream_full_rands[875]  = 1'b1;
    stream_full_rands[876]  = 1'b0;
    stream_full_rands[877]  = 1'b0;
    stream_full_rands[878]  = 1'b1;
    stream_full_rands[879]  = 1'b0;
    stream_full_rands[880]  = 1'b0;
    stream_full_rands[881]  = 1'b0;
    stream_full_rands[882]  = 1'b0;
    stream_full_rands[883]  = 1'b1;
    stream_full_rands[884]  = 1'b1;
    stream_full_rands[885]  = 1'b0;
    stream_full_rands[886]  = 1'b1;
    stream_full_rands[887]  = 1'b1;
    stream_full_rands[888]  = 1'b1;
    stream_full_rands[889]  = 1'b0;
    stream_full_rands[890]  = 1'b1;
    stream_full_rands[891]  = 1'b1;
    stream_full_rands[892]  = 1'b1;
    stream_full_rands[893]  = 1'b1;
    stream_full_rands[894]  = 1'b0;
    stream_full_rands[895]  = 1'b1;
    stream_full_rands[896]  = 1'b0;
    stream_full_rands[897]  = 1'b1;
    stream_full_rands[898]  = 1'b1;
    stream_full_rands[899]  = 1'b0;
    stream_full_rands[900]  = 1'b0;
    stream_full_rands[901]  = 1'b1;
    stream_full_rands[902]  = 1'b0;
    stream_full_rands[903]  = 1'b1;
    stream_full_rands[904]  = 1'b1;
    stream_full_rands[905]  = 1'b0;
    stream_full_rands[906]  = 1'b0;
    stream_full_rands[907]  = 1'b0;
    stream_full_rands[908]  = 1'b1;
    stream_full_rands[909]  = 1'b0;
    stream_full_rands[910]  = 1'b0;
    stream_full_rands[911]  = 1'b0;
    stream_full_rands[912]  = 1'b1;
    stream_full_rands[913]  = 1'b0;
    stream_full_rands[914]  = 1'b1;
    stream_full_rands[915]  = 1'b1;
    stream_full_rands[916]  = 1'b1;
    stream_full_rands[917]  = 1'b0;
    stream_full_rands[918]  = 1'b0;
    stream_full_rands[919]  = 1'b0;
    stream_full_rands[920]  = 1'b0;
    stream_full_rands[921]  = 1'b0;
    stream_full_rands[922]  = 1'b1;
    stream_full_rands[923]  = 1'b1;
    stream_full_rands[924]  = 1'b0;
    stream_full_rands[925]  = 1'b0;
    stream_full_rands[926]  = 1'b0;
    stream_full_rands[927]  = 1'b1;
    stream_full_rands[928]  = 1'b1;
    stream_full_rands[929]  = 1'b0;
    stream_full_rands[930]  = 1'b1;
    stream_full_rands[931]  = 1'b0;
    stream_full_rands[932]  = 1'b0;
    stream_full_rands[933]  = 1'b0;
    stream_full_rands[934]  = 1'b0;
    stream_full_rands[935]  = 1'b0;
    stream_full_rands[936]  = 1'b1;
    stream_full_rands[937]  = 1'b0;
    stream_full_rands[938]  = 1'b1;
    stream_full_rands[939]  = 1'b0;
    stream_full_rands[940]  = 1'b1;
    stream_full_rands[941]  = 1'b1;
    stream_full_rands[942]  = 1'b1;
    stream_full_rands[943]  = 1'b1;
    stream_full_rands[944]  = 1'b1;
    stream_full_rands[945]  = 1'b0;
    stream_full_rands[946]  = 1'b1;
    stream_full_rands[947]  = 1'b0;
    stream_full_rands[948]  = 1'b0;
    stream_full_rands[949]  = 1'b0;
    stream_full_rands[950]  = 1'b1;
    stream_full_rands[951]  = 1'b1;
    stream_full_rands[952]  = 1'b1;
    stream_full_rands[953]  = 1'b1;
    stream_full_rands[954]  = 1'b1;
    stream_full_rands[955]  = 1'b0;
    stream_full_rands[956]  = 1'b0;
    stream_full_rands[957]  = 1'b0;
    stream_full_rands[958]  = 1'b1;
    stream_full_rands[959]  = 1'b0;
    stream_full_rands[960]  = 1'b1;
    stream_full_rands[961]  = 1'b0;
    stream_full_rands[962]  = 1'b1;
    stream_full_rands[963]  = 1'b0;
    stream_full_rands[964]  = 1'b0;
    stream_full_rands[965]  = 1'b1;
    stream_full_rands[966]  = 1'b1;
    stream_full_rands[967]  = 1'b0;
    stream_full_rands[968]  = 1'b0;
    stream_full_rands[969]  = 1'b0;
    stream_full_rands[970]  = 1'b0;
    stream_full_rands[971]  = 1'b1;
    stream_full_rands[972]  = 1'b0;
    stream_full_rands[973]  = 1'b0;
    stream_full_rands[974]  = 1'b0;
    stream_full_rands[975]  = 1'b1;
    stream_full_rands[976]  = 1'b1;
    stream_full_rands[977]  = 1'b1;
    stream_full_rands[978]  = 1'b0;
    stream_full_rands[979]  = 1'b1;
    stream_full_rands[980]  = 1'b0;
    stream_full_rands[981]  = 1'b1;
    stream_full_rands[982]  = 1'b1;
    stream_full_rands[983]  = 1'b0;
    stream_full_rands[984]  = 1'b1;
    stream_full_rands[985]  = 1'b1;
    stream_full_rands[986]  = 1'b1;
    stream_full_rands[987]  = 1'b1;
    stream_full_rands[988]  = 1'b1;
    stream_full_rands[989]  = 1'b1;
    stream_full_rands[990]  = 1'b0;
    stream_full_rands[991]  = 1'b0;
    stream_full_rands[992]  = 1'b0;
    stream_full_rands[993]  = 1'b1;
    stream_full_rands[994]  = 1'b0;
    stream_full_rands[995]  = 1'b0;
    stream_full_rands[996]  = 1'b0;
    stream_full_rands[997]  = 1'b1;
    stream_full_rands[998]  = 1'b1;
    stream_full_rands[999]  = 1'b1;
    //stream_full_rands[1000] = 1'b1;
  end // initial begin

  always @(posedge clk) begin // @(negedge clk) begin
    ctr <= ctr + 1;

    pass <= 0;
    fail <= 0;

    if (reset) begin
      ctr <= 0;
      state <= start;
      counts_equal <= 0;
      counts_equal_ctr <= 0;

      
    end else begin
      size_idx <= (size_idx + 1) % RANDS;
      pu_id_idx <= (pu_id_idx + 1) % RANDS;
      d_type_idx <= (d_type_idx + 1) % RANDS;

      inbuf_empty_idx <= (inbuf_empty_idx + 1) % RANDS;
      buffer_full_idx <= (buffer_full_idx + 1) % RANDS;
      stream_full_idx <= (stream_full_idx + 1) % RANDS;

      case(state)
        idle : begin
          // don't do anything here
        end

        // Initialize all the relevant values
        start : begin          
          rd_req <= 0;
          rd_req_size <= 0;
          rd_req_pu_id <= 0;
          rd_req_d_type <= 0;
          d_0_count <= 0;
          d_1_count <= 0;
          rd_pointer <= 0;
          read_info_pop_count <= 0;
          d0_pop_count <= 0;
          d1_pop_count <= 0;
          read_count <= 0;
          reqs_sent <= 0;

          size_idx <= 0;
          pu_id_idx <= 0;
          d_type_idx <= 0;
          inbuf_empty_idx <= 0;
          buffer_full_idx <= 0;
          stream_full_idx <= 0;

          ctr <= 0;
          state <= send_reqs_init;
          counts_equal <= 0;
          counts_equal_ctr <= 0;
        end
  
        send_reqs_init : begin
          if (read_info_full) begin
            // wait here until it's not full
            reqs_sent <= reqs_sent;
          end else if (reqs_sent < TESTCASES) begin
            //$display("State: send_reqs_init. Reqs_sent <= %d\n", reqs_sent);

            
            rd_req <= 1;
            rd_req_size <= rd_req_size_urands[size_idx];
            rd_req_pu_id <= rd_req_pu_id_urands[pu_id_idx];
            rd_req_d_type <= rd_req_d_type_urands[d_type_idx];

            read_count <= read_count + rd_req_size;
            //$display ("Requesting %d reads of type %d", rd_req_size, rd_req_d_type);
            if (rd_req_d_type == 0)
              d_0_count <= d_0_count + rd_req_size;
            else
              d_1_count <= d_1_count + rd_req_size;

            ctr <= 0;
            state <= send_reqs_complete;

          end else begin // if (reqs_sent < 1000)
            //$display("State: send_reqs_init going to finish. Reqs_sent <= %d\n", reqs_sent);
            ctr <= 0;
            state <= finish;
          end
        end // case: send_reqs_init

        send_reqs_complete : begin
          //$display("State: send_reqs_complete. Reqs_sent <= %d\n", reqs_sent);
          rd_req <= 0;
          reqs_sent <= reqs_sent + 1;
          ctr <= 0;
          state <= send_reqs_init;
        end
  
        finish : begin
          if ((ctr % 1000) == 0) begin
            $display("State: finish. Reqs_sent: %d, read_info_pop_count: %d, read_count: %d\n", reqs_sent, read_info_pop_count, read_count);
            if (ctr > 10000) $finish;

          end

          if (counts_equal && ((ctr - counts_equal_ctr) >= 200)) begin
            $display("State: finish. Now getting test result.\n");
            $display("d0_pop_count: %d, d_0_count: %d, d1_pop_count: %d, d_1_count: %d", d0_pop_count, d_0_count, d1_pop_count, d_1_count);

            if (d0_pop_count == d_0_count && d1_pop_count == d_1_count) begin
              pass <= 1;
              fail <= 0;

            end else begin
              pass <= 0;
              fail <= 1;
            end

            ctr <= 0;
            state <= idle;

          end else if (!counts_equal && (read_info_pop_count == read_count)) begin // if (counts_equal && ((counts_equal_ctr - ctr) >= 50))
            $display("State: finish. Reqs_sent <= %d\n", reqs_sent);
            counts_equal <= 1;
            counts_equal_ctr <= ctr;
          end
          
        end // case: finish
        
        default : begin
        end
      endcase // case (state) 
    end // else: !if(reset)
  end // always @ (negedge clk)


  //task send_random_read_req;
  //  begin
  //    @(negedge clk);
  //    repeat (1000)
  //    begin
  //      if (read_info_full) begin
  //        wait (!read_info_full);
  //        @(negedge clk);
  //      end
  //
  //      rd_req = 1;
  //      rd_req_size = $urandom%10 +1;
  //      rd_req_pu_id = $urandom % NUM_PU;
  //      rd_req_d_type = $urandom % 2;
  //      //rd_req_d_type = 0;
  //      read_count = read_count + rd_req_size;
  //      //$display ("Requesting %d reads of type %d", rd_req_size, rd_req_d_type);
  //      if (rd_req_d_type == 0)
  //        d_0_count = d_0_count + rd_req_size;
  //      else
  //        d_1_count = d_1_count + rd_req_size;
  //      @(negedge clk);
  //      rd_req = 0;
  //    end
  //    wait (read_info_pop_count == read_count);
  //    repeat (100) @(negedge clk);
  //    if (d0_pop_count == d_0_count && d1_pop_count == d_1_count)
  //      status.test_pass;
  //    else
  //      status.test_fail;
  //  end
  //endtask // send_random_read_req

  always @(posedge clk)
    if (reset)
      inbuf_empty <= 0;
    else
      inbuf_empty <= (read_count == read_info_pop_count) || (inbuf_empty_rands[inbuf_empty_idx] == 0);

  always @(posedge clk)
    if (reset)
      read_info_pop_count <= 0;
    else
      read_info_pop_count <= read_info_pop_count + inbuf_pop;

  always @(posedge clk)
    if (reset)
      d0_pop_count <= 0;
    else
      d0_pop_count <= d0_pop_count + (stream_push && !stream_full);

  always @(posedge clk)
    if (reset)
      d1_pop_count <= 0;
    else
      d1_pop_count <= d1_pop_count + (buffer_push && !buffer_full);

  always @(posedge clk)
    buffer_full <= buffer_full_rands[buffer_full_idx];
  always @(posedge clk)
    stream_full <= stream_full_rands[stream_full_idx];


endmodule
