//---------------------------------------------------------------------------------------
//  Project:  ADPCM Encoder / Decoder
//
//  Filename:  tb_ima_adpcm.v      (April 26, 2010 )
//
//  Author(s):  Moti Litochevski
//
//  Description:
//    This file implements the ADPCM encoder & decoder test bench. The input samples
//    to be encoded are read from a binary input file. The encoder stream output and
//    decoded samples are also compared with binary files generated by the Scilab
//    simulation.
//
//---------------------------------------------------------------------------------------
//
//  To Do:
//  -
//
//---------------------------------------------------------------------------------------
//
//  Copyright (C) 2010 Moti Litochevski
//
//  This source file may be used and distributed without restriction provided that this
//  copyright statement is not removed from the file and that any derivative work
//  contains the original copyright notice and the associated disclaimer.
//
//  THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES,
//  INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND
//  FITNESS FOR A PARTICULAR PURPOSE.
//
//---------------------------------------------------------------------------------------
// Refactored to run on Cascade in April 2019 by Tiffany Yang

include ima_adpcm_enc.v;
include ima_adpcm_dec.v;

module test(clk);
  parameter BUFFER_BYTES = 32;

  // Truncated for development
  parameter TOTAL_IN_BYTES = 348160;
  parameter TOTAL_ENC_BYTES = 174080; 
  parameter TOTAL_DEC_BYTES = 348160;

  parameter MAIN0 = 0;
  parameter MAIN1 = 1;
  parameter MAIN2 = 2;

  parameter IN0 = 0;
  parameter IN1 = 1;
  parameter IN2 = 2;
  parameter IN3 = 3;
  parameter IN4 = 4;
  parameter IN5 = 5;

  parameter ENC0 = 0;
  parameter ENC1 = 1;
  parameter ENC2 = 2;
  parameter ENC3 = 3;
  parameter ENC4 = 4;

  parameter DEC0 = 0;
  parameter DEC1 = 1;
  parameter DEC2 = 2;
  parameter DEC3 = 3;
  parameter DEC4 = 4;

  parameter TESTS_TO_RUN = 1;

  
  input wire clk;

  //---------------------------------------------------------------------------------------
  // internal signal
  reg rst;        // global reset
  reg [15:0] inSamp;    // encoder input sample
  reg inValid;      // encoder input valid flag
  wire inReady;      // encoder input ready indication
  wire [3:0] encPcm;    // encoder encoded output value
  wire encValid;      // encoder output valid flag
  wire decReady;     // decoder ready for input indication
  wire [15:0] decSamp;  // decoder output sample value
  wire decValid;      // decoder output valid flag
  integer sampCount, encCount, decCount;

  reg [7:0] intmp, enctmp, dectmp;
  reg [3:0] encExpVal;
  reg [15:0] decExpVal;
  reg [31:0] dispCount;

  reg inDone, encDone, decDone;

  reg[31:0] testCount;

  reg[7:0] inReg, decReg;

  // Variables to read file input into before copying to in-mem buffer
  reg[(BUFFER_BYTES << 3) - 1:0] inVal;
  reg[(BUFFER_BYTES << 3) - 1:0] encVal;
  reg[(BUFFER_BYTES << 3) - 1:0] decVal;

  reg[15:0] inIdx, encIdx, decIdx;

  // Buffers to hold file content
  reg[(BUFFER_BYTES << 3) - 1:0] inBuf [(TOTAL_IN_BYTES / BUFFER_BYTES) - 1:0];
  reg[(BUFFER_BYTES << 3) - 1:0] encBuf [(TOTAL_ENC_BYTES / BUFFER_BYTES) - 1:0];
  reg[(BUFFER_BYTES << 3) - 1:0] decBuf [(TOTAL_DEC_BYTES / BUFFER_BYTES) - 1:0];
  reg[31:0] inBytesRead, encBytesRead, decBytesRead;


  reg[3:0] mainState;
  reg[3:0] inState;
  reg[3:0] encState;
  reg[3:0] decState;

  reg[31:0] mCtr;
  reg[31:0] iCtr;
  reg[31:0] eCtr;
  reg[31:0] dCtr;

  initial begin
    $display("Initializing");

    testCount = 0;

    mCtr = 0;
    mainState = 0;

    iCtr = 0;
    inState = 0;

    eCtr = 0;
    encState = 0;

    dCtr = 0;
    decState = 0;

    
    inBuf[0] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[1] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[2] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[3] = 256'h0000000000000000000000000000000000000000000000000000000000000000;    
    inBuf[4] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[5] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[6] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[7] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[8] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[9] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[10] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[11] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[12] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[13] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[14] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[15] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[16] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[17] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[18] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[19] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[20] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[21] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[22] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[23] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[24] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[25] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[26] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[27] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[28] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[29] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[30] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[31] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[32] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[33] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[34] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[35] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[36] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[37] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[38] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[39] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[40] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[41] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[42] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[43] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[44] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[45] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[46] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[47] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[48] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[49] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[50] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[51] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[52] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[53] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[54] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[55] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[56] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[57] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[58] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[59] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[60] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[61] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[62] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[63] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[64] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[65] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[66] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[67] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[68] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[69] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[70] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[71] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[72] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[73] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[74] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[75] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[76] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[77] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[78] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[79] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[80] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[81] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[82] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[83] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[84] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[85] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[86] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[87] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[88] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[89] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[90] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[91] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[92] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[93] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[94] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[95] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[96] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[97] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[98] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[99] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[100] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[101] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[102] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[103] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[104] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[105] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[106] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[107] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[108] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[109] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[110] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[111] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[112] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[113] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[114] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[115] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[116] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[117] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[118] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[119] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[120] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[121] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[122] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[123] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[124] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[125] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[126] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[127] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[128] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[129] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[130] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[131] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[132] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[133] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[134] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[135] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[136] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[137] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[138] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[139] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[140] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[141] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[142] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[143] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[144] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[145] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[146] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[147] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[148] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[149] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[150] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[151] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[152] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[153] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[154] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[155] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[156] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[157] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[158] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[159] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[160] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[161] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[162] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[163] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[164] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[165] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[166] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[167] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[168] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[169] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[170] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[171] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[172] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[173] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[174] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[175] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[176] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[177] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[178] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[179] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[180] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[181] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[182] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[183] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[184] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[185] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[186] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[187] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[188] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[189] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[190] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[191] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[192] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[193] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[194] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[195] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[196] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[197] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[198] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[199] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[200] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[201] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[202] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[203] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[204] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[205] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[206] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[207] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[208] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[209] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[210] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[211] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[212] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[213] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[214] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[215] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[216] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[217] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[218] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[219] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[220] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[221] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[222] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[223] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[224] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[225] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[226] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[227] = 256'h000000000000ffff000000000000000000000000000000000000000000000000;
    inBuf[228] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[229] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[230] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[231] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[232] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[233] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[234] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[235] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[236] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[237] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[238] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[239] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[240] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[241] = 256'h0000000000000000ffff00000000000000000000000000000000000000000000;
    inBuf[242] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[243] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[244] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[245] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[246] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[247] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[248] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[249] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[250] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[251] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[252] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[253] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[254] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[255] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[256] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[257] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[258] = 256'h0000000000000000000000000000010001000000000000000000ffff00000000;
    inBuf[259] = 256'h0000000000000000ffff00000000000000000000ffffffff0000000000000000;
    inBuf[260] = 256'h00000000000000000000ffff000000000000000000000000000000000000ffff;
    inBuf[261] = 256'h0000000000000000000000000000ffff00000000ffffffff0000000000000000;
    inBuf[262] = 256'h0000ffff00000000000000000000000000000000010000000000000000000000;
    inBuf[263] = 256'h0000000000000100010000000000010000000000000000000000000001000000;
    inBuf[264] = 256'h0000000000000000000000000000000000000000ffffffff0000010000000000;
    inBuf[265] = 256'h00000000ffff0000010001000000000000000000ffff00000000000000000000;
    inBuf[266] = 256'h00000000000000000000000000000000ffff0000000000000000000000000000;
    inBuf[267] = 256'h00000000ffff0000000000000000010000000000000000000000000000000000;
    inBuf[268] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[269] = 256'h000000000000000000000000ffffffff000001000100ffffffff000000000000;
    inBuf[270] = 256'h000000000000ffff0000000000000000010000000000ffff0000010001000000;
    inBuf[271] = 256'h0000000000000000000000000000000001000000000000000000000000000100;
    inBuf[272] = 256'h0000ffff00000000ffff00000000000000000000000000000000000000000000;
    inBuf[273] = 256'h0000ffff0000010001000000000000000000ffff0000010001000000ffff0100;
    inBuf[274] = 256'h0100000000000000000000000000010000000000000000000000000000000000;
    inBuf[275] = 256'h0000000001000000000000000000000000000000000000000100010000000000;
    inBuf[276] = 256'h00000000010000000000000000000000000000000000000000000000ffff0000;
    inBuf[277] = 256'h00000000000000000000ffffffff000001000000000000000000000000000000;
    inBuf[278] = 256'h0000000000000000ffff00000100000000000000000000000100010000000000;
    inBuf[279] = 256'h00000000000000000000000001000100ffffffff00000000ffffffff00000000;
    inBuf[280] = 256'h00000000000000000000ffff0000010000000000000000000000000000000000;
    inBuf[281] = 256'h0000000000000000010000000000000000000000000000000000000000000000;
    inBuf[282] = 256'h00000000000000000000ffff0000000000000000000000000000000000000000;
    inBuf[283] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[284] = 256'h00000000000000000000000000000000ffff0000000000000000000000000000;
    inBuf[285] = 256'h0000000000000000000000000000000000000000000001000100000000000000;
    inBuf[286] = 256'h00000000000000000000010000000000000001000000ffff0000000000000000;
    inBuf[287] = 256'h000000000000000000000000ffffffff00000000000000000000000000000000;
    inBuf[288] = 256'h0000000000000100010000000000000000000000000000000000000000000000;
    inBuf[289] = 256'h00000000000000000000ffff000000000000ffff000000000000ffff00000000;
    inBuf[290] = 256'h0000000000000000000000000000ffff0000010001000000ffff000000000000;
    inBuf[291] = 256'h00000000000001000000000000000000ffff000001000100000001000000ffff;
    inBuf[292] = 256'h00000000010000000000000000000000ffff0000000000000000000000000000;
    inBuf[293] = 256'h0000ffffffff00000000000000000000000000000000000000000000ffffffff;
    inBuf[294] = 256'h00000100000000000000000000000000ffffffff00000100000000000000ffff;
    inBuf[295] = 256'hffff000001000000000000000000000000000000000000000000000001000000;
    inBuf[296] = 256'h000000000000ffff000000000000000000000000000000000000000001000100;
    inBuf[297] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[298] = 256'hffff000000000000000001000100000000000000000000000000000000000100;
    inBuf[299] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[300] = 256'h000000000000000000000000ffffffff000001000000ffffffffffff00000000;
    inBuf[301] = 256'h0000000000000000000000000000000000000000000000000000000001000000;
    inBuf[302] = 256'h0000000000000000010000000000000000000000000000000000000000000000;
    inBuf[303] = 256'h000000000000ffffffff000000000000ffff0000000000000000000000000000;
    inBuf[304] = 256'h0000000000000000000000000000000000000000000000000100000000000000;
    inBuf[305] = 256'h0000ffff00000100010000000000000000000000000000000000000000000100;
    inBuf[306] = 256'h0100000000000000000000000000000000000000000000000000000000000000;
    inBuf[307] = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    inBuf[308] = 256'h000000000000010001000000ffff000000000000000000000000000000000000;
    inBuf[309] = 256'h0000000000000000000000000000000000000000000000000000000001000000;
    inBuf[310] = 256'h0000000000000000000000000000000000000100000000000000000000000000;
    inBuf[311] = 256'h00000000000000000000000000000000000000000000ffffffff00000000ffff;
    inBuf[312] = 256'hffff00000000000000000000000000000000ffff000000000000000000000100;
    inBuf[313] = 256'h010000000000000001000000000000000000000001000100000000000000ffff;
    inBuf[314] = 256'hffff000000000000000000000000000000000000000000000000000000000000;
    inBuf[315] = 256'h0000000000000000000000000000ffff00000000ffffffff010001000000ffff;
    inBuf[316] = 256'h000000000000000000000000000000000000000000000000000001000000ffff;
    inBuf[317] = 256'hffff000000000000010000000000ffffffff0000000000000000010000000000;
    inBuf[318] = 256'h000000000000000000000000000000000000000000000000000000000000ffff;
    inBuf[319] = 256'h0000000000000000010000000000000000000000000000000000000000000000;
    inBuf[320] = 256'h0000010000000000000000000000000000000000000000000000000000000000;
    inBuf[321] = 256'h000000000000010000000000000000000000000000000100000000000000ffff;
    inBuf[322] = 256'h00000000000000000000000000000000ffffffff0000ffff0000010000000000;
    inBuf[323] = 256'h00000000ffffffffffffffffffff000000000000000001000000ffff00000100;
    inBuf[324] = 256'hffffffff00000000000000000000000001000100ffffffff0000000000000000;
    inBuf[325] = 256'h01000000000000000000ffffffff00000000000001000100010000000000ffff;
    inBuf[326] = 256'h00000000ffff000000000000010000000000ffff000001000000000000000100;
    inBuf[327] = 256'h01000000ffff000001000100000000000000ffffffff00000000000000000000;
    inBuf[328] = 256'h000000000000000000000000000000000000ffff000001000000ffff00000000;
    inBuf[329] = 256'h0000000001000000000000000000000000000100000000000000000000000000;
    inBuf[330] = 256'h00000000000000000100000000000000000000000000ffffffff000001000000;
    inBuf[331] = 256'h00000000ffffffff000000000000ffffffff0000000000000000000000000000;
    inBuf[332] = 256'h0000000000000100fffffffffffffefffbfffbff00000d0019001200f7ffe9ff;
    inBuf[333] = 256'hf8ff0000ecffdfffedfffcff02000f0019000a00f4ffeffff9ff03000b000f00;
    inBuf[334] = 256'h0c0009000a000c000f001a0027002e002a001600ffff0a002e002800f0ffd1ff;
    inBuf[335] = 256'he2ffedffe3fff8ff250032002200240033002d0015000600040009000e000700;
    inBuf[336] = 256'hf8fff2fff7fffcfff9ffe7ffcbffc3ffd5ffd5ffbeffceff0b0028001c002d00;
    inBuf[337] = 256'h48001900c1ffb6fff0ff0300d9ffb2ffaaffb4ffcaffe0ffe8ffeaffebffe2ff;
    inBuf[338] = 256'hdaffe4fff9ff140031002400e0ffb1ffcefff9ff0e0047008300580003002300;
    inBuf[339] = 256'h7600370091ff58ffaaff020025002a00190008000f0012000400fdfff0ffc4ff;
    inBuf[340] = 256'h9fff9aff8cff95ff00005900280007005b004400a2ffc0ff6000d1ff46ff2202;
    inBuf[341] = 256'h87078d0aec093e09120a4e0a6b093609bb099e094909b709220abd0949092909;
    inBuf[342] = 256'hb6080108ba079a072f070507590771072b072d075207ee064506eb05a5054605;
    inBuf[343] = 256'h5805f0056706770664063f0610062006680688068406a406cb06d20608079b07;
    inBuf[344] = 256'h4e080209bb092d0a270afa09ec09e209e609390ac50a4d0bc80b260c3b0c360c;
    inBuf[345] = 256'h5f0c790c3b0cea0bc30b880b3a0b450b9b0bc30bb60bba0ba90b540bfb0abe0a;
    inBuf[346] = 256'h640afb09c409a1095e092f0938092d09ee08b5087808ff0773072207ff06e906;
    inBuf[347] = 256'hf6061b072b07340754076d076b0776078c078207640767077d079407cf073a08;
    inBuf[348] = 256'ha108f8085d09bb09ee09090a1e0a1d0a0a0a0f0a3c0a800ad50a330b780b960b;
    inBuf[349] = 256'h9a0b810b430b030be30ad70ad00ad50adf0ad00aa50a740a420a0b0ada09b809;
    inBuf[350] = 256'h920963093a091409e708bc0894085e081008bc076e07330723073e0761077007;
    inBuf[351] = 256'h6c0757072907f006cd06ca06dc06ff062d075607720786079807a807bd07d707;
    inBuf[352] = 256'hed07fe070f081f082f08410854085e08620864086308630870088b089f089e08;
    inBuf[353] = 256'h86084c08eb0778071607d706b806af06ad069b066f062606c4055405ee049b04;
    inBuf[354] = 256'h5f043b042b04220413040204f403e203cc03b6039c037403470326031c032b03;
    inBuf[355] = 256'h50038103ab03be03b903a6039803a103c603ff0344048704b804d204e004ec04;
    inBuf[356] = 256'h09053c057605ae05d805ed05ee05e305d305c105ad058e0559051005b8046404;
    inBuf[357] = 256'h2104f303d103ac036e03100398021602a10146010901df00ba008d0052000e00;
    inBuf[358] = 256'hc5ff81ff45ff0dffd5fe9efe6afe3ffe20fe0efe04fef8fddffdb6fd86fd58fd;
    inBuf[359] = 256'h3bfd39fd59fd95fde0fd2cfe73feaffeddfe05ff32ff6bffb0ffffff51009e00;
    inBuf[360] = 256'hd700f600ff00f800e700d400c600bd00b2009b00760048001100daffabff87ff;
    inBuf[361] = 256'h69ff4dff2cff0affecfecdfeaefe88fe4ffefefd9bfd32fdd8fc98fc6dfc4efc;
    inBuf[362] = 256'h2dfcf9fbb2fb65fb1cfbe1fab6fa90fa69fa3efa0cfae0f9c8f9c4f9dbf908fa;
    inBuf[363] = 256'h39fa68fa8cfa9dfa9efa9afa94fa9cfab9fae5fa22fb6efbb6fbf7fb29fc3efc;
    inBuf[364] = 256'h35fc12fcd9fba3fb81fb73fb7efb9afbacfbabfb94fb63fb2cfbf9facafaaffa;
    inBuf[365] = 256'ha6fa9dfa94fa86fa64fa30faf1f9abf973f954f946f94df95ff95cf93ff906f9;
    inBuf[366] = 256'hacf849f8eff7a9f791f7adf7e7f739f88df8bdf8c1f896f840f8e5f7a4f78cf7;
    inBuf[367] = 256'hb5f71bf897f815f978f9a0f998f96ef92ff900f9f4f802f933f97cf9c0f9fef9;
    inBuf[368] = 256'h2efa3bfa34fa1bfae6f9adf97df952f93df93cf932f920f9fbf8b1f85cf811f8;
    inBuf[369] = 256'hd3f7b7f7b7f7b2f7a3f77df72df7cff67bf62ef6fff5f3f5f6f50df62ff642f6;
    inBuf[370] = 256'h4df648f61cf6e0f5a8f573f560f57af5abf5f4f541f671f692f6a9f6a7f6a7f6;
    inBuf[371] = 256'hb7f6c6f6e7f61bf750f795f7e5f720f856f887f89bf8acf8c8f8e3f810f94bf9;
    inBuf[372] = 256'h74f992f99ef982f95bf93cf91af909f907f9f9f8e9f8daf8b6f896f87bf848f8;
    inBuf[373] = 256'h0cf8ccf779f737f715f701f708f71af70ef7f0f6c3f67ef645f625f608f6fcf5;
    inBuf[374] = 256'hfbf5e6f5cef5bef5a5f5a0f5b1f5bef5d7f5fbf512f630f65ef684f6b1f6e5f6;
    inBuf[375] = 256'h05f729f757f77ef7b8f709f84ff891f8ccf8e5f8f1f8f7f8e7f8ddf8dff8d6f8;
    inBuf[376] = 256'hddf8fcf81af945f978f991f99ef99ef981f96af966f95ff966f977f96ff958f9;
    inBuf[377] = 256'h36f9fbf8c7f8a3f875f850f830f8f8f7c2f799f771f762f769f767f767f769f7;
    inBuf[378] = 256'h5af759f773f793f7c6f703f82cf851f879f895f8bdf8f5f81ff947f96cf97bf9;
    inBuf[379] = 256'h91f9b9f9e1f916fa52fa74fa89fa96fa8ffa92faa5faaffabbfac6fabafab0fa;
    inBuf[380] = 256'hb5fac0fae3fa15fb33fb42fb43fb24fb05fbf3fae0fad5facafaa6fa7afa4ffa;
    inBuf[381] = 256'h1bfaf8f9eaf9d6f9c2f9acf984f95ff946f932f936f950f966f986f9b0f9d6f9;
    inBuf[382] = 256'h07fa42fa76faabfadffa02fb2cfb65fb9ffbe3fb29fc56fc71fc80fc81fc91fc;
    inBuf[383] = 256'hbbfcf1fc37fd82fdb6fdd8fdecfde8fde2fddefdd0fdc7fdc1fdb2fda9fdaafd;
    inBuf[384] = 256'ha9fdb0fdb9fdb0fd98fd71fd34fdf6fcc5fc9dfc8ffc91fc8ffc88fc78fc54fc;
    inBuf[385] = 256'h2dfc0afceafbd8fbd2fbccfbcefbd4fbd2fbd3fbd9fbdefbeefb0efc37fc71fc;
    inBuf[386] = 256'hb5fcf6fc3afd7dfdb8fdf3fd2efe65fe9efed3fefffe29ff4eff6cff8effbaff;
    inBuf[387] = 256'hedff280066009a00c000d200cc00bb00a5008b0076006400530046003a003300;
    inBuf[388] = 256'h340039003b00380028000300cdff8aff43ff06ffddfecefeddfe00ff2dff58ff;
    inBuf[389] = 256'h72ff74ff5eff31fff5feb7fe81fe5dfe58fe70fea5fef3fe4affa0ffe9ff1c00;
    inBuf[390] = 256'h3800440045004b0062008d00d10029018401d80119023a024302390227022002;
    inBuf[391] = 256'h2a023f025d027a02870289028102740271027a028902a302be02cf02d902d702;
    inBuf[392] = 256'hc502af0296027d027302780283029502a2029902800256022202fc01eb01f101;
    inBuf[393] = 256'h180250028602b702d702df02dc02d002be02b802c002d40208035403ad030f04;
    inBuf[394] = 256'h6104890489045c040e04c50392037f039a03d30310044d0476047e0476045a04;
    inBuf[395] = 256'h2c040204da03b503a603a503aa03c203e003f803170431043d04480446043004;
    inBuf[396] = 256'h1904fd03de03d403da03e8030a042d044204580463046504750488049b04b904;
    inBuf[397] = 256'hd404e9040c0538056b05b50501063e0672068d068e0692069806a406ca06f606;
    inBuf[398] = 256'h1b07400753074c0740072307f506cc06a3067e0676067e068c06a706b2069e06;
    inBuf[399] = 256'h79063e06f305b805890561055105430531052c0527051d051f051805ff04e604;
    inBuf[400] = 256'hbf049004750466045d04660469045e045b04560456047604a104cd04fe041605;
    inBuf[401] = 256'h11050605f004dc04ea040d0544059a05f40548069c06d306e606e606c7069806;
    inBuf[402] = 256'h7c0672067e06b006e5060e07310739072c0727071e07140715070907ee06d806;
    inBuf[403] = 256'hbd06a606a806ad06af06b406a4068006600637060e06f705da05b8059e057d05;
    inBuf[404] = 256'h5d05570556055a05690565054a052905f804c404a6048e047d047d0474046304;
    inBuf[405] = 256'h5b044d043c043704290412040404f103e203e903f203fa030b040d0403040104;
    inBuf[406] = 256'hfb03f503fe03fb03ec03dc03be039f039a03a503c403fe033204540469045b04;
    inBuf[407] = 256'h36041404f103dc03e803ff031e044904650472047b04740464045d0454044f04;
    inBuf[408] = 256'h5a0464046d04800489048d0499049e04a404b604c104c604cb04be04a1047f04;
    inBuf[409] = 256'h4d041304e403ba039f03a103ae03c003d003c0038c033e03d6026a021902e301;
    inBuf[410] = 256'hd201e801080226023a022f020502cc0180013401fd00d700ca00d800ed00fe00;
    inBuf[411] = 256'h0801f900d500aa00790051003f003b0043005700660071007f008b009b00b800;
    inBuf[412] = 256'hd600f5001701310146015d01710185019d01b001c201d701e901fd0113022202;
    inBuf[413] = 256'h270223021002f701e001cb01bf01bc01bc01bb01bc01b501aa019e018b017501;
    inBuf[414] = 256'h60014901330120010901ef00d200af008e007300600054004d0040002600fdff;
    inBuf[415] = 256'hc4ff85ff4dff25ff13ff15ff22ff30ff33ff26ff0affe5febffe9dfe86fe7afe;
    inBuf[416] = 256'h7afe83fe92fea5feb3febafeb4fea1fe88fe72fe67fe6dfe83fe9dfeb3febbfe;
    inBuf[417] = 256'hb0fe98fe7cfe65fe5bfe5ffe6bfe7efe8ffe98fe9afe93fe85fe74fe66fe5cfe;
    inBuf[418] = 256'h61fe76fe98fec7fef8fe1eff36ff39ff27ff0ffffbfef5fe08ff30ff5eff8aff;
    inBuf[419] = 256'ha3ffa1ff8bff6aff49ff3bff42ff57ff76ff92ff9fffa1ff97ff85ff78ff70ff;
    inBuf[420] = 256'h68ff64ff5dff4cff3bff25ff08ffecfecbfea0fe76fe4cfe25fe11fe0efe11fe;
    inBuf[421] = 256'h16fe0bfee1fda0fd4ffdfdfcc7fcb5fcc0fce6fc10fd28fd2dfd1cfdf5fccffc;
    inBuf[422] = 256'hadfc92fc8bfc94fca9fcd1fc03fd30fd5cfd78fd7dfd79fd6ffd65fd70fd8efd;
    inBuf[423] = 256'hb8fdeffd27fe52fe78fe97feaffecffef2fe11ff32ff4cff58ff62ff68ff69ff;
    inBuf[424] = 256'h72ff7cff81ff88ff8bff85ff7eff72ff56ff37ff10ffe0febcfea6fe9dfeabfe;
    inBuf[425] = 256'hc2fed2fedbfed1feadfe7efe4afe15fef5fdeafdedfd05fe20fe2efe2efe17fe;
    inBuf[426] = 256'he6fdaefd77fd46fd30fd31fd40fd62fd85fd9cfdacfdaefd9efd8efd7ffd73fd;
    inBuf[427] = 256'h79fd8bfda0fdbffddcfdedfdfbfd02fefcfdf8fdf4fdecfdecfdf0fdeefdf0fd;
    inBuf[428] = 256'hedfddffdd1fdc1fdacfda3fda1fd9ffda5fda9fda1fd97fd87fd71fd68fd6dfd;
    inBuf[429] = 256'h7ffda7fdd9fd04fe28fe39fe31fe21fe0efefffd04fe1bfe3bfe66fe8ffea9fe;
    inBuf[430] = 256'hb8feb7fea4fe8ffe7ffe79fe8bfeb4fee5fe1fff50ff6bff75ff6eff59ff45ff;
    inBuf[431] = 256'h36ff28ff25ff28ff27ff28ff24ff13fffbfed8fea9fe7efe5bfe43fe41fe4bfe;
    inBuf[432] = 256'h53fe53fe41fe13fedafd9ffd6cfd52fd4ffd56fd60fd60fd49fd27fdfefcd5fc;
    inBuf[433] = 256'hb9fcadfca9fcb3fcc6fcddfcfffc28fd4cfd6bfd7dfd7efd7dfd82fd95fdbffd;
    inBuf[434] = 256'hfdfd3ffe7ffeb0feccfedafee2fee4feecfef7fe00ff0aff16ff22ff36ff54ff;
    inBuf[435] = 256'h71ff8fffa4ffa7ff9eff8dff78ff6dff71ff7eff95ffadffbfffcbffd1ffcdff;
    inBuf[436] = 256'hc3ffb0ff8dff61ff2ffffafecffeb5fea6fea4fea8fea5fe9dfe8dfe74fe5afe;
    inBuf[437] = 256'h43fe2cfe1cfe16fe16fe23fe3cfe5bfe7efea2febbfecbfed1fecbfec0feb4fe;
    inBuf[438] = 256'ha5fe9bfe97fe99fea3feb7fecffeeafe04ff11ff11ff05ffebfecffebcfeb5fe;
    inBuf[439] = 256'hc2fee0fe04ff29ff47ff54ff51ff3fff1efff8fed5feb7feaafeb1fec7fee9fe;
    inBuf[440] = 256'h0eff29ff36ff35ff23ff0bfff3fee1feddfeeafe06ff32ff67ff9affc5ffdfff;
    inBuf[441] = 256'he6ffdeffcfffbfffb9ffc2ffd6fff2ff11002b003f004c005300590063007000;
    inBuf[442] = 256'h7f008e0098009d0099008f00820079007300730078007c007c00710053002300;
    inBuf[443] = 256'he3ff99ff50ff13ffeafedbfee4fefafe14ff26ff25ff0fffe5feaffe7afe54fe;
    inBuf[444] = 256'h43fe4ffe72fea2fed5fefbfe0cff0bfffbfee6fed6fed4fee3fe05ff33ff65ff;
    inBuf[445] = 256'h94ffb7ffcbffd1ffd0ffd4ffe7ff0f0048008e00d00003012001280123012001;
    inBuf[446] = 256'h2a0145017001a101c901de01d901bd019501690145012e0122011f0120011c01;
    inBuf[447] = 256'h11010001e600c2009a006f004b00390039004d006f008d009a008d0064002b00;
    inBuf[448] = 256'hf4ffccffbdffcaffe8ff09002100260018000100e5ffd3ffd6ffedff1b005700;
    inBuf[449] = 256'h9400ca00f10001010001f700ef00f4000e0136016b01a201cb01e001dd01c401;
    inBuf[450] = 256'h9e0177015501410141014f0166017f018e01900186016e015101390128012201;
    inBuf[451] = 256'h23012501250125011f011c01200129013701480153015a015e015b0153014901;
    inBuf[452] = 256'h39012a01230126013f016e01a801e301110224021d020402e501d301dc01fd01;
    inBuf[453] = 256'h34027302a802ce02e102dd02cc02b7029e028802760266025d025d025f026502;
    inBuf[454] = 256'h6a0262024d022902f801c5019a0179016801620160015e015601460132012001;
    inBuf[455] = 256'h0d01ff00f500ed00eb00ec00ef00f9000a0120013a01580174019001a901bb01;
    inBuf[456] = 256'hc901d501dd01e401ec01f101f90104021002240240025e027c0294029d029d02;
    inBuf[457] = 256'h95028a0287029202aa02cf02f8021c0339034a034a033b031c03eb02b0027102;
    inBuf[458] = 256'h3702120207020e021e0223020c02d80189012d01de00a7008c008b009500a100;
    inBuf[459] = 256'had00b900c600dc00f5000a01150112010301f500f000f8000c01240136013d01;
    inBuf[460] = 256'h38012e012e013b0152016f0185018e018c01840182019301ba01ef012b025d02;
    inBuf[461] = 256'h7e028c028702760266025b02560259025e02620264025e0249022802f701b901;
    inBuf[462] = 256'h770138010501e700da00d500d300c700ac008600560029000a00fafff9ff0500;
    inBuf[463] = 256'h15002400310039003d0044004b0055006200720083009900ad00bd00ce00da00;
    inBuf[464] = 256'he200eb00f6000801250147016c019301b301c801d201ce01c301b901b201b201;
    inBuf[465] = 256'hba01c401c701c201ab01870161013b011c010901fb00ef00e000c600a5008200;
    inBuf[466] = 256'h5f00400027001000fcffeaffd7ffc6ffbcffb4ffafffacffa7ffa2ffa2ffa4ff;
    inBuf[467] = 256'hacffbeffd3ffedff090021003800510066007b009200a700bb00cf00dd00ea00;
    inBuf[468] = 256'hf9000401110122013201450157016201650162015401400129011001f900e800;
    inBuf[469] = 256'hd800cc00c300b600a3008800600031000000cfffa6ff88ff71ff5fff4fff3bff;
    inBuf[470] = 256'h29ff1bff0fff08ff07ff03fffefef6feeafee4fee9fef7fe10ff30ff4dff66ff;
    inBuf[471] = 256'h7aff87ff96ffa9ffbdffd2ffe7fff5ff02000f001c003200520075009900b800;
    inBuf[472] = 256'hcc00da00e100e300e600ef00f700000105010201fa00f000df00cd00b8009a00;
    inBuf[473] = 256'h750047000f00d8ffa6ff78ff53ff35ff17fff9fedafeb6fe97fe7efe67fe57fe;
    inBuf[474] = 256'h4cfe45fe47fe52fe65fe84fea9fecdfeecfe02ff0aff0cff08fffffefafefbfe;
    inBuf[475] = 256'hfefe08ff16ff26ff3bff51ff63ff74ff80ff86ff88ff86ff80ff81ff88ff96ff;
    inBuf[476] = 256'hb1ffd4fff9ff1d00370043004300380021000500e3ffbcff95ff6dff47ff2bff;
    inBuf[477] = 256'h1aff0fff0bff07fffcfeeffeddfeccfec6fecefee0fefcfe19ff2fff3dff40ff;
    inBuf[478] = 256'h39ff2fff25ff1cff17ff12ff0dff0cff0aff05ff02fffafeebfed4feb3fe8afe;
    inBuf[479] = 256'h61fe3cfe21fe17fe1cfe2ffe4afe66fe7efe92fe9ffea5fea9fea8fea4fe9efe;
    inBuf[480] = 256'h95fe8bfe85fe84fe8bfe9cfeb5fed3fef8fe1aff36ff4eff5dff65ff6aff6dff;
    inBuf[481] = 256'h72ff7fff91ffa6ffbcffcfffddffe7ffe9ffe4ffddffceffb7ff9aff76ff4dff;
    inBuf[482] = 256'h23fff5fec6fe98fe68fe38fe0dfee8fdcafdb5fda5fd98fd8dfd82fd7afd78fd;
    inBuf[483] = 256'h7cfd87fd99fda8fdb3fdb6fdb2fda8fd9efd96fd93fd9afda8fdbffde0fd09fe;
    inBuf[484] = 256'h39fe6cfe99febdfed2fed7fecefebffeb0feabfeb2fec4fedffefefe18ff2aff;
    inBuf[485] = 256'h32ff2eff20ff08ffe5feb8fe82fe45fe03fec2fd86fd52fd28fd06fdecfcd8fc;
    inBuf[486] = 256'hc7fcb8fca8fc95fc81fc69fc4efc32fc16fcfefbedfbeafbf7fb18fc4efc95fc;
    inBuf[487] = 256'he9fc45fda1fdf9fd49fe8dfec5feeffe09ff12ff0dfffffeeefee4fee8fe00ff;
    inBuf[488] = 256'h28ff5aff89ffa8ffb0ff9dff72ff36fff0fea7fe60fe1ffee7fdb9fd97fd80fd;
    inBuf[489] = 256'h72fd66fd54fd37fd0bfdd3fc94fc59fc27fc03fceafbd5fbbdfb9bfb6efb3bfb;
    inBuf[490] = 256'h0afbe4fad3fadafafafa2efb6ffbb5fbf8fb33fc63fc89fca6fcc2fce3fc10fd;
    inBuf[491] = 256'h4ffda0fdfffd63fec2fe10ff44ff5aff52ff32ff01ffc7fe8bfe51fe1efef4fd;
    inBuf[492] = 256'hcefdacfd94fd83fd76fd66fd50fd32fd0cfde6fcc7fcb6fcbafcd1fcf5fc1dfd;
    inBuf[493] = 256'h3dfd4cfd46fd2bfd00fdccfc96fc66fc3ffc26fc1bfc1ffc31fc4ffc70fc8cfc;
    inBuf[494] = 256'h9afc94fc79fc50fc26fc0bfc0bfc2efc71fcc9fc28fd7ffdc6fdf8fd18fe2bfe;
    inBuf[495] = 256'h35fe3afe3afe34fe2bfe1ffe15fe12fe17fe25fe3afe51fe68fe7ffe96feaefe;
    inBuf[496] = 256'hc9fee3fef7fe00fffcfeebfed5fec2febcfec7fee1fe03ff21ff33ff36ff30ff;
    inBuf[497] = 256'h2bff36ff59ff97ffe7ff3c008600bc00de00f600130140018301d6012a027002;
    inBuf[498] = 256'h9902a1028f026d024b022f021e0213020802fa01ec01e201e401f3010d022902;
    inBuf[499] = 256'h3e0246024102380236024a027802c2021f038203db031e0440043c041304cc03;
    inBuf[500] = 256'h6e030b03b3026c0239021602f901d801b101810151012c011201ff00e900bb00;
    inBuf[501] = 256'h6a00faff72ffedfe8cfe59fe5afe83feb5fed9fee0fec9fea1fe76fe5bfe55fe;
    inBuf[502] = 256'h55fe55fe4cfe31fe18fe11fe27fe71feedfe83ff2b00ca004701ae01fd013902;
    inBuf[503] = 256'h7a02b702e60206030403dc029d024e020e02f40102024202a50207035a038803;
    inBuf[504] = 256'h840361032603e402b5029002740268025a0251025c027e02c8023a03bd034a04;
    inBuf[505] = 256'hbd04f104f104b6044404ca034f03db028f025c023d02450262028f02dd023403;
    inBuf[506] = 256'h8e03ec03300451045b044e043804260425043d04560475049e04b104bc04d304;
    inBuf[507] = 256'hd904dc04e804d704b90491043704c40342039002d6012f018d00280025005f00;
    inBuf[508] = 256'hf900e101e502f103d1046d05c405d105b505830541051805fd04e004e8040705;
    inBuf[509] = 256'h2d058405fb0580062607c4074108a908e208e908d708ae0877083c08fc07b307;
    inBuf[510] = 256'h5a070607c1068f06a106f5066e071708b40808092909e9084108740767063405;
    inBuf[511] = 256'h2a041c033902d001a001cd0171021a03c4034b043d04c703c7020f012eff16fd;
    inBuf[512] = 256'hb8fac6f817f77df576f48af380f2c8f1eaf011f004f075f0aaf126f4fdf6c5f9;
    inBuf[513] = 256'h73fc14fea7feddfed9fe59ff1b0109043308550dc3123918671d042212264829;
    inBuf[514] = 256'h822ba52c6f2c3f2b9c29ec273c273e28ee2a8f2fcd358e3c1d43c248764cd34d;
    inBuf[515] = 256'hd14c49496343bf3bd9321e297b1f9816790eb0075f0288fdeff834f4d9ed95e5;
    inBuf[516] = 256'hdddb22d056c33cb7e4ab80a2419c9098a0978399189d5fa240a9b9b0ccb840c1;
    inBuf[517] = 256'h30c984d017d7b5dcc3e191e6cbeb07f23af9dc01d40b10167f20a12a2a33533a;
    inBuf[518] = 256'hfe3f4443b8446c44ab413c3d6e37fe2f1d287820f1187412430d94083a04d4ff;
    inBuf[519] = 256'h65fa8ef36bebeae148d734cc22c148b645ac8da33b9c03975394d493aa958d99;
    inBuf[520] = 256'h389e10a39ea7e3aaccacc9adf5ade0ad5faed8af85b2a0b632bcdcc250ca7ed2;
    inBuf[521] = 256'hc7dab8e26fea3bf19ff616fb2cfeb7ffd500780191016602d10346057107ca09;
    inBuf[522] = 256'h620b970c080d1d0c560a9507700349fefaf735f086e730de42d48fcac5c102ba;
    inBuf[523] = 256'hcab384afcaac61ab17ab12abe6aa87aa91a951a856a795a6bfa655a8efaa51af;
    inBuf[524] = 256'h87b5efbce0c51ed091da04e50fef7bf75afec80369071d0a5d0c060ed70f9c11;
    inBuf[525] = 256'h96122813e5123c110d0f5a0cd8085a059601e5fcb8f79ef110eacde1f1d871cf;
    inBuf[526] = 256'h53c6fdbd62b631b0aeab88a8dea6c9a6cfa76da974ab69ad7daec0ae95aeb5ad;
    inBuf[527] = 256'hb0acbeacc3adb3af69b333b8d0bc6bc161c56cc725c800c88ec61dc5c5c4f3c4;
    inBuf[528] = 256'h7cc60bca15ceebd225da37e275e987f06bf72dfe1806680f021a9126b6347b43;
    inBuf[529] = 256'h72529560906cc075bf7b587efc7d9e7b27784c74e970476eab6b9b687c64cf5d;
    inBuf[530] = 256'hfb532647c13642231c0ee6f7c8e19acdfabb7fad0fa3419c7e987d972798a799;
    inBuf[531] = 256'hcd9b349e40a1e4a54daca9b46abf30cc71daede9fef9160a371a1b2a5939f747;
    inBuf[532] = 256'h6f555261b26bf673d8798e7d127f6a7e257cab781474c46e0e69d5620b5cc654;
    inBuf[533] = 256'hdd4c2644bd3aae30e825a71a500f080437f996ef63e7c8e04bdcd7d9f9d8ced9;
    inBuf[534] = 256'hf6db94dea6e113e522e8feeaf7ed83f0c3f226f536f702f90bfbeefca8feb400;
    inBuf[535] = 256'ha2023c04e7053407bb07d20739079d057e030a011dfe39fbcff8e0f6bef5bbf5;
    inBuf[536] = 256'hcaf6d3f8e5fbc1ffe7031e08170c5a0fd811b713f114d615e6162b18c319ed1b;
    inBuf[537] = 256'h651ed4202e23162525265b268f2574231020721b81156d0e92063cfedef5ebed;
    inBuf[538] = 256'h9fe638e0dada55d68bd278cfe6ccc2ca31c928c8b7c71ec854c947cb22ceded1;
    inBuf[539] = 256'h71d602dc82e2c4e9bbf116fa7602ac0a67126619a01fef243b29ba2c772f6831;
    inBuf[540] = 256'hbc3274336833b5328331c42f8d2d0e2b46282225ab21d91d8d19d014c00f740a;
    inBuf[541] = 256'h3205520001fc60f897f594f32ff25ef100f1e4f01af199f117f288f2edf20ff3;
    inBuf[542] = 256'h01f31bf370f328f49af5b7f750fa61fd97009e037b0615095b0b990df70f6612;
    inBuf[543] = 256'hf814a5172d1a721c681ef11f13210022d4228f234b241525ba2516261b268125;
    inBuf[544] = 256'h2b243522821f0f1c2418c513fb0e240a5905ac007dfcd2f879f580f2aeefa9ec;
    inBuf[545] = 256'h6de9f6e54ae2c6deaddb2ed99cd70ad755d764d801daf1db21de85e020e305e6;
    inBuf[546] = 256'h29e978ecd5ef11f313f6cef839fb75fd92ff8a017e036105020761086309da09;
    inBuf[547] = 256'hf309c40925093908fc062505d1021e00ecfc9bf992f6bff363f1afef3fee02ed;
    inBuf[548] = 256'h00ecc7ea51e9d4e716e62ee467e2a2e0f5de8cdd34dc06db35da9cd95cd998d9;
    inBuf[549] = 256'h0fdabbda87db1ddc84dcbfdcb6dcb6dce1dc24ddd0dddede0de08ae137e3d1e4;
    inBuf[550] = 256'ha3e6b0e8bbea13eda5ef0ef26ff4a8f65af8b9f9d0fa62fbb4fbddfba5fb45fb;
    inBuf[551] = 256'hcffa15fa4bf97ff870f738f6d4f4f4f2a2f0dfed7deab7e6cbe2c4de07dbd4d7;
    inBuf[552] = 256'h1bd51dd3e1d119d1e9d046d1d3d1bdd208d45bd5ebd6b6d85eda24dc24de17e0;
    inBuf[553] = 256'h67e242e55ae8ecebe7efb6f36ef7fafae0fd5e008002ed03dd044005be04a503;
    inBuf[554] = 256'hfc0198fffafc3ffa41f769f4a7f1a9eebbebb6e842e5ade1fcdd01da2fd6bad2;
    inBuf[555] = 256'h8fcf07cd44cb1fcabec92bca2ccba4cc76ce63d033d2d5d34fd58cd6a9d7f6d8;
    inBuf[556] = 256'h5bdad0db9bdd75dfe9e02ae209e312e3abe20fe2f1e0d1df2cdfc3defbde40e0;
    inBuf[557] = 256'h07e24ae43fe716ea81ecf2eefdf09ff2e0f410f87dfc3a038d0c281809266135;
    inBuf[558] = 256'hc8443b53985fc4685a6e7c709c6f7a6c12685e63d65ebf5a39579f53394fa649;
    inBuf[559] = 256'hf0416f37692acc1af8086bf60ae4cdd277c4aab97bb260afaaaf4fb2e0b654bc;
    inBuf[560] = 256'hfbc114c84aceb1d412dc56e4a1ed86f85b048310271dd82961360743414fac5a;
    inBuf[561] = 256'h5a65986edc75457b6a7e007f7e7d157ad2744b6e0767415f5957c24f9a48cf41;
    inBuf[562] = 256'h713b5d35232f9528b921611ab612430b400406fe43f90bf62ef4e6f3e9f491f6;
    inBuf[563] = 256'hfbf8fbfbc9fe81013f043f068e078d089e08d107ca062e051d035f01b7ff23fe;
    inBuf[564] = 256'h40fdb8fc49fc55fc81fc7cfc9afc9dfc38fcb8fb20fb65fae0f9eaf9bffa96fc;
    inBuf[565] = 256'h91ffba03c7085f0e3e14d319a61ea5229325562748287f280d28562770266125;
    inBuf[566] = 256'h7424a323c022d621af20df1e431cbc1811144c0eb407820009f9cdf12aeb4ce5;
    inBuf[567] = 256'h71e0b1dcfcd960d8ced726d872d988db32de6fe106e5c1e8b7ecc9f0e1f43cf9;
    inBuf[568] = 256'hcbfd84029e07e80c3712a917e61c9f21e4256129bf2b1f2d582d432c322a5027;
    inBuf[569] = 256'hb823d81f031c581809153912e70ffc0d660c0c0bb9094c08d0063a05a6036102;
    inBuf[570] = 256'h860126017d01830211043206cf08920b5f0e1a115c13f714fc154116c815ed14;
    inBuf[571] = 256'hb9132a1299100f0f5f0dc30b4b0ada08ba070e07b506ca063807b6074308d908;
    inBuf[572] = 256'h6909140aef0a0a0c6d0d040fd810e312fa1436179619d61b031efe1f5321f421;
    inBuf[573] = 256'hc5216d20121ef11a1317e312b40e9a0ad0065a030b00ebfcdef9bcf69cf36ef0;
    inBuf[574] = 256'h34ed27ea4ee7d3e412e311e2eee1d6e28be4dfe6bae9b7ec9cef67f2ecf42cf7;
    inBuf[575] = 256'h56f969fb6cfd64ff3001b602df039304e204d3045f04a903c502af017a0018ff;
    inBuf[576] = 256'h6cfd82fb50f9c6f61bf472f1c5ee47ec11eaf4e70de67fe424e31fe29ee16de1;
    inBuf[577] = 256'h89e100e27ee2ede267e3b1e3e0e336e492e402e5a5e539e6afe607e710e7f2e6;
    inBuf[578] = 256'hcce67ce63ee60ee69de507e535e4eee29ae165e047dfbfdedcde59df67e0c4e1;
    inBuf[579] = 256'hf7e23ee48be5a4e6fce7a2e957eb5eed8fef7ef149f3d9f4faf5f5f6d3f764f8;
    inBuf[580] = 256'hd6f815f9e7f86ff8b2f78df630f5aaf3def1efefebedb2eb60e910e7b8e492e2;
    inBuf[581] = 256'hbfe022dfe5dd13dd63dcf7dbeddb0cdc93dcb1dd1adff0e050e3c6e554e8f9ea;
    inBuf[582] = 256'h41ed43ef14f173f2c1f33bf5a2f63bf80afa9cfb12fd54fef3fe2cfff9fe14fe;
    inBuf[583] = 256'hd5fc2cfbd6f844f67ff367f09fed4beb39e9cce7e5e602e642e58fe496e3a1e2;
    inBuf[584] = 256'he2e143e1f0e0f8e020e158e1aae104e273e233e351e49fe51fe7afe8c3e93dea;
    inBuf[585] = 256'h3bea73e9ede72de62ce4dfe1c0dfd8dde6db3bda09d918d8a9d7fcd7bed8e6d9;
    inBuf[586] = 256'h8edb2bdd8fde04e039e12ce2a3e3c5e5c0e88fed81f471fdbd082216b724e733;
    inBuf[587] = 256'hd04232503b5b3e63bf67da68fd66e4627d5da1571452264dc048a144f73fd139;
    inBuf[588] = 256'hb531f9265e199f0962f881e699d5b7c699ba36b2b1adb5ac05afc1b302ba37c1;
    inBuf[589] = 256'h75c85bcf0bd648dc6fe243e9c4f033f90203b40df918d624a830123c20474951;
    inBuf[590] = 256'h2d5ac4617467c06abf6b556a7266a6609c59b9519149da41c93a5a34d42e202a;
    inBuf[591] = 256'hc125a321aa1d5619a514d90fdb0aed05ab0127fe7bfb23fa0efae1fab8fc4aff;
    inBuf[592] = 256'hd6015704b1062208bf08c808b3079505e90263ff26fbd4f659f2dced0feafee6;
    inBuf[593] = 256'hb5e49be389e33de4b6e59ce793e985eb4cedcfee2df0acf199f322f68ef915fe;
    inBuf[594] = 256'h7c0395094510f816391dda225327522adf2bcd2b2a2a5c279e235b1f101bdd16;
    inBuf[595] = 256'heb124f0fd60b6a08e8041301dafc33f810f389edb0e7bee107dcc2d645d2e3ce;
    inBuf[596] = 256'habccc3cb40ccf6cdd2d0a4d413d9f5ddfee2d1e771ecb5f065f4c1f7d1fa79fd;
    inBuf[597] = 256'h0f00b40267058a084a0c95108c15eb1a2020cf2475287c2ace2a8529c2260023;
    inBuf[598] = 256'he01eba1ad7168a13ef10ec0e810d990cea0b410b790a3f095807c5049001eefd;
    inBuf[599] = 256'h65fa78f78df500f5f1f512f8fffa55fe7f0126044e06c7078508d608a808cb07;
    inBuf[600] = 256'h8c060005230383018100440037015f035906ef09b70d30114414e416fe18c81a;
    inBuf[601] = 256'h631cd41d211f47204c212b22e822c223c224d5251d275928fb28d0288027b124;
    inBuf[602] = 256'h9d20801b9b158e0fb70939045fff1bfb45f704f444f1f9ee51ed27ec3deb7cea;
    inBuf[603] = 256'h94e953e8e6e674e552e410e4ece4f4e628ea2bee89f2faf631fbfafe69029105;
    inBuf[604] = 256'h6808dd0ad80c270ea10e4c0e540df10b6b0a16091a086207cd061e06f6042903;
    inBuf[605] = 256'hbf00c1fd7afa40f71bf42ff19aee14eca3e992e7c5e571e408e45ce446e5cee6;
    inBuf[606] = 256'h63e896e960ea77eadee901e9f9e7fce64fe6bde539e5cbe442e4bde370e352e3;
    inBuf[607] = 256'h97e33ee4f3e49de5ece578e577e418e388e176e042e0eee0aee23ae5fae7c9ea;
    inBuf[608] = 256'h6ced9eef89f130f382f4a9f586f6e1f6d9f673f6c2f52cf5daf4c5f40ff589f5;
    inBuf[609] = 256'hc4f59df5f3f496f3c2f1b0ef70ed4ceb64e98fe7e6e569e4dce27de18ee0f9df;
    inBuf[610] = 256'h05e0e4e045e227e472e6abe8d4eaefecacee42f0d9f130f37df4d3f5e9f6f8f7;
    inBuf[611] = 256'h0ef9f0f9e8faf8fbd4fca5fd3bfe36feccfde3fc58fba2f9d9f7fef596f495f3;
    inBuf[612] = 256'hbcf249f2f9f172f1f3f066f0abef1fefc5ee6cee40ee27eee2ed82ed0ded70ec;
    inBuf[613] = 256'hd0eb58eb09ebe6ea08eb69ebe2eb82ec3fedc6ed16ee36eebceda3ec38eb4be9;
    inBuf[614] = 256'hefe6ace47ce24be093de52dd3ddc90db4adb02dbddda04db28db8bdb91dcf7dd;
    inBuf[615] = 256'hdfdfa7e2d6e52de903ed21f187f507fb1502f40a3616cc230c332443db52cb60;
    inBuf[616] = 256'hd36b21736676ca75ef71ee6bbd64435d69566750204b8546b641bc3b27341e2a;
    inBuf[617] = 256'h231dd20da2fc7bea37d926ca59be09b751b4beb5d9ba47c2d7cad5d335dcb6e3;
    inBuf[618] = 256'hbfea1cf135f7eefd1f05e70ccb15561f4c29ef33a73e17496353d25cd4646d6b;
    inBuf[619] = 256'hf96ff371a4710e6f2e6ab663425c2454e94b2e443c3d39376832d62e282c0c2a;
    inBuf[620] = 256'h402828264f23da1fd91b73177a137510690ebf0d750ec20f79116513a8144d15;
    inBuf[621] = 256'hac152e15ee136f120b109c0cb508ee0340fe8af8dff27bed45e956e6aae4aee4;
    inBuf[622] = 256'h1ce69ee847ecadf06cf573fa5dffdf03e807570b5a0e4a116a143318da1c3622;
    inBuf[623] = 256'h3328532ec7331e38df3a8f3b553a7d373d33142e7d28b722021d7e173612350d;
    inBuf[624] = 256'h7508fa03ceffe0fb24f890f403f166edc1e927e6c0e2c1df58dd9bdb9fda6eda;
    inBuf[625] = 256'h01db70dce0de40e292e6c9eb5df1cff6d7fbddff97024b040305f804dd04eb04;
    inBuf[626] = 256'h34051d0695075209700bb00da80f47114a12491258118f0ff10ce909fc067104;
    inBuf[627] = 256'h9902ba01c1016c0296030d058606fa078c09350bf60cda0ead102d124613ed13;
    inBuf[628] = 256'h28144814a5145d157e16f1174a192e1a6d1ad11957183e1691135110af0c9808;
    inBuf[629] = 256'hfd0339ff99fa6ef648f36cf1d8f084f10df3f6f4f7f6c6f85cfa02fcdbfd1900;
    inBuf[630] = 256'hf30231069609fe0c1c10e2127915ec17721a3c1d1420b622c524b82548257423;
    inBuf[631] = 256'h6720981c8918a7143b113f0ea50b6009340726056f03f901cf00030019ffcafd;
    inBuf[632] = 256'hf6fb78f9a4f617f442f26cf1dff160f367f58df74af926fa20fa63f91ff8b4f6;
    inBuf[633] = 256'h63f524f4d2f249f162ef0ced76ea05e802e693e4e6e3dee314e45ae48de48ae4;
    inBuf[634] = 256'h9ce414e5f7e56ee777e98eeb83ed49ef9af0aff1f4f26df456f6def884fbf3fd;
    inBuf[635] = 256'he0ffa3001a0073feaefb42f8bff43af1faed0deb05e8e7e4b1e12ddec9dae2d7;
    inBuf[636] = 256'h63d59cd38ed2aad1e4d029d031cf71ce61ce12cfe7d0e7d383d773db5adfbee2;
    inBuf[637] = 256'hb1e554e8a8eaf5ec39ef2ff1bff29df38df3cbf27cf1dcef7dee82edd3ec8cec;
    inBuf[638] = 256'h5eecccebd8ea68e95fe73ee553e39ae172e0dedf6cdf30df23dfe9ded4de37df;
    inBuf[639] = 256'he0df0de1d5e2aee47de62be83fe9dde948ea5aea66ea9feab6eabdeaacea2dea;
    inBuf[640] = 256'h7ce9bde8cde713e7a3e631e6f5e5bae509e52ae41fe3c0e1b8e04de04ee028e1;
    inBuf[641] = 256'hb8e255e416e6d9e729e964eacaeb14ed7eee0df039f1e3f1fcf138f1c2ef01ee;
    inBuf[642] = 256'h23ec6aea1de92be862e7a4e6c1e567e47de216e018dd8fd9e2d52ed26cce08cb;
    inBuf[643] = 256'h24c882c570c329c25ac121c1b0c185c281c3dbc432c69cc7aec94dcc96cf1bd4;
    inBuf[644] = 256'h7cd953dfe6e5deecf2f3d5fbe4043b0f5f1b3529fc37f546f954c0606a69476e;
    inBuf[645] = 256'h266f756cdd66625f10579f4eae466a3f8738c1318a2a1c2228185e0c90fe50ef;
    inBuf[646] = 256'h4edf66cffcc032b5deaccca8fba8efacf6b3c7bc55c607d00dd961e18ce96ef1;
    inBuf[647] = 256'h4af9bf01690a0613e41b87249e2c8e34303c53434f4ad5505456b05a7b5d205e;
    inBuf[648] = 256'hb65c74595454ba4d6746b13eef36fa2f452acc25f922ed21ef218c2261236323;
    inBuf[649] = 256'h0822871fe31b8717831357101f0e2c0d300d5a0d5d0dee0c700b02090f067402;
    inBuf[650] = 256'h6afe72fa3df698f1d8ecd0e76fe253ddc2d8e7d452d23bd1a7d1c5d376d786dc;
    inBuf[651] = 256'hd7e206eabbf1a5f93b011e08150eed12de164a1a8a1d1c2132259729102e0a32;
    inBuf[652] = 256'hc834da35f334fd31512d562791208e199412f30bd5051200cefa29f6e7f124ee;
    inBuf[653] = 256'h0beb56e8f7e508e44ae2a2e034df06de24ddbfdcf1dca8ddd9de8ce094e2ebe4;
    inBuf[654] = 256'hd5e739ebf6ee3df3abf7a6fb2affd00117036003e602b1018400daffadff6300;
    inBuf[655] = 256'h14024804e906c9096b0cb50ea4100e1200139613d313cc13b613d5136d14c815;
    inBuf[656] = 256'h1a183e1bd71e72225b25f026fd266f257222a31e8c1a8c1602130010640d2b0b;
    inBuf[657] = 256'h43099c075d068b05f1047304d903d0024a0177ff84fdd6fbf1fa1afb7bfc1bff;
    inBuf[658] = 256'ha002a406da0adb0e8312fd155019861cc71fdf2273255f2773289228f027eb26;
    inBuf[659] = 256'hdb25fd2472241f24a923c3224f212d1f741c74194c161113de0f910c2909bd05;
    inBuf[660] = 256'h7d02a6ffa0fdb2fcd2fc14fe1200370233049e052f062006a805ed0453040204;
    inBuf[661] = 256'hd803d203d703b4037f0360035c0396030a0467045d04ae032102c4ffe0fcdef9;
    inBuf[662] = 256'h33f72df5f9f39bf3d4f376f465f56af67bf7b8f801fa46fb81fc61fdb7fd85fd;
    inBuf[663] = 256'hb2fc71fb2cfa09f93ff801f80ff82cf82bf8a7f77cf6d3f4c5f299f0a6eefdec;
    inBuf[664] = 256'h98eb5deaffe867e7abe5e3e36ae2a0e18ce12de268e3d0e422e653e73ce8fae8;
    inBuf[665] = 256'hd6e9d1eaf5eb54eda9eed2efe9f0d9f1cdf220f4d0f5daf735fa75fc3afe3cff;
    inBuf[666] = 256'h29ff05fe0bfc8bf910f7fcf47bf3b1f25bf223f2f4f18ef1e6f055f0e3efa4ef;
    inBuf[667] = 256'hceef13f037f044f0f3ef56efdfeea9eee8eedbef3bf1ccf260f4a0f588f62df7;
    inBuf[668] = 256'h9cf72df8eaf8c3f9b9fa8dfbf9fb04fca9fb0afb7efa3ffa78fa2cfb2efc47fd;
    inBuf[669] = 256'h15fe68fe4cfe9efda3fcbefbcbfafef981f9dcf838f8cdf746f708f75bf7c9f7;
    inBuf[670] = 256'h7cf85df9c5f9dff9a0f9c2f8d0f7f1f611f6b4f5b4f5b8f5eaf5e1f555f587f4;
    inBuf[671] = 256'h5af3f5f1baf0a7efeeee8dee36eeeeed62ed60ec55eb14eab8e8e9e733e75ae6;
    inBuf[672] = 256'hdde524e5ebe3efe2f8e1e3e05ae02ae0f2df01e032e030e03ee0aae057e165e2;
    inBuf[673] = 256'h4ee4d2e68ae9f1ece3f0f2f40cfaa1006e0854127e1ef22b643ae848cc554460;
    inBuf[674] = 256'h8d67116b416b9c68f063465e0c58df51024cf745d53f4e3984319f28671e4112;
    inBuf[675] = 256'he704c4f611e853da8dce59c5e9bf60be55c086c5b7ccefd4a4ddc2e53ced77f4;
    inBuf[676] = 256'h1dfbbb01e30812105f17df1edf25692cac327638103ea74306490a4e6052b655;
    inBuf[677] = 256'hb2570e58fe5675547050a04b2446fe3f083a8e349a2ff62bcd29cb28ec28b129;
    inBuf[678] = 256'h542a5a2a682973278324fa20941d681aa917d11538146e12aa101d0e9a0aea06;
    inBuf[679] = 256'hb00214fef0f9b8f542f116edade809e4d3dff8dbdad805d763d63cd79fd940dd;
    inBuf[680] = 256'h4ce292e8b2efc4f74600a408b310d117a81d6d220726be281b2b372d502f7231;
    inBuf[681] = 256'h3d337634a33441334e30ae2b9725bf1e76172b107309390381fd82f80af426f0;
    inBuf[682] = 256'h16ede0ea8ee906e911e97ee9e9e936ea8ceacbea30eb12ec25ed59eebbefcaf0;
    inBuf[683] = 256'h6ff1e9f116f22bf2a6f285f3b1f43ff6f2f748f91bfa70fa17fa4ff9bdf878f8;
    inBuf[684] = 256'haff8d5f9a2fbbefd66004b0323064809970ccc0f0413e8150e187319031ade19;
    inBuf[685] = 256'h76191a192019ad19941aaa1b841ca91c001c611ac5178d14ea10030d29095705;
    inBuf[686] = 256'h7901a2fdcff925f6e8f23ff065ee66ed0ded4aede0ed8fee6def8af0f7f1f4f3;
    inBuf[687] = 256'h92f6c8f983fd77017e0583095b0d2011dd146818c11ba81ebc20f4211d220221;
    inBuf[688] = 256'hf61e181c7a18b114fd10650d3f0a91071505dc02d900ddfe05fd64fbd6f963f8;
    inBuf[689] = 256'h0ff7b3f54ef40ff305f25df165f113f240f3ddf47af6b0f77ff8ccf89af842f8;
    inBuf[690] = 256'hd6f754f7d7f628f62df5faf367f2a0f0edee39edceebe5ea3deaf0e902eafee9;
    inBuf[691] = 256'hfce908eacfe9a2e9bbe9dde95cea5ceb6decaded20ef59f07af1abf2a5f378f4;
    inBuf[692] = 256'h12f50ef567f41df30ef18beee2eb25e9a6e682e46ce26fe07bde3fdce9d9b5d7;
    inBuf[693] = 256'h89d5b2d36cd266d1afd04cd0d3cf65cf42cf35cf8ccf92d0edd1a7d3cbd5c8d7;
    inBuf[694] = 256'h9ed967dbcedc16de79dfa9e0d7e1f9e293e3dae3e2e370e313e308e30fe38de3;
    inBuf[695] = 256'h6ee422e5e1e590e6c5e6f0e622e715e733e76fe761e750e71ae762e686e586e4;
    inBuf[696] = 256'h34e3fde1efe0e0df21df9dde11deb1dd6cdd1cdd12dd58ddcadd99dea6df9ce0;
    inBuf[697] = 256'h8fe175e21fe3d4e3cde4ece567e74ce943eb49ed54ef0af177f2a3f33cf461f4;
    inBuf[698] = 256'h23f447f31ef2e0f06bef24ee32ed4becb6eb72eb1debf6eaebea97ea44eadde9;
    inBuf[699] = 256'h0fe946e88ae7a2e610e6e6e5e4e56fe687e7d9e899eaaaeca6ee8ff030f237f3;
    inBuf[700] = 256'hb1f39ef3faf2faf1bff059efdced56ecd7ea5be9f0e7b4e67fe53ae4f4e268e1;
    inBuf[701] = 256'h6cdf35ddbcda03d87cd569d3d3d108d131d110d293d3b2d50dd880da26ddc6df;
    inBuf[702] = 256'h4fe210e5d8e77eea71edaef036f4cff8dcfe710609107f1b0a280f3585413b4c;
    inBuf[703] = 256'h7d54b459a05b955afe568f51254b4e44aa3d9037d231642ceb26b42085190f11;
    inBuf[704] = 256'hff06bbfbaaef4be3c5d7f0cd7ac644c26ac1a0c399c84bcfcdd69cdedde569ec;
    inBuf[705] = 256'ha8f262f8dafda3035409ce0e6914bb19ae1eb823af288a2d9e32af377f3c2741;
    inBuf[706] = 256'h5f45bf482f4b774c3d4c764a64473f43603e76390f356431c92e6f2d052d452d;
    inBuf[707] = 256'h012eb12ed72e5a2e022d902a4e278f23471fd21a97164312da0da40937059b00;
    inBuf[708] = 256'h5bfc3ef857f42ff15deeafeb7be94ee700e508e334e1a1dfefde15df57e041e3;
    inBuf[709] = 256'h9ee772eddff43afd1106210f8717c71ec2241229c02b372da62d672df02c6c2c;
    inBuf[710] = 256'he42b552b9f2a8229c4276d258022fa1e2e1b55176e13c90f9c0cca098107de05;
    inBuf[711] = 256'ha904dd039e03ca0343042805610681076b081809160950081d074705d3024400;
    inBuf[712] = 256'h59fd09faf9f60bf445f157ef2bee8cedceed77eef0ee65ef9aef70ef72efc6ef;
    inBuf[713] = 256'h89f038f2e0f4a6f8ecfd9204750c7715e01e022863304737443c5c3f88400140;
    inBuf[714] = 256'h433ea53b7e3838351c325c2f142d362b7b297827d1244a21e51cf317fb127b0e;
    inBuf[715] = 256'hd60a5108ef067c06d406d00711097c0a130c740d800e600fb40f600fce0ed20d;
    inBuf[716] = 256'h6b0c1c0bbc092908cf06930577040c0454044e054d070c0a3a0dca103e143617;
    inBuf[717] = 256'h9919221be71b331c241c2c1c901c431d831e3e201a221824ef252827d427d027;
    inBuf[718] = 256'hf2269125bd236321d21efd1bcd1889151f128c0e1f0bcd078d04a601fbfe71fc;
    inBuf[719] = 256'h3dfa5af8c1f6a8f5fbf481f41bf48ef3aef2a6f1c1f03ef077f0a1f194f311f6;
    inBuf[720] = 256'hdcf886fbb5fd4eff34005c00efff1bff06fee5fcf2fb5afb23fb51fbddfb79fc;
    inBuf[721] = 256'hf2fc51fd65fd34fd0bfdd1fc7cfc47fcfbfb8afb43fbf9fa94fa43faadf992f8;
    inBuf[722] = 256'h20f72ef5cbf25af0e7ed8eeb6fe94fe71fe5d3e23fe0aadd55db4ed9ffd789d7;
    inBuf[723] = 256'hbcd7bad85fda53dca6de21e171e3b6e5cee791e951eb1aede3eefdf060f3e2f5;
    inBuf[724] = 256'h95f83bfb85fd64ff9700fc00bf00e1ff89fe12fd8dfb05faadf869f70cf6b0f4;
    inBuf[725] = 256'h49f3b9f135f0d2ee71ed2cec08ebcce995e884e779e6ade550e533e575e529e6;
    inBuf[726] = 256'h03e70de850e982eab5ebfbec1fee44ef6ff063f136f2c7f2d4f296f20bf225f1;
    inBuf[727] = 256'h65f0dcef6aef64ef9eefbdeffdef43f068f0dcf09df188f2dff360f5aaf6dbf7;
    inBuf[728] = 256'hc1f822f956f982f9a3f905fac7fab3fba6fc73fdbdfd3cfde7fbc8f9faf6e2f3;
    inBuf[729] = 256'hdbf003ee8eeb85e99ce7c6e513e44ee29de04fdf2ede1ddd3ddc34dbb9d90cd8;
    inBuf[730] = 256'h3fd64ed4aad2a5d12ad168d180d223d44ad616d93ddcc0dfe5e363e820ed5ef2;
    inBuf[731] = 256'hcef747fd2d0388097d10aa184522492da739aa464653615eb066526be86b7468;
    inBuf[732] = 256'hb661b8586f4e04443c3a4b315e293722431b2d147d0cd7034cfae5eff7e44cda;
    inBuf[733] = 256'h7ad050c8c9c248c019c158c542cc23d542df47e989f2edfae0019907ef0cd211;
    inBuf[734] = 256'h67163e1bec1f0024be27e62a422d562f55312d3335357d37a2398a3b253d123e;
    inBuf[735] = 256'h2c3eb13da33c083b5139d0378136bb35d4358e36ce37a5398a3bef3cc43da33d;
    inBuf[736] = 256'h0e3c42396a356730b22aaf24281e371700102208b4ff2af799ee7ee685dfbcd9;
    inBuf[737] = 256'h46d552d276d079cf5ecfcdcfccd095d208d553d8b1dce7e111e850ef3ef7c8ff;
    inBuf[738] = 256'hde08cc11281ab821cd270d2c9c2e612f7a2e6a2c972937269822f51e311b2017;
    inBuf[739] = 256'hd412470e6909a40450007bfc89f9aaf782f615f666f6f0f6b0f7e6f843fabefb;
    inBuf[740] = 256'h9bfd97ff660114037104230520056b04d8025f0033fd5bf9d7f4f4efdceaa0e5;
    inBuf[741] = 256'hade057dcb4d828d6e2d4abd484d55ad7c0d9a0dc03e0b9e3d5e77eec9cf128f7;
    inBuf[742] = 256'h08fdfe02e4087a0e8313f217981b4a1e242030216e212a219a20c31fcb1ebf1d;
    inBuf[743] = 256'h751cd31ad018471627138a0f800b2407bf028ffec0faa0f764f503f48cf3f5f3;
    inBuf[744] = 256'heef443f6d9f76bf9cffa16fc46fd5dfe7fffd60061021204f105e007a409320b;
    inBuf[745] = 256'h7d0c670d070e6e0e980ea30e960e490ec70d0c0df30b980a2709b20765067605;
    inBuf[746] = 256'hf904ec043f05ea05c00692075d080b097509ac099a090e091e08c106eb04f302;
    inBuf[747] = 256'hfc0012ff7ffd2ffcecfacaf99bf836f7d7f57cf421f303f20bf128f07cefe5ee;
    inBuf[748] = 256'h78ee6eeeacee4bef6bf0bdf130f3c9f43cf690f7dcf8eaf9d7faa7fb20fc6bfc;
    inBuf[749] = 256'h9bfc85fc65fc53fc14fccdfb7ffbebfa3dfa7df981f87df774f62df5d4f36ef2;
    inBuf[750] = 256'hcaf023ef92ede2eb3aeaaae8f1e631e596e3fee194e08edfb5de0ade9edd27dd;
    inBuf[751] = 256'ha3dc37dcbbdb4edb1fdbfadaeada05db07db09db2ddb41db70dbc4dbeddb0fdc;
    inBuf[752] = 256'h2ddcffdbe0db06dc3ddcf0dc3bdeb1df84e1a5e39ae59de7b0e973eb28edcaee;
    inBuf[753] = 256'hf5efeaf0b0f108f252f29ef2b4f2c8f2b0f209f2f7f05bef12ed87eae0e719e5;
    inBuf[754] = 256'h98e25de031de4edcb2da36d92dd8bbd7bfd770d8e0d9c8db2ede16e12ae459e7;
    inBuf[755] = 256'h98ea8bed1bf03ff2b3f38ff4f5f4caf44ff4b1f3c3f2bff1bcf07bef44ee30ed;
    inBuf[756] = 256'hf7ebe5ea05eaf7e817e888e7f6e6d6e652e701e82ee9e1ea8fec66ee66f01bf2;
    inBuf[757] = 256'hb5f33cf553f628f7bcf7c1f76ff7d5f6c7f58ef44af3e6f1a5f0a8efd5ee43ee;
    inBuf[758] = 256'heaed8ded0ced56ec54eb10eac1e893e798e6fce5bee596e579e562e50ce590e4;
    inBuf[759] = 256'h42e4fde3bae3b2e39ee326e374e28de14ee011df2ede8bdd4fddb6dd6dde5ddf;
    inBuf[760] = 256'hbae029e286e32ee5efe6ade808eb2aee34f2fef7ebfffb096816cb243334b443;
    inBuf[761] = 256'h0a52ee5d7666ec6a346bc467516117594850ab47024063393b33212d4826d81d;
    inBuf[762] = 256'hbf13f707c6fa3bed2de06cd424cbcac4a9c124c2c1c5fccb70d4dfdd7ce7f6f0;
    inBuf[763] = 256'h56f97300e306610c2b111316c31afc1e16238426df28a12acd2b802c842d1b2f;
    inBuf[764] = 256'h2931e0330537e9393a3ccf3d573ee23dfd3c153c783b9f3bbd3c883eb8401443;
    inBuf[765] = 256'h1e457046fd46a4463445de42c93fd43b3a374332ca2cff263221141b9814e90d;
    inBuf[766] = 256'h9a06b7fedcf620ef14e8aae2ecdef9dc08dd52de53e0e9e250e57ce7f2e988ec;
    inBuf[767] = 256'ha2efe8f3ebf888feea044b0b4f1119171e1c21205b237c256326602668258023;
    inBuf[768] = 256'h01211a1ede1a7c172f14fe10dc0d0b0bbf08f10601064d06b707570a3e0edf12;
    inBuf[769] = 256'hc917b01cdd20ce238225e125e924062391208a1d131a6e167112030e67098c04;
    inBuf[770] = 256'h4affe6f962f49eeef6e89ce3afdec0da27d801d78ed7a6d9eedc25e1dce5e5ea;
    inBuf[771] = 256'h60f037f6b0fc2c04610c2b156e1e3b27df2e203548391f3b303ba239bd364233;
    inBuf[772] = 256'h5f2f0b2b972602221e1d1e181e13120e160941048cff06fbe3f67df343f1b5f0;
    inBuf[773] = 256'h57f253f66dfc3b04f90c96155e1dd4237a286a2b1e2db12d692dba2c712b4f29;
    inBuf[774] = 256'h8826f6228d1ee0193d15cf100d0d080a9107b70559045803e202170323043606;
    inBuf[775] = 256'h3d09240da6113716a81ac51e2222ec244e27ef28e7294f2a9c29b827d924cf20;
    inBuf[776] = 256'he91bcf16c411280d56092906720301018afe09fc97f962f7c7f5f3f4eff4dbf5;
    inBuf[777] = 256'h81f79bf931fc17ff120241057f08710bfd0def0ffa102b11ac109a0f370eb90c;
    inBuf[778] = 256'h300b9609d007c70562038d0074fd46fa24f76df462f2f8f04ff067f0e1f0a7f1;
    inBuf[779] = 256'hc1f2dcf3fcf460f6def76bf939fb0cfda7fe1f004701ec012502dd01ec0051ff;
    inBuf[780] = 256'hfafce6f93df631f216ee3beac4e6dde37fe160df75ddaadbd3d93bd838d7d6d6;
    inBuf[781] = 256'h6ad727d9b8dbfcded3e2c7e6b5eaa8ee71f218f6a5f9e2fcbaff06028a035204;
    inBuf[782] = 256'h58048f033b026300f5fd2efb0cf87cf4dbf04eede2e906e7dbe443e382e282e2;
    inBuf[783] = 256'hece2e0e34ae5d0e69de8c9ea0ced7fef2ff2b4f4e6f6b3f8caf92afa0cfa8df9;
    inBuf[784] = 256'he9f862f8fef7b1f74cf773f613f52bf3bcf02beec6eb95e9e2e7aee6aae5f0e4;
    inBuf[785] = 256'h87e435e443e4dde4cae537e728e940eb95ed29f0aef240f5cef7faf9c6fb05fd;
    inBuf[786] = 256'h68fd23fd44fcc6fa2af99df70ef6daf4e5f3cef2b2f166f099ee9aec94ea87e8;
    inBuf[787] = 256'he8e6ebe56be57fe507e697e61ae784e7aae7b0e7d4e70ee867e8fae89ee914ea;
    inBuf[788] = 256'h64ea88ea43eaa6e9e8e8cce735e666e43ee28ddfc6dc2adaabd7bcd5a4d41bd4;
    inBuf[789] = 256'h2cd4e6d4d7d5f1d66cd802dab3dbd5dd20e06ce212e513e88feb4bf0d0f679ff;
    inBuf[790] = 256'hb70a6d18f42760384a4844560c618c676169d26679609957a94dcb430d3bfd33;
    inBuf[791] = 256'h652edc29a525c220961ab512fb08e4fd08f239e6aadb39d3a7cdb3cb53cd30d2;
    inBuf[792] = 256'hc1d9bce212ec0ff5a5fca0028b07400b1f0e0e11cd132c16a818de1a831c251e;
    inBuf[793] = 256'hc41f582171230b26ec28422cce2f153304366e38f6398d3a663aa53977385137;
    inBuf[794] = 256'haa368a3609374b38e1395b3b943c073d503c943ac337e933932f052b5e260422;
    inBuf[795] = 256'hf61de719c6154611ff0b06067aff75f896f161ebf9e5c1e1d7ded5dca0db22db;
    inBuf[796] = 256'hf7da33db14dc71dd75df52e2a8e55fe98dedbff1cff5ebf9b5fde9009f038e05;
    inBuf[797] = 256'h8406c4067406bf050d059504560441043304e5031103bc01050004fe24fcecfa;
    inBuf[798] = 256'h84fa2ffb24fd0a008f036f07fd0ace0dc70f9b104110050fe50cf90988069b02;
    inBuf[799] = 256'h4afed1f955f5f6f0c8ecc2e8dee401e126dd7bd934d6a6d33cd221d268d305d6;
    inBuf[800] = 256'h97d9bfdd37e2a6e6f6ea40ef90f31df80dfd4202ac070f0de711f215ef18861a;
    inBuf[801] = 256'hd11a021a2b18b115f21201101f0d820a0e08db05090471020301c2ff89fe49fd;
    inBuf[802] = 256'h17fc0dfb57fa2bfab8fa10fc14fe99005e03f5051408a2096f0a8d0a4f0ad109;
    inBuf[803] = 256'h3209bf086b0804089e071a073d062e050e04d402b301e1005a00360096007101;
    inBuf[804] = 256'hb3027704a6060409810bf80d1a10cd111513d3130f140014a51302133a122a11;
    inBuf[805] = 256'hb30fe00d920bd108de05ca02bcffecfc3bfaa4f73bf5cef276f074eeb6ec6beb;
    inBuf[806] = 256'hd1eaa4ead1ea5bebd7eb3cecc5ec51ed0dee3fefb4f05cf225f4a9f5d9f6b3f7;
    inBuf[807] = 256'h02f8f8f7b5f718f767f6b4f5bef4d0f3f2f2daf1d7f0faeff4ee21ee9fed1bed;
    inBuf[808] = 256'he3ec0eed21ed43ed85ed7aed5eed6eed61ed63ed9bedb0eda0ed7eed10ed69ec;
    inBuf[809] = 256'ha9ebb9eab3e995e83ee7b9e5f8e3ede1d2dfb1dd8cdbaad911d8b3d6c9d549d5;
    inBuf[810] = 256'h17d560d507d6d6d6edd728d953daaadb1cdd81de20e0f1e1b2e39ae59be762e9;
    inBuf[811] = 256'h0ceb91eca7ed79ee19ef5aef76ef81ef4def12efdfee7dee34ee16eed7ede0ed;
    inBuf[812] = 256'h12ee18ee45ee68ee49ee0deec6ed44edc4ec70ec21ecf8eb10ec2eec58ec94ec;
    inBuf[813] = 256'hb7ecd0ece8ecf3ec16ed58ed9dedf9ed55ee7cee7aee59ee06eeb0ed7eed57ed;
    inBuf[814] = 256'h53ed7aed84ed5eed16ed7deca6ebdeea31ead5e913ead1ea03ec99ed38efc0f0;
    inBuf[815] = 256'h22f22bf306f4cbf467f515f6bcf611f745f727f77cf6baf5d7f4a8f3b3f2d5f1;
    inBuf[816] = 256'haff0b0efb9ee7fed8fecf4eb69eb50eb9debeceb56ecc8ec04ed16ed17ed15ed;
    inBuf[817] = 256'h21ed5eedf2edb7ee9cefa3f04ef165f11af123f0a1ee4bed1cec19ebafea81ea;
    inBuf[818] = 256'h0aea50e911e823e6e5e3aae1aadf3ede89dd76dde6ddb1de8fdf56e024e1f5e1;
    inBuf[819] = 256'hcfe228e450e685e980eec5f57fffe30baa1a072beb3bd24b5c595c63c3689269;
    inBuf[820] = 256'h33664f5f6d56f24ccd43f73bce35d6309c2c5c280a23431cd313cb0902ff40f4;
    inBuf[821] = 256'h74eadae2f7dd38dc02deb9e2d7e9eff296fcf305bb0ec815d41a7b1e6c20ef20;
    inBuf[822] = 256'h1e21ea205b202320fe1fa11f791f7a1f921f3520802147238a252128972aa72c;
    inBuf[823] = 256'h602eb72fa4309f31f53287349f367639a03cfd3f9343d4465949184bba4bf64a;
    inBuf[824] = 256'h0049034608426c3d8f387733502e50293a24f91eae1909140c0e18080f0238fc;
    inBuf[825] = 256'h33f7e7f276ef43edceebe7eac5eadcea32eb48ecc9ede1ef09f39af658fa6bfe;
    inBuf[826] = 256'hfd01be0401076508f1082e09090997083808ea07b707b407ef077a082f090e0a;
    inBuf[827] = 256'h220b010cac0c620dc60d0a0ebe0eb40f15114913e615b818ae1b2e1efe1fe820;
    inBuf[828] = 256'hbe208f1f621d6f1ae616f012b10e760a3f061d025afee2faadf7e8f46cf23ff0;
    inBuf[829] = 256'h8eee52edcbec1bed29ee31f006f343f6fbf9cffd4f01bd04e5079b0a740d5910;
    inBuf[830] = 256'h1313131602195d1b5f1db51ef31e751e3e1d371be418891643146f123811a810;
    inBuf[831] = 256'hd0109211ca123f14a615e116cf175518be185719501a1e1c181f1d230228712d;
    inBuf[832] = 256'h9332a33626398a399e37d933ac2e9f289422ff1c0218e2138310940d160bea08;
    inBuf[833] = 256'hfe06780549047a0334035603fb0364057d076f0a610ef812ff17251dab214025;
    inBuf[834] = 256'hb327a0284028f526bd24eb21c31e201b1c17ca12140e4509b4049e0078fd83fb;
    inBuf[835] = 256'hbdfa36fbaffccdfe5e01fd03620698087b0af60b3a0d2c0ead0ee70ec80e260e;
    inBuf[836] = 256'h510d370c930a8e080f06ea0240ff27fbbbf64ef227ee8aeabde7d3e5cce487e4;
    inBuf[837] = 256'hb2e42ce5e7e5b9e6b4e700e98fea6beca2ee08f17ef3e8f50bf8d1f935fb0efc;
    inBuf[838] = 256'h57fc27fc81fb87fa5df90af8adf652f5eaf389f234f1dbefa3ee94ed8feca7eb;
    inBuf[839] = 256'hdaeaf6e91de96de8d5e78ee7b7e721e8d2e8b8e985ea38ebc9eb0cec36ec65ec;
    inBuf[840] = 256'h7deca6ecdfeceaece7ecd7ec96ec65ec56ec47ec6fecbbeceaec1fed45ed24ed;
    inBuf[841] = 256'h02ede7ecbbecccec13ed57edc8ed4bee97eee6ee3aef5bef87efcdeff6ef2ef0;
    inBuf[842] = 256'h77f095f0b0f0d5f0cdf0c2f0d0f0c7f0caf0f6f01bf151f1adf1eff11ef242f2;
    inBuf[843] = 256'h16f2abf115f119f0e3ee9eed1cec92ea38e9dee7b3e6e2e522e597e460e42ce4;
    inBuf[844] = 256'h21e45ce491e4e4e464e5c5e537e6bfe60be75de7c9e705e852e8b4e8d5e8f9e8;
    inBuf[845] = 256'h20e9ffe8dfe8bfe85de80ee8d7e772e741e74de758e7bde782e852e95cea8feb;
    inBuf[846] = 256'h8dec74ed43eeb1eedfeee4ee9aee21ee9aedeeec20ec40eb36eae6e85ae79de5;
    inBuf[847] = 256'h9fe37ce17cdf9ddddfdb95dabfd91cd9d1d8dcd8ddd8ead825d94bd971d9d2d9;
    inBuf[848] = 256'h3ddabfda99db97dcb2dd31dfefe0f4e2b7e55fe914ee50f43efcd6050d11761d;
    inBuf[849] = 256'h6f2a2e379e42e24b445221558454e950d74a5a43963b2f34c62da22861249620;
    inBuf[850] = 256'hbe1c1e185e12720b860340fb5df3a6ecf8e7cfe57ae60feaf9ef9ef75300d908;
    inBuf[851] = 256'h60108316751a261c2d1c8f1acd17ed141512770fac0d840ccd0bc10b1c0cb70c;
    inBuf[852] = 256'he10d750f45117b13f1157e18311bfb1dd520cd23f126592af22d9d315e35e238;
    inBuf[853] = 256'hc53bf23d223f0b3fd33d863b28381734892f982a93259520981bbe16f211150d;
    inBuf[854] = 256'h4b08790389fec3f938f5f1f04fed64ea20e8c4e636e622e69de678e74ae83be9;
    inBuf[855] = 256'h4dea24ebf6ebf8ecdcedadee93ef3af08bf0a5f05ef0b5efe6ee0eee49edbbec;
    inBuf[856] = 256'h70ec62ec85ecd7ec4eedd1ed76ee4def39f05cf1d7f290f4a4f635f91afc50ff;
    inBuf[857] = 256'hd00247068609590c630e7f0f970f920e9e0ce5099006020370fff6fbd2f8f5f5;
    inBuf[858] = 256'h45f3dff0aaee97ecdeea82e994e850e8b7e8cbe9a6eb23ee2ef1bcf47ff845fc;
    inBuf[859] = 256'he0fff802720543074f08d208f408b7085d08020887071507b1062e06af053b05;
    inBuf[860] = 256'hc20466042604f90309046204fc04ec052c079d082b0aae0b0e0d460e3d0f0510;
    inBuf[861] = 256'hbf1061110112ae123e139e13c1137713bb12a21133109c0e110dad0b8f0acb09;
    inBuf[862] = 256'h580935095909c1096f0a500b5f0c9a0ddc0e1210471170128f13bf14f9152c17;
    inBuf[863] = 256'h4d183519be19c9192a19dd17f8158913b710bb0db10abc07ff0474021e0006fe;
    inBuf[864] = 256'h1bfc5afacbf85ff71af611f53af495f32bf3f1f2e1f208f35bf3ccf34ff4c5f4;
    inBuf[865] = 256'h1ff55cf571f569f55af549f537f525f504f5d5f4a1f462f41af4dbf3adf398f3;
    inBuf[866] = 256'h97f3a2f3b7f3d3f3eff3fff3f5f3cff397f348f3e8f28cf241f20cf2f4f1f3f1;
    inBuf[867] = 256'hfef10bf20cf2fbf1dff1bcf19af182f178f178f175f161f139f101f1bdf06bf0;
    inBuf[868] = 256'h23f0eaefabef6def22efb5ee1cee60ed88eca4ebcbea08ea6be9fee8b3e88de8;
    inBuf[869] = 256'h8ee8afe8fee886e933ea04ebfbebf2ece2edd5eebbefa1f0a7f1c8f20df47df5;
    inBuf[870] = 256'he8f639f863f93efacffa38fb79fbacfbeefb2ffc73fcb9fce0fce6fcd2fc8bfc;
    inBuf[871] = 256'h28fcc0fb3ffbb5fa2dfa8bf9e6f852f8bef740f7e2f688f647f62cf619f628f6;
    inBuf[872] = 256'h73f6d4f658f711f8d0f895f965fa15fbabfb32fc7dfc8ffc74fc06fc5bfb96fa;
    inBuf[873] = 256'ha5f9a1f8a7f792f66ff549f4fbf2a7f173f04def6deef6edc1ede8ed6dee09ef;
    inBuf[874] = 256'hccefb2f073f126f2cdf220f34cf363f328f3ddf2acf260f238f25cf28cf2ecf2;
    inBuf[875] = 256'h87f3fff355f482f42cf463f34af2d3f04aef02ee04ed87eca6ec31ed05eef8ee;
    inBuf[876] = 256'hb6ef0ff0e8ef37ef0eee7eecc4ea0be954e7e1e5d3e4fae37ce362e34be346e3;
    inBuf[877] = 256'h51e317e3c3e279e201e2aae1afe1cce145e25de3cae4c8e6b3e970ed3cf26ff8;
    inBuf[878] = 256'he8ffab08b6128a1dbf28d033c83def45bd4b844e2d4e1e4bc145f43ec737eb30;
    inBuf[879] = 256'hf82a4726a522c31f2d1d571afd16f6123f0e43095e040f001efde2fba8fcd0ff;
    inBuf[880] = 256'hde04480baf12cd19b51f38246a260f26f8231320c91a84157610ec0b01098707;
    inBuf[881] = 256'h3c07a0081e0b2b0e09121f16031a0c1edb214225ad28f32b112f6032bc352039;
    inBuf[882] = 256'h9b3cce3f8d42ac44b5459c456844ee416e3e3f3a83358c30b12b1427e7224c1f;
    inBuf[883] = 256'h461cdb19ee174b16de147913e1111710210ef50bc809cd0702069904af031403;
    inBuf[884] = 256'hc702d202da02d8020003cf025202db01e8007fff12fe3ffc17fa2cf845f673f4;
    inBuf[885] = 256'h3df37af21df273f244f35ef4d2f562f7e1f853faacfbe9fc13fe3aff6d00a601;
    inBuf[886] = 256'hf902840443064408980a230dc00f341234147815af15cb14ea121310af0c3609;
    inBuf[887] = 256'hcd05e002c60053ff9efea9fef9fe74ff0b005a00710073003f0024006100ec00;
    inBuf[888] = 256'h0802b603b8050908650a730c2d0e510fbd0fb40f2d0f3c0e420d400c300b4e0a;
    inBuf[889] = 256'h8309b208f7074a07a4062b06eb05f805630621072a087209dd0a510cb10ddf0e;
    inBuf[890] = 256'hcd0f6c10bc10d110bd109e109110ac10f6106211dc11491275124d12cf11f610;
    inBuf[891] = 256'he10fbf0eab0dda0c7d0c910c190d190e680fe5107112dc130415e7158816e516;
    inBuf[892] = 256'h1f174f177a17a717c617c2178a170f1745162d15d01329124610380efd0ba109;
    inBuf[893] = 256'h4207ee04bd02c30004ff8efd61fc6ffbc3fa68fa43fa48fa77faacfad2fae7fa;
    inBuf[894] = 256'hcffa88fa23fa8ff9d2f811f847f77cf6cff52bf58af4fff368f3b4f201f238f1;
    inBuf[895] = 256'h5cf09feff7ee79ee53ee66eea7ee2fefcfef7ef055f128f2f2f2bef352f4abf4;
    inBuf[896] = 256'hd8f4b9f471f427f4ccf392f389f380f38ef3aaf39af383f369f329f3f4f2c3f2;
    inBuf[897] = 256'h65f204f28ef1d5f013f04bef5eee8bedccecf3eb28eb66ea82e9b4e80fe87fe7;
    inBuf[898] = 256'h38e73ae74ee785e7d9e710e84ee8aee80ce986e92deac0ea45ebc8eb10ec34ec;
    inBuf[899] = 256'h5bec5bec52ec60ec54ec49ec5cec5fec7aecc9ec18ed86ed19ee8fee06ef7eef;
    inBuf[900] = 256'he3ef65f0e0f01bf14df179f16cf173f19bf1b6f105f285f2f6f287f32df4aff4;
    inBuf[901] = 256'h3cf5c5f512f647f658f61af6c5f569f5f8f4adf495f48ff4aef4e2f4f8f4fcf4;
    inBuf[902] = 256'he6f490f410f466f372f256f134f007ef0fee7fed3bed4fedb1ed02ee27ee16ee;
    inBuf[903] = 256'h96edcdecf7eb12eb64ea27ea35eaaeea99ebadecf7ed6befb9f0f1f101f3a1f3;
    inBuf[904] = 256'hfbf313f4c2f357f3eaf253f2ddf189f11af1c3f078f0fdef81ef03ef5beebeed;
    inBuf[905] = 256'h30ed98ec1fecc4eb70eb3eeb1eebfdeae7eac8ea9bea6cea25eacfe977e900e9;
    inBuf[906] = 256'h81e812e89ee745e725e71ee73de78be7dae72ce88fe8e6e840e9bee94deaffea;
    inBuf[907] = 256'hf7eb21ed95ee88f0fbf213f60afacefe5c04b60a84117f18691faf25e82ad42e;
    inBuf[908] = 256'h013156311030522d90297c257321dc1d111bf81867172d16d9142c130311430e;
    inBuf[909] = 256'h200bdf07d30486024b015e01ff02ef05ca09460e9e123516da180f1aad191818;
    inBuf[910] = 256'h5915b411df0d170ab00650040c03f6024f04c606ff09dc0dd1117c15d518951b;
    inBuf[911] = 256'had1d5c1f9c2088216e22472329243e255a2663275028ce28af28f02766261f24;
    inBuf[912] = 256'h5c213b1efb1aed172d15e1122911f50f440f0b0f0e0f300f480f0e0f780e880d;
    inBuf[913] = 256'h290c970a06096c070106da04b903b202cc01c400c1fff0fe20fe7afd28fde4fc;
    inBuf[914] = 256'hb4fcabfc7cfc28fcccfb3cfb93fa06fa8df94df96ef9cbf958fa02fb88fbd7fb;
    inBuf[915] = 256'hedfbc3fb7afb34fbfdfaecfa05fb3cfb99fb26fcebfcfbfd5fff0901d0028704;
    inBuf[916] = 256'hf705e3063107e7060406ac0418036301bdff62fe62fdd4fccefc2cfdc9fd8afe;
    inBuf[917] = 256'h2fff95ffc2ffb4ff89ff75ff98ff0c00de00ff015c03d8044b06a107ba087309;
    inBuf[918] = 256'hc0099909f208e8079f063405da03bb02df014e010501e100ce00c100a7008500;
    inBuf[919] = 256'h6e0069007e00b7000d017001d5012e027202940294027e0258022c0219022702;
    inBuf[920] = 256'h5302aa0219038303e5032a043c042c04ff03b20366032403ec02d602ed022d03;
    inBuf[921] = 256'ha4034f041b05f705cd068f073508c5085309e909860a300bd30b560cb50cda0c;
    inBuf[922] = 256'hbc0c6b0cda0b070b030ab9082a077805a003b701ebff36fe9ffc44fb08faeef8;
    inBuf[923] = 256'h17f86bf7eaf6aff68df669f650f617f6abf531f59cf4eef350f3c2f23ff2e4f1;
    inBuf[924] = 256'ha6f176f15cf143f119f1e2f094f031f0d3ef86ef5cef6aefa9ef1df0bdf070f1;
    inBuf[925] = 256'h3cf21df3fbf3e8f4ddf5b2f675f71df883f8c6f8f3f8f6f803f92bf950f995f9;
    inBuf[926] = 256'hf1f924fa3efa31fabef90cf92df8fef6c0f592f45bf352f284f1c2f02bf0bbef;
    inBuf[927] = 256'h38efc5ee66eef0ed8fed4ded04edd7ecc7ecb2ecb6ecd6ecfbec47edb6ed26ee;
    inBuf[928] = 256'ha9ee28ef74efa5efbaefacefb0efd9ef20f0aaf06df145f23ff341f41ff5eff5;
    inBuf[929] = 256'ha3f61bf785f7e8f731f893f816f994f92afacafa3afb95fbd9fbe1fbe6fbf8fb;
    inBuf[930] = 256'heefbf6fb0bfceefbbefb7ffbfafa5dfabaf9ebf822f87af7d5f666f642f63ef6;
    inBuf[931] = 256'h75f6e2f64af7bcf738f896f8f4f85cf9b2f90afa5ffa8cfaa3faa3fa77fa43fa;
    inBuf[932] = 256'h0cfabcf96df920f9baf85af810f8c4f792f77cf757f72ff703f7aff654f610f6;
    inBuf[933] = 256'hd3f5caf50df671f6fcf6a5f726f883f8bdf8b0f883f84df8fcf7bbf791f757f7;
    inBuf[934] = 256'h29f7fff6aff65ef613f6b5f574f553f533f52cf528f5fdf4b9f442f480f390f2;
    inBuf[935] = 256'h70f12df000eff6ed2eedd4ecd7ec3aedffede6eee1efdff09df11cf26ef270f2;
    inBuf[936] = 256'h4cf236f221f238f29ff232f3f6f3eaf4dbf5c7f6b9f79ef891f9b3fa02fc99fd;
    inBuf[937] = 256'h8dffd8018a04a107ff0a940e2d1281156918ac1a161cb81c9a1cc51b7f1aee18;
    inBuf[938] = 256'h1f174d158413b8110e10850e0a0dc80bbb0ad40947090e091c09a7099b0ae00b;
    inBuf[939] = 256'ha20db60ff6118a142b17a319101c1b1e8c1f98200321b9202220301ff41def1c;
    inBuf[940] = 256'h191c781b621b991bf01b861c001d341d541d301dd81ca41c791c701cc61c391d;
    inBuf[941] = 256'hca1d9b1e5d1f1c20ff20b9215422f522462353234b23ef225422bb21f4201520;
    inBuf[942] = 256'h571f821e981dba1c9f1b391aa918b5166e141a12ab0f560d720bee09e5088508;
    inBuf[943] = 256'h8908e808b309970a890bae0cb50da20ea60f7d102911e5116e12b912fc12ec12;
    inBuf[944] = 256'h7912d411bf103a0f8a0d930b72097c07a005f503b802c5011b01df00e3002601;
    inBuf[945] = 256'hc3018e028603c1040a065807b908f109ed0abc0b2d0c320ceb0b450b410a1609;
    inBuf[946] = 256'hc5075606f904b50385029401e80072004f007500c1003d01e3019c028603aa04;
    inBuf[947] = 256'hfd058d073f09ec0a8b0cf00d020fda0f6710a710c210a2103610a50fd90ed60d;
    inBuf[948] = 256'hd60cd70bdd0a150a6409b9083408ba074507f806c0069106810677066c067706;
    inBuf[949] = 256'h8906a806e8062f077707c607f80708080608dd0794074107d3064d06c3052e05;
    inBuf[950] = 256'h98041f04c60394039803c60313047c04f2046b05e7056806f60699075d084909;
    inBuf[951] = 256'h550a6e0b8c0c8c0d4e0ece0efa0ebd0e280e3a0de70b500a820885068a04b302;
    inBuf[952] = 256'h0a01b9ffc4fe09fe82fd0ffd7efcd2fb09fb1dfa3af975f8d2f76df736f70ff7;
    inBuf[953] = 256'hf7f6c9f66ef6fcf56ef5c7f42ef49bf309f388f205f27cf103f18ff02df0f3ef;
    inBuf[954] = 256'hd1efd4ef0ef06ef009f1e8f1f3f22cf482f5c1f6e6f7e6f8a2f942fad7fa51fb;
    inBuf[955] = 256'hcbfb43fc87fc9dfc80fc10fc6bfba4faacf99ff88cf75bf628f502f4dcf2d2f1;
    inBuf[956] = 256'hf4f02cf086efffee79eef8ed7fedfaec7fec1fecd4ebbdebeeeb56ec05edf4ed;
    inBuf[957] = 256'hf3eef1efd8f078f1d0f1eaf1b7f156f1e3f05df0ecefaeef9defd5ef5df009f1;
    inBuf[958] = 256'hd1f19cf232f397f3d1f3d5f3d0f3e2f302f450f4d3f465f516f6e6f6aaf770f8;
    inBuf[959] = 256'h30f9b3f9f7f9f7f98ef9def80df81ff746f6a4f51ff5bdf47af41ff4a9f326f3;
    inBuf[960] = 256'h7af2bdf116f175f0e9ef8fef49ef1fef2fef5fefbcef63f02cf110f21af317f4;
    inBuf[961] = 256'hfcf4e2f5a6f651f705f8a2f826f9a6f9f4f90efa10fad9f97ef927f9b5f83bf8;
    inBuf[962] = 256'hd6f75af7d6f667f6e1f55cf5f5f486f427f4f4f3bcf393f385f356f313f3caf2;
    inBuf[963] = 256'h48f2abf111f154f09befffee57eec1ed4bedc4ec4aece5eb64ebe4ea70ead9e9;
    inBuf[964] = 256'h47e9d0e851e8f4e7c8e79de78ce79ae799e7b2e7f7e74be8d3e890e94dea11eb;
    inBuf[965] = 256'hcdeb4deca9ece9ecfdec0fed2bed3fed69ed9fedc2edebed0cee06eef7edd1ed;
    inBuf[966] = 256'h79ed19edadec2beccdeb96eb7eebbbeb3fecf3ecfbed36ef7ef0eaf150f386f4;
    inBuf[967] = 256'ha3f57ff605f759f76ef74ef738f728f729f767f7b8f707f860f891f898f89ef8;
    inBuf[968] = 256'h9cf8b0f810f9a8f97dfa96fbbefcecfd2aff5b009501ef025604d6056a07e808;
    inBuf[969] = 256'h570aa30bb20c9e0d620ef30e7b0ff70f5610c01026116e11b811f111fc11fd11;
    inBuf[970] = 256'he4119e1159111311c710ad10c61008119a1165124a13571467155c164c171f18;
    inBuf[971] = 256'hc6186719ed194b1aac1af61a201b521b6e1b591b2f1bc41a021a1519f017a016;
    inBuf[972] = 256'h6a1547143e137a12d8114c11f910c110a610d4102b11a7115b121013b5135a14;
    inBuf[973] = 256'hc614fd141b15f3148d140c143d132612e810570f860da90bb309d50752061e05;
    inBuf[974] = 256'h4e04f403d003cc03df03d803bf03b503ae03c40308045504a404ea04ff04ec04;
    inBuf[975] = 256'hbf046a040804ab034103d9027e021f02c70180013201dc007e00030075ffe7fe;
    inBuf[976] = 256'h63fe03fedffdf7fd47fec4fe50ffd6ff46009200bd00cb00be00a10073002d00;
    inBuf[977] = 256'hd9ff77ff0affa9fe5dfe26fe0dfe06fef9fde2fdb1fd64fd10fdc5fc97fca0fc;
    inBuf[978] = 256'he2fc56fdf7fda7fe51ffebff58009700ad0094006200360016001a005300a900;
    inBuf[979] = 256'h10017901bd01d601cc01a20178016f018f01e70177022303dc038b0410056505;
    inBuf[980] = 256'h840566052205c70460040d04d703b803be03e003090440047c04a304b604a604;
    inBuf[981] = 256'h5404c6030103080201010f0038ff93fe1dfeb3fd4cfdd8fc43fc9efb01fb6ffa;
    inBuf[982] = 256'h06fad2f9c3f9dff921fa6dfaccfa3afb9cfbfffb5ffca2fcd6fcfafcf5fcd8fc;
    inBuf[983] = 256'ha3fc43fccefb4dfbbafa37fad3f989f973f98ff9caf92dfaaafa27fbaffb33fc;
    inBuf[984] = 256'ha2fc0cfd69fdacfdeafd18fe2bfe35fe31fe12fef5fdd8fdb5fda6fda6fda6fd;
    inBuf[985] = 256'hb4fdc3fdbefdb2fd94fd54fd05fda5fc2efcbafb50fbedfaaafa8afa82fa9ffa;
    inBuf[986] = 256'hd6fa10fb50fb84fb96fb91fb70fb30fbecfaa9fa66fa30fafef9bdf975f920f9;
    inBuf[987] = 256'hc0f870f83df828f83ef874f8b3f8faf83ef97bf9c1f917fa76fadffa43fb8dfb;
    inBuf[988] = 256'hb9fbc7fbb5fb95fb70fb41fb0cfbcbfa72fa0afa9cf92ff9d3f892f864f845f8;
    inBuf[989] = 256'h32f81df806f8f8f7ecf7e7f7f1f7fbf704f814f825f83df870f8b6f814f98ef9;
    inBuf[990] = 256'h12fa97fa1dfb8efbe6fb27fc43fc3afc1afcdbfb87fb32fbd0fa66fafcf97bf9;
    inBuf[991] = 256'he2f836f868f786f6a5f5c5f400f470f310f3edf20ef356f3bff33cf4a9f403f5;
    inBuf[992] = 256'h48f569f57ef599f5b4f5e5f531f680f6d5f622f749f74df72ef7e1f682f61ff6;
    inBuf[993] = 256'hb8f563f520f5daf49af454f4f9f39bf33af3d4f282f241f20ff204f21ff261f2;
    inBuf[994] = 256'he1f290f35cf443f51ff6d6f670f7dcf727f875f8c4f822f9a6f936facefa79fb;
    inBuf[995] = 256'h19fcb4fc58fde6fd65fedefe2eff63ff91ffa6ffc4ff0a006500f200b9018c02;
    inBuf[996] = 256'h76036c043d05fe05b8064c07e8079c084a09160aff0ad90bc60cc50daf0eb20f;
    inBuf[997] = 256'hc810c511cc12c71382142615a315d215ed15ea15ab1573154015ff1400154015;
    inBuf[998] = 256'ha1155b1647172a182b19211ae11ab01b791c231df51dcf1e8a1f66203921e021;
    inBuf[999] = 256'h9b223d23a02300242b240224d2237a23f12291223622d221ae21972174218c21;
    inBuf[1000] = 256'ha621ae21e4210722fe210422d7216b210b218d20f81fa51f681f401f6b1f9a1f;
    inBuf[1001] = 256'hb21fd91fbc1f4c1fca1e021e0a1d321c4b1b5e1aa419d418eb171c172b162915;
    inBuf[1002] = 256'h5e149d13fc12b01272123d122912e7117511fe104e10810fce0e060e3c0d960c;
    inBuf[1003] = 256'hd90b150b750ac7092709bc084c08e10791071e079a062c06af0545051305eb04;
    inBuf[1004] = 256'hda04ee04f004f20408050c05120527051905ef04b3044004b8033c03c0026902;
    inBuf[1005] = 256'h4c024402590285029d02a902ac028a0256021502b3014401cf004900cbff65ff;
    inBuf[1006] = 256'h0fffe4feecfe17ff72ffefff7300f7006b01b501dd01e201c301970163012a01;
    inBuf[1007] = 256'hfb00d300af00990089007d007a0076006b005c0041001700e5ffa1ff4efff4fe;
    inBuf[1008] = 256'h90fe2ffee8fdbffdc7fd0bfe7afe0cffafff3e00b000010128013c0154017301;
    inBuf[1009] = 256'haf010c027902f4027403de03350476048d0482045804fa037703d20202021f01;
    inBuf[1010] = 256'h3a004bff6dfea9fdeffc50fccefb55fbf5fab3fa74fa43fa19fad2f977f907f9;
    inBuf[1011] = 256'h6bf8bff713f75df6bef545f5e1f4acf4b1f4d4f428f5a7f520f695f6f7f614f7;
    inBuf[1012] = 256'h00f7c5f650f6cef55bf5e5f491f469f448f43ff44df441f430f421f4f1f3caf3;
    inBuf[1013] = 256'hc4f3c8f3fbf365f4d1f448f5bbf5ecf5ecf5c4f54ff5bcf425f471f3d0f25bf2;
    inBuf[1014] = 256'hf0f1b8f1bbf1c0f1d5f1eff1caf17ef11cf18af00af0c9efb3eff9efa1f065f1;
    inBuf[1015] = 256'h4df23ff3edf364f4a4f479f40ff481f3b4f2eaf148f1b7f06cf077f09cf0ecf0;
    inBuf[1016] = 256'h54f187f192f177f108f179f0ebef44efbbee67ee1beefeed18ee36ee7ceef4ee;
    inBuf[1017] = 256'h68eff5ef9df025f1acf139f29ef200f36df3aff3e2f30af4eef3b5f377f314f3;
    inBuf[1018] = 256'hc8f2b2f2abf2d4f22ef375f3b8f3f5f3f0f3cef39ff340f3e0f29df257f23bf2;
    inBuf[1019] = 256'h60f298f2fff296f31af497f407f52cf521f5f4f485f408f4a3f344f320f352f3;
    inBuf[1020] = 256'haaf339f4eef478f5d3f5f0f596f5e9f40af4f0f2e2f110f169f01df034f076f0;
    inBuf[1021] = 256'hedf085f1fef163f2b5f2caf2caf2c8f2aaf296f299f28af281f27df24df209f2;
    inBuf[1022] = 256'hb1f123f183f0deef1def6aeed2ed36edb7ec53ece8eb94eb56eb14ebefeae7ea;
    inBuf[1023] = 256'he1eaf9ea2ceb63ebc1eb47ece1eca8ed8bee63ef36f0e6f055f19bf1b6f1a9f1;
    inBuf[1024] = 256'ha2f1aaf1c3f10ef27cf2fbf295f327f499f4f1f41af513f502f5f0f4f9f44bf5;
    inBuf[1025] = 256'he3f5c6f6f5f745f99dfaf5fb26fd34fe32ff1300ec00d101ac02890370044705;
    inBuf[1026] = 256'h22060e07f307e808e909d10aa80b5d0ccc0c0f0d280d0e0df00cdd0cc60cd40c;
    inBuf[1027] = 256'h020d320d850ded0d510edb0e850f3c1034115f12a4132515bb1631189719ba1a;
    inBuf[1028] = 256'h701be51b081cdc1bb11b861b591b631b7a1b781b7a1b481bc91a341a72199018;
    inBuf[1029] = 256'he41765171f175817e417aa18c619ec1af31bf61cb41d1d1e661e5e1e0b1eaa1d;
    inBuf[1030] = 256'h121d541cb11b061b601af51988190f19a61807182c1747163015031407131612;
    inBuf[1031] = 256'h4511bd103b10bc0f590fd10e2e0e9b0dec0c3d0cbf0b440be10ab60a850a550a;
    inBuf[1032] = 256'h3a0af50992092b099308e50746079006e1055505c0043604c8034503c3025302;
    inBuf[1033] = 256'hcc014c01e7007f00330018000c00250064009900c200cd008700faff2eff1dfe;
    inBuf[1034] = 256'hfffc02fc37fbccfacffa1efbadfb52fcd0fc16fd11fdb2fc1bfc69fbb6fa32fa;
    inBuf[1035] = 256'hf3f9fdf957faeefaa0fb55fce7fc33fd2ffdc9fc06fcfbfabef972f83ff73cf6;
    inBuf[1036] = 256'h7ff511f5e3f4ecf419f552f599f5e9f53ef6a5f614f778f7c8f7e9f7c7f771f7;
    inBuf[1037] = 256'hf1f662f6fdf5ddf512f6aef68ff784f866f9ecf9dcf924f9a7f76df5b3f2aeef;
    inBuf[1038] = 256'hb9ec4eeac1e863e875e9e5eb7aefdff376f8a7fcf6ffe70147023401e3fecafb;
    inBuf[1039] = 256'h8ef8acf59bf3b8f201f354f46bf6c4f8e5fa76fc17fdabfc51fb2ff9a3f62af4;
    inBuf[1040] = 256'h22f2eef0e1f005f246f46df7fdfa72fe5001150375036a021100c6fc18f98af5;
    inBuf[1041] = 256'h9cf2baf00cf08ff01ff265f4fbf68bf9b5fb37fdf9fdf1fd32fdf3fb6cfad3f8;
    inBuf[1042] = 256'h6cf75ef6baf58cf5c4f537f6cbf65bf7bef7f4f701f8ecf7e0f700f855f8fcf8;
    inBuf[1043] = 256'hf3f917fb58fc95fd9efe67ffe4fffbffbcff34ff5afe4efd2dfcfcfae6f90af9;
    inBuf[1044] = 256'h61f801f8e5f7e3f7f4f70af801f8ecf7dcf7c5f7cbf7f8f730f87df8d3f807f9;
    inBuf[1045] = 256'h21f91ff9e2f881f805f857f796f6d0f5f5f42ef48cf3fdf29ef272f251f24cf2;
    inBuf[1046] = 256'h5bf25bf26af28df2b1f2f8f268f3e3f382f43bf5ecf5a7f664f701f894f814f9;
    inBuf[1047] = 256'h62f998f9b3f9a1f986f96bf949f945f963f991f9e6f955fac0fa38fbaefb0afc;
    inBuf[1048] = 256'h65fcb6fcedfc22fd4cfd5afd64fd64fd52fd4ffd5afd70fdacfdfffd56febafe;
    inBuf[1049] = 256'h10ff42ff5fff59ff35ff11fff0feddfef0fe21ff67ffc7ff27007800bc00e000;
    inBuf[1050] = 256'he400da00be00a00096009e00c400150181010a02ae025303f5038d0403055905;
    inBuf[1051] = 256'h91059c058b0564051d05c8046404e3035603bf0217027e01ff009b0071007e00;
    inBuf[1052] = 256'hb10011018701f0015702a802d502fa0214031c0332034a035a037f03ae03e003;
    inBuf[1053] = 256'h3704a7042405c6056f0603079207fc07300852085a08490856087a08af081e09;
    inBuf[1054] = 256'hac09430a010bc30b740c3a0df70d9d0e550f011093103811d1115112e5126a13;
    inBuf[1055] = 256'hcf133c148c14b014da14ee14e514fa140d1512153a1557155515671565154815;
    inBuf[1056] = 256'h50155f157415cd154316c9168f175d181719e719911afe1a641b951b8c1b911b;
    inBuf[1057] = 256'h7d1b551b611b761b911bf31b631cd41c771d061e691ecf1ef51ed11ea91e521e;
    inBuf[1058] = 256'hdd1da11d7a1d761ddc1d6c1e161f0320d7207a21122252223a220d229821ef20;
    inBuf[1059] = 256'h5f20b31ff71e6f1edb1d431de61c821c211cf71bbb1b6d1b3c1bdc1a571ae619;
    inBuf[1060] = 256'h4b199e181e188e170117ab164816eb15c2158c155c155e1548152a152515ec14;
    inBuf[1061] = 256'h91143c14ab1301136d12b9110c1191101010a80f760f340ff40ec50e600ede0d;
    inBuf[1062] = 256'h570d9b0cd70b300b7f0af0099d095209320948095c098809c709db09d309a609;
    inBuf[1063] = 256'h200964088107600639051d04f302e601f600070040ffa3fe1afec9fda1fd7efd;
    inBuf[1064] = 256'h6efd53fd0bfdaefc31fc8cfbe8fa44fa99f90df990f819f8c3f777f72ff700f7;
    inBuf[1065] = 256'hd3f6a7f697f691f698f6c4f6f6f629f765f784f78bf78df776f75cf755f744f7;
    inBuf[1066] = 256'h32f71ef7e0f682f610f67af5e4f46cf4fef3b4f391f367f342f31df3d5f287f2;
    inBuf[1067] = 256'h3df2dff18bf143f1e2f083f023f0a8ef39efe1ee8eee6fee86eebaee2eefd5ef;
    inBuf[1068] = 256'h8bf067f155f22af3fff3bff449f5bcf50ff624f623f604f6b1f55bf505f5a5f4;
    inBuf[1069] = 256'h73f46df47ff4c6f428f579f5cef50ef620f62ef636f62df641f66ff6a1f6fcf6;
    inBuf[1070] = 256'h72f7e4f76cf8f1f849f985f98ef946f9d4f83cf87bf7caf635f6b2f569f54ef5;
    inBuf[1071] = 256'h3ef54bf55df54bf528f5eaf477f4f9f37df3fbf2a4f284f284f2bef229f396f3;
    inBuf[1072] = 256'h16f49ef406f56cf5d4f524f67ff6eff64ff7bcf732f883f8c0f8e6f8cbf88bf8;
    inBuf[1073] = 256'h37f8b2f728f7b0f629f6b6f561f5f9f497f445f4d8f378f33df308f303f33ef3;
    inBuf[1074] = 256'h80f3d8f339f453f431f4d3f305f3faf1d9f08def57ee5ded79ecdaeb8beb50eb;
    inBuf[1075] = 256'h47eb6eeb7deb8beb92eb4eebe4ea64eaaae9fce884e827e825e88fe824e9fce9;
    inBuf[1076] = 256'h04ebe8ebbfec81edf3ed45ee89ee92ee9beeb5eeb2eec9ee02ef25ef62efb4ef;
    inBuf[1077] = 256'hdeef0ef042f04bf05ff085f08ff0aff0dcf0def0e2f0e2f0b3f092f085f067f0;
    inBuf[1078] = 256'h6df08df093f0a8f0bdf0a5f093f081f04bf023f000f0bcef88ef5cef1aeff6ee;
    inBuf[1079] = 256'he5eec6eec5eed1eecaeedeee03ef24ef71efdaef46f0d9f07af10df2b6f25ff3;
    inBuf[1080] = 256'hf3f396f433f5b8f546f6c7f62ef79cf7fef74cf8a5f8f7f83af98cf9d8f917fa;
    inBuf[1081] = 256'h60fa9afac0fae7fafbfa00fb13fb29fb4bfb93fbeffb61fcf3fc8bfd27feccfe;
    inBuf[1082] = 256'h63ffefff7b00f5006601d8013a029502ef0235037203ab03d503030440048604;
    inBuf[1083] = 256'heb0473050e06c7068e074a080209a909320ab30a2e0ba00b240cb60c4b0df90d;
    inBuf[1084] = 256'hb40e760f57104f1155127613941491156916f616231704179416e21521155a14;
    inBuf[1085] = 256'ha1131d13c51292129512b012cf120013241335134e1360137413af1301146a14;
    inBuf[1086] = 256'hfb148d150b167816a91694165616de154115ae141b1496133a13e8129a126212;
    inBuf[1087] = 256'h1e12cf118e114111ef10b310751042103c1050108a1003118f112112b7121b13;
    inBuf[1088] = 256'h42134113ff1292122212a0111e11b7104f10ed0fa70f580f040fb30e380e940d;
    inBuf[1089] = 256'hd70cec0bef0a100a4709ad0856081308d907a3074207c4064706c10556052305;
    inBuf[1090] = 256'h0a050f052d0530051805eb048c0415049f031e03ad0263022902120224023b02;
    inBuf[1091] = 256'h580277026d024202fb018501fb007300e4ff69ff0effbffe8bfe77fe6afe75fe;
    inBuf[1092] = 256'h98febafee5fe12ff27ff2fff29ff03ffd0fe93fe3bfedcfd74fdf3fc6bfcd8fb;
    inBuf[1093] = 256'h2bfb74faaef9d0f8f3f721f75ff6d3f57ef55af56df59cf5cbf5f9f515f620f6;
    inBuf[1094] = 256'h34f654f683f6cef61bf756f77cf776f744f7fef6a4f648f604f6d2f5b7f5bff5;
    inBuf[1095] = 256'hd9f505f647f685f6bdf6edf6fcf6f0f6d5f6a0f667f638f608f6e3f5cef5b6f5;
    inBuf[1096] = 256'ha6f5a2f59af59af5a2f59af58df579f550f52af513f504f511f538f55ef587f5;
    inBuf[1097] = 256'ha5f5a7f5a2f5a0f5a3f5c6f506f64af692f6c0f6b8f688f635f6cdf580f563f5;
    inBuf[1098] = 256'h80f5ebf595f65ff745f829f9f2f9a5fa35fb96fbd9fbf8fbf2fbe4fbd3fbcafb;
    inBuf[1099] = 256'he4fb1efc6efcd6fc37fd78fd94fd77fd1dfd9afcf2fb31fb74fabef918f995f8;
    inBuf[1100] = 256'h32f8f3f7e3f7f7f729f879f8d1f828f97cf9bef9eef913fa27fa30fa34fa30fa;
    inBuf[1101] = 256'h2ffa3dfa61faaafa25fbccfb9cfc82fd60fe1effa5ffe8ffeaffb6ff5efffafe;
    inBuf[1102] = 256'h9cfe50fe21fe0cfe0ffe29fe4ffe7cfeaefed9fefefe1fff34ff46ff59ff6aff;
    inBuf[1103] = 256'h83ffa8ffd6ff14006400ba0016016c01a701be01a7015701d90038007dffc0fe;
    inBuf[1104] = 256'h12fe74fdf9fca2fc67fc4dfc4bfc50fc59fc59fc3efc10fccffb7dfb30fbf0fa;
    inBuf[1105] = 256'hbffaaafaacfabafad9fa03fb31fb6bfbadfbeefb34fc77fcb0fceafc24fd63fd;
    inBuf[1106] = 256'haffd05fe5bfeacfee8fe03ff02ffe6febcfe98fe84fe88fea7fed8fe12ff47ff;
    inBuf[1107] = 256'h6cff77ff64ff2fffd9fe66fedefd4ffdc2fc46fce5fb9bfb67fb40fb13fbddfa;
    inBuf[1108] = 256'h9cfa4efa00fac0f98df973f976f98af9b8f902fa5cfacffa57fbd9fb51fcb0fc;
    inBuf[1109] = 256'hdbfcdffcc9fc97fc71fc67fc6bfc8bfcbdfcdbfcf4fc09fd10fd33fd86fdfefd;
    inBuf[1110] = 256'hb6fe9fff8b007c015a02fc028003e70325046804b504f6044d05b20508067506;
    inBuf[1111] = 256'hf60674071b08e208a4097e0a530bf80b8b0cfa0c2a0d520d6d0d6b0d820da80d;
    inBuf[1112] = 256'hc20dfe0d480e800ed50e320f7c0fe40f5610b4103011b01114128f1209136c13;
    inBuf[1113] = 256'hf3138d142715fa15e716cd17d118c619821a2e1ba21bc51bcf1ba71b431be51a;
    inBuf[1114] = 256'h791afb19ae197c1956197319a619d419201a581a621a6b1a4e1a021ac0196c19;
    inBuf[1115] = 256'h0419c2188918541858186c188118ba18de18d718c3187118db1732175b166315;
    inBuf[1116] = 256'h8814b413f4127b122812f7110612201234125612571234121412e011a8119811;
    inBuf[1117] = 256'h95119f11d011ff1126125c127e128e12a112941266122b12c9114d11d8105910;
    inBuf[1118] = 256'hde0f750ffb0e690ec00de80cf00bf80a040a300992081408af075707ea066306;
    inBuf[1119] = 256'hca051a056804c8033603bc025c020302b5016c011f01d10082002a00ceff6dff;
    inBuf[1120] = 256'h03ff98fe2cfebefd56fdf2fc94fc45fc04fcd5fbbcfbacfb9ffb8efb6afb35fb;
    inBuf[1121] = 256'hfcfac4faa6fab4fae5fa37fb99fbe0fbfcfbddfb75fbdafa28fa6af9c7f84cf8;
    inBuf[1122] = 256'hedf7aef780f743f7f9f699f615f680f5e6f43ff4a9f32cf3bcf270f24bf23af2;
    inBuf[1123] = 256'h50f289f2cff22df39af3f7f34df493f4b2f4c1f4c6f4b5f4acf4aff4a5f49cf4;
    inBuf[1124] = 256'h88f449f4f5f393f319f3b3f272f24af253f282f2aef2dcf2fdf2eef2caf29af2;
    inBuf[1125] = 256'h52f21af202f2f9f11df272f2d7f25ef3fdf38af40ef57ff5b4f5c1f5adf564f5;
    inBuf[1126] = 256'h0cf5bbf462f423f407f4ebf3dff3e0f3c2f39bf370f328f3e4f2b6f285f26bf2;
    inBuf[1127] = 256'h71f26ff278f290f292f29bf2bcf2dcf21cf38ef30ff4b0f472f51ef6baf642f7;
    inBuf[1128] = 256'h84f794f785f739f7d9f688f62bf6e8f5d4f5c5f5cff5f9f50cf616f61df6ebf5;
    inBuf[1129] = 256'h96f52ef590f4e1f344f39bf210f2b8f166f12bf10ff1dcf0a9f08bf05df045f0;
    inBuf[1130] = 256'h59f069f089f0baf0c0f0aef095f04af0f9efc0ef79ef45ef34ef13effaeef9ee;
    inBuf[1131] = 256'he2eed6eee6eee2eee3eeeeeeceee9eee74ee30ee03ee12ee40eeb4ee76ef4af0;
    inBuf[1132] = 256'h33f122f2cef244f389f376f33ef300f3acf270f25df248f243f249f226f2f2f1;
    inBuf[1133] = 256'hb7f157f1f9f0acf04df0f5efa4ef30efb8ee47eec9ed6ded47ed41ed7aededed;
    inBuf[1134] = 256'h6eee0aefb3ef3ff0c0f031f173f19ff1b6f1a2f185f169f145f140f165f1a6f1;
    inBuf[1135] = 256'h1bf2b9f25ff312f4b9f434f58ff5c3f5c9f5c6f5c3f5c9f5f6f547f6b0f637f7;
    inBuf[1136] = 256'hc7f74df8d0f844f9a5f905fa5efaaefa04fb56fba5fb04fc6efcebfc88fd33fe;
    inBuf[1137] = 256'he5fe95ff26009000d800f6000301180137017701da014602b502140344034c03;
    inBuf[1138] = 256'h3103f302b90299029602cd023b03c3036a041705a9052e069906df061f075907;
    inBuf[1139] = 256'h8407bf07030842089b0804097209050ab10a620b330c060dc00d760e0c0f6e0f;
    inBuf[1140] = 256'hc10ff70f0c102f1055107610ba1008115011b71123128612091391130d149d14;
    inBuf[1141] = 256'h1b156f15b815d415b81596155b150815d314a6147a147d149114ab14f8145215;
    inBuf[1142] = 256'hac1528169a16ec1640176d17681762173a17f016b51667160016b1155515ed14;
    inBuf[1143] = 256'ha914681425140b14ed13be13a413751330130813e012c112df1211135213be13;
    inBuf[1144] = 256'h19144f147c146b142014d0136413f512be129e129812c312e012db12c7127212;
    inBuf[1145] = 256'he5115311a110e80f560fc20e330ec00d3a0da50c210c8a0bf10a780afd098d09;
    inBuf[1146] = 256'h49090c09e808fc0826097409fa09870a1c0bbe0b370c890cc20cbd0c920c5f0c;
    inBuf[1147] = 256'h100cc50b970b670b440b310b000bb90a5f0ad60937099b08f3076307fd06aa06;
    inBuf[1148] = 256'h7d06770673067b06860670064506020693051805a1043004ed03e20300045104;
    inBuf[1149] = 256'hbb0410054c054f0502057d04c103d602e601f40003002fff6cfeb4fd1cfd98fc;
    inBuf[1150] = 256'h25fcd9fba2fb7afb6efb61fb48fb31fb03fbc2fa88fa4bfa16fa02faf9f9f9f9;
    inBuf[1151] = 256'h08fa02fae1f9b4f964f906f9b9f874f84bf851f863f883f8aff8bef8b8f8aaf8;
    inBuf[1152] = 256'h7ef84ef830f810f8fef702f8faf7f0f7e9f7c7f79ef77df748f715f7ecf6abf6;
    inBuf[1153] = 256'h60f611f69ef520f5a8f422f4b1f368f32ef31af331f34cf377f3aff3cdf3e0f3;
    inBuf[1154] = 256'heff3dbf3c3f3b6f3a0f3a5f3d1f30bf464f4d9f43df594f5d8f5e0f5c3f58ef5;
    inBuf[1155] = 256'h33f5d8f493f455f43af44bf469f4a5f401f55af5c0f534f691f6e6f635f75bf7;
    inBuf[1156] = 256'h6ef778f765f753f757f75ef783f7cff71ef879f8dcf81bf943f95df950f93af9;
    inBuf[1157] = 256'h36f92bf931f94ef956f94af928f9cbf845f8b2f704f765f6f5f5a2f580f597f5;
    inBuf[1158] = 256'hbcf5f1f538f666f688f6adf6b7f6bdf6d3f6ddf6f0f620f749f780f7d0f713f8;
    inBuf[1159] = 256'h56f8a3f8cdf8e5f8f5f8dbf8b2f894f86af856f86ff893f8d3f82ef971f9a0f9;
    inBuf[1160] = 256'hbcf99bf959f909f997f828f8d1f775f72ef701f7c4f68cf65bf609f6b1f55bf5;
    inBuf[1161] = 256'hecf487f43df4f6f3d8f3e5f3f9f325f459f467f462f445f4faf3aff373f33ff3;
    inBuf[1162] = 256'h3ff374f3c0f335f4b7f41cf570f59af583f54ff5fff494f445f416f407f43df4;
    inBuf[1163] = 256'ha1f41bf5b5f547f6baf61ff75df772f784f783f776f780f78bf799f7c6f7f4f7;
    inBuf[1164] = 256'h23f86bf8a6f8d7f811f92df935f942f934f924f92ff938f958f9a5f9f8f962fa;
    inBuf[1165] = 256'hebfa63fbdcfb5cfcb5fc06fd5bfd8cfdc1fd05fe30fe6afebdfefdfe5affdbff;
    inBuf[1166] = 256'h59000301db01b102aa03b904a00582064e07d1073f089708b908ef083b097f09;
    inBuf[1167] = 256'hfc09a30a440b130cf20cae0d810e550f0410d210ac1169124b133114ed14bf15;
    inBuf[1168] = 256'h82160d17a7172e188018e6183b195c198f19ad1998199a199019631966197319;
    inBuf[1169] = 256'h7819c119201a791a0b1b9c1b0a1c941c021d401d9b1de61d181e801eed1e4c1f;
    inBuf[1170] = 256'hde1f5f20b72020215d2162217621662135212a211321ec20f720f920ed201221;
    inBuf[1171] = 256'h2a213221632179216f21782154210321c1205920d71f791f0a1f911e3f1ed81d;
    inBuf[1172] = 256'h5d1dfb1c761cd61b491b981acd1915193b184f177d169615ad14f0132e137a12;
    inBuf[1173] = 256'hf91177110211b6105d10ff0fb40f470fc60e4f0ebb0d280dbb0c560c130c0c0c;
    inBuf[1174] = 256'h150c360c760c9d0caf0cb20c780c110c900bd90a090a3e0964089c07f8065b06;
    inBuf[1175] = 256'hd6056605e6045f04d20325037402ca011c0185000f00a5ff59ff28fffafedbfe;
    inBuf[1176] = 256'hc5fea0fe7afe48fef6fd93fd1afd7ffcddfb32fb7bfad4f935f99af814f895f7;
    inBuf[1177] = 256'h16f7a7f63bf6d0f57bf530f5f3f4d5f4c5f4c2f4d7f4eef406f52df551f579f5;
    inBuf[1178] = 256'hb7f5f9f542f6a0f6f1f634f76df779f75cf722f7b6f62bf69cf5fdf469f4f9f3;
    inBuf[1179] = 256'h99f356f338f314f3ebf2bbf25af2d9f14af19ef0f9ef7cef14efdceeddeee9ee;
    inBuf[1180] = 256'h06ef30ef33ef1feffeeeb0ee56ee06eea6ed58ed2cedfdece4ece9ece0ece1ec;
    inBuf[1181] = 256'hf4ecebece7eceeecd9eccaecccecb7ecb2ecc9ecd6ecfdec47ed85edd4ed36ee;
    inBuf[1182] = 256'h76eeb7eefeee25ef59efa8efe8ef41f0aff0f9f036f161f144f10bf1c8f05ff0;
    inBuf[1183] = 256'h0cf0e4efc3efceef02f01df039f04cf01ff0dfef9aef2fefdceeb1ee8cee9bee;
    inBuf[1184] = 256'he1ee27ef8eef0df069f0c6f022f14ef178f1a9f1b8f1d8f10ef22df261f2aaf2;
    inBuf[1185] = 256'hd9f218f367f39cf3dff332f467f4a3f4e6f401f51df53cf534f532f53af524f5;
    inBuf[1186] = 256'h1cf527f51ef52ff560f589f5d4f53cf691f6eff64cf773f787f785f74bf708f7;
    inBuf[1187] = 256'hc9f676f641f631f625f63df673f694f6b7f6cff6aff678f62ff6bbf54df5f5f4;
    inBuf[1188] = 256'h9ff473f473f475f48ff4b3f4b0f49cf472f414f4aaf341f3c8f26ef23ef21bf2;
    inBuf[1189] = 256'h21f248f261f27ef293f27ff262f246f21bf209f219f231f267f2b1f2e6f215f3;
    inBuf[1190] = 256'h36f32af30ef3e9f2a8f26ff244f211f2f2f1e2f1c7f1b3f1a0f175f147f116f1;
    inBuf[1191] = 256'hcff08df052f00ff0dfefbfef9def91ef93ef8fef98efa3ef9cef99ef92ef80ef;
    inBuf[1192] = 256'h81ef98efc2ef19f095f021f1c3f15ef2d7f236f36ef37df384f389f39af3d7f3;
    inBuf[1193] = 256'h39f4b9f461f512f6bbf65ff7e4f749f8a1f8e1f819f962f9b0f90efa87fa04fb;
    inBuf[1194] = 256'h86fb16fc9afc21fdb9fd50fefafebeff840055013202fb02c10389043c05f405;
    inBuf[1195] = 256'hb90671073408fe08af095f0a0b0b980b2a0cc00c400dcb0d5a0ec80e340f920f;
    inBuf[1196] = 256'hc40ff80f2b104e1099100a11881140121b13ed13d814bc1573162c17d7175f18;
    inBuf[1197] = 256'h0519ba19681a461b341c0c1dfb1dd91e851f3720ce203721b32121226c22d222;
    inBuf[1198] = 256'h2a235c23a823e523022445248424b1240b256325a32508265c268c26d6260527;
    inBuf[1199] = 256'h0c272c272f270b270127d92688265026f62574250c258724e1236123ca221c22;
    inBuf[1200] = 256'h9621f9204320b31f0a1f4c1ebb1d171d671ce41b4a1b9e1a181a7919cf185a18;
    inBuf[1201] = 256'he017721748171c17f016ed16c41678163616bd151f159914f1134513ca124312;
    inBuf[1202] = 256'hc41174110b1195103510a40ff70e570e8c0db50c000c360b750ae1093e09a408;
    inBuf[1203] = 256'h3008a7072107ba063706b3054405b3041a048f03e1022f029201dd003400aeff;
    inBuf[1204] = 256'h23ffb3fe70fe2dfe03fefbfde2fdcefdc6fda0fd79fd5efd2dfd09fdfafce1fc;
    inBuf[1205] = 256'hdbfceafceffc03fd26fd38fd4efd63fd56fd3cfd13fdc1fc65fc02fc8cfb23fb;
    inBuf[1206] = 256'hcafa74fa3dfa1ffa0bfa12fa2bfa41fa63fa83fa92faa2faa9fa9ffa9cfa97fa;
    inBuf[1207] = 256'h8cfa8ffa95fa98faa8fab6fabcfac7fac6fab6faa1fa79fa3ffa04fabef974f9;
    inBuf[1208] = 256'h3bf909f9e5f8dff8e8f804f939f974f9b2f9f5f926fa45fa59fa52fa3dfa2afa;
    inBuf[1209] = 256'h10fa01fa09fa17fa34fa64fa8dfab5fae0faf5fa01fb07fbf3fad4fab1fa7bfa;
    inBuf[1210] = 256'h48fa23fa01faf5f905fa17fa30fa49fa3dfa14fad0f95ff9dff866f8ecf792f7;
    inBuf[1211] = 256'h64f746f747f75ef765f768f765f743f71df7fff6d5f6bdf6bdf6b9f6c5f6e1f6;
    inBuf[1212] = 256'hfaf626f759f779f79ef7cff7f0f71bf84ef86bf884f89bf892f884f878f85ef8;
    inBuf[1213] = 256'h4ef855f85af86df892f8a9f8bff8d8f8daf8d3f8cdf8aef886f865f832f802f8;
    inBuf[1214] = 256'he6f7c8f7b8f7c6f7d0f7def7f9f7fbf7eaf7daf7aff777f74ef720f7fdf6faf6;
    inBuf[1215] = 256'hf7f6f9f613f719f713f71bf70ff7fcf609f718f736f77ef7c3f706f85af890f8;
    inBuf[1216] = 256'habf8cdf8d1f8cbf8e8f806f935f997f9f8f95ffae5fa4efb9dfbeffb10fc10fc;
    inBuf[1217] = 256'h12fcecfbb9fba0fb71fb49fb4cfb3cfb2bfb35fb1cfbf5fad9fa92fa3efafaf9;
    inBuf[1218] = 256'h96f936f9f9f8abf86ef858f82df809f8f5f7bbf782f75ef721f7fbf6fbf6edf6;
    inBuf[1219] = 256'hf5f616f716f712f707f7c7f680f638f6d7f597f57bf562f582f5cdf50bf66ef6;
    inBuf[1220] = 256'hc9f6eff61af71cf7e5f6b2f671f616f6dff5c6f5b2f5caf5f9f52cf67ef6cef6;
    inBuf[1221] = 256'h11f75cf78bf798f79ff782f74ef72ff714f711f74ef7b3f748f814f9e9f9c3fa;
    inBuf[1222] = 256'h97fb37fcb7fc1dfd4efd76fdadfde5fd46fed7fe79ff42002001ed01c5029403;
    inBuf[1223] = 256'h3a04e1047905ed056d06e4064607c5074808c1086609170ac60aa40b850c570d;
    inBuf[1224] = 256'h3e0e090fac0f5710da103711a71100124b12c3123713ad135814fb149b156516;
    inBuf[1225] = 256'h1517b2176418ea184e19be19fd19251a6b1a931ac11a251b7c1be01b761cf11c;
    inBuf[1226] = 256'h611de11d241e491e731e651e4d1e561e461e471e7d1e9d1eca1e161f361f4c1f;
    inBuf[1227] = 256'h6c1f531f2d1f141fce1e891e601e151ed51daf1d631d171dd91c6a1cf71b911b;
    inBuf[1228] = 256'h071b881a201a9a192019bc183218a91728177416ba15071526144f138f12b311;
    inBuf[1229] = 256'hf3105510a00f020f7b0ecd0d260d860cb60bed0a330a56099408f10734079506;
    inBuf[1230] = 256'h0e066405ce0442048d03e8024e028d01e200460087ffe4fe58feb4fd31fdc0fc;
    inBuf[1231] = 256'h35fcc4fb5bfbc9fa45fac0f913f97df8f2f74ff7cff663f6ecf596f549f5e3f4;
    inBuf[1232] = 256'h91f438f4c0f360f309f3abf279f261f24ff260f26df263f25ff23ff200f2c7f1;
    inBuf[1233] = 256'h82f137f10ef1eef0d3f0d2f0cdf0c8f0d0f0c7f0b4f0adf096f07bf06ef053f0;
    inBuf[1234] = 256'h39f02ff01ef018f02af036f04ff081f0a4f0c7f0eff0f7f0f6f0fbf0ecf0ecf0;
    inBuf[1235] = 256'h08f121f155f1a6f1e7f12cf27af2a3f2bef2daf2d9f2def2f8f205f32cf35ff3;
    inBuf[1236] = 256'h7ff3acf3d0f3c8f3b2f394f34bf307f3dbf29ff27ef288f288f299f2bbf2b7f2;
    inBuf[1237] = 256'haaf2a2f270f23cf21af2e1f1b9f1aff194f185f18df177f162f159f130f108f1;
    inBuf[1238] = 256'hf1f0b9f082f05af011f0c6ef88ef30efdfeea6ee5cee21ee03eed4edb1eda2ed;
    inBuf[1239] = 256'h74ed42ed19edd1ec8eec60ec24ecfeebfdebf5eb01ec28ec3bec53ec71ec74ec;
    inBuf[1240] = 256'h73ec79ec6cec62ec66ec57ec58ec6cec6fec8becc8ecf8ec3fed99edd4ed0fee;
    inBuf[1241] = 256'h47ee52ee56ee5dee4aee4dee6cee83eebdee18ef67efc9ef30f070f0aff0e7f0;
    inBuf[1242] = 256'hfaf018f147f167f1a3f1f6f13df296f2f3f234f380f3d5f316f46cf4ccf415f5;
    inBuf[1243] = 256'h61f5a6f5c0f5ccf5c8f5a8f597f598f59ef5caf516f65ff6b5f60af73ff769f7;
    inBuf[1244] = 256'h82f77bf777f77df77df793f7bff7eef72cf874f8aef8e9f824f94af96ff99bf9;
    inBuf[1245] = 256'hb9f9dff90ffa36fa61fa96fac3faf8fa34fb63fb93fbc7fbebfb0cfc28fc2cfc;
    inBuf[1246] = 256'h28fc20fc07fceafbcefbabfb91fb83fb73fb73fb83fb94fbaefbc8fbd2fbd8fb;
    inBuf[1247] = 256'hd6fbc3fbadfb97fb82fb80fb8dfba5fbcdfbf5fb0ffc1ffc18fcf7fbc8fb89fb;
    inBuf[1248] = 256'h46fb0cfbd8fab1fa9efa8ffa84fa80fa77fa72fa7afa83fa9afac4faf3fa31fb;
    inBuf[1249] = 256'h80fbcffb2cfc96fcfefc77fdfcfd79fefdfe82fff1ff5f00ce002c0194010802;
    inBuf[1250] = 256'h7b020803a3033304cd046205d00537069506d6062a079007f70789083709da09;
    inBuf[1251] = 256'h920a430bc90b540cd20c2a0d9c0d1b0e880e1d0fc10f4c10f3109f113012e612;
    inBuf[1252] = 256'ha813561435152016e816ca179b183219db19751ae61a841b311cd21cb21d9c1e;
    inBuf[1253] = 256'h621f43200621862117228d22d5224e23cc233224d3246f25dc256426ca26f926;
    inBuf[1254] = 256'h4d279427c2273328a72802298f29fc29272a5e2a632a2e2a232a0f2aef291e2a;
    inBuf[1255] = 256'h532a782acc2af72ae62ae22aa52a302adf297329f528b6286b280b28db278d27;
    inBuf[1256] = 256'h1527b72637269d253025a324ff238323e02220228521c620fb1f5f1fa91ef11d;
    inBuf[1257] = 256'h6b1dca1c201c981be41a1c1a6f199618b317f5161b1643158f14b813d9120b12;
    inBuf[1258] = 256'h0e110610120ff90dea0c020c050b160a4509550863077c067005670473036a02;
    inBuf[1259] = 256'h7601a100c1fff6fe3ffe71fdadfcf5fb2afb73fad4f932f9aaf836f8b9f747f7;
    inBuf[1260] = 256'hcff63af6a6f50cf567f4dbf367f304f3cbf2a9f290f287f271f245f20ff2bef1;
    inBuf[1261] = 256'h5cf103f1aff071f05ef061f082f0c5f006f145f17ef196f19af193f16ff14cf1;
    inBuf[1262] = 256'h32f10ef1fcf001f100f110f130f145f167f191f1a8f1caf1f2f105f221f240f2;
    inBuf[1263] = 256'h47f259f272f27af294f2bff2e4f225f37df3ccf329f488f4cdf414f556f57ef5;
    inBuf[1264] = 256'hb7f5fff53bf68ef6f4f64ef7b8f72af888f8eff857f9a7f9f9f944fa6bfa89fa;
    inBuf[1265] = 256'h9afa86fa6efa58fa32fa20fa28fa2ffa4cfa7afa95faa9faaffa89fa50fa0cfa;
    inBuf[1266] = 256'hacf955f913f9d1f8acf8a7f89af892f88bf866f837f805f8b9f76bf72af7dcf6;
    inBuf[1267] = 256'h98f664f61df6d7f59ef556f51df5fff4e1f4d9f4f0f4fff40df518f5fbf4c6f4;
    inBuf[1268] = 256'h87f428f4d0f398f36df36cf39df3d2f311f451f464f457f431f4d9f374f318f3;
    inBuf[1269] = 256'hb2f264f237f206f2e7f1d8f1b4f196f183f15bf13ef132f116f102f1f2f0c1f0;
    inBuf[1270] = 256'h8bf054f003f0c7efaaef90ef9fefd4ef03f03cf072f07af073f063f035f018f0;
    inBuf[1271] = 256'h18f018f03df07ef0aef0e6f01df12df140f15bf160f17cf1b1f1d9f111f24ef2;
    inBuf[1272] = 256'h67f27cf28ff283f288f2a7f2c3f204f369f3c1f323f483f4b5f4daf4f7f4f3f4;
    inBuf[1273] = 256'hf9f416f529f552f58cf5aef5d1f5f2f5f2f5f5f504f605f618f640f658f671f6;
    inBuf[1274] = 256'h8bf68bf68af694f697f6b5f6f9f647f7b1f72ff896f8eff833f946f93ef92af9;
    inBuf[1275] = 256'h00f9e0f8d9f8def8fdf836f96ff9acf9e7f908fa1ffa2ffa2bfa25fa25fa23fa;
    inBuf[1276] = 256'h2bfa42fa5ffa8cfac4fafdfa3ffb82fbbbfbf1fb1efc39fc48fc45fc31fc13fc;
    inBuf[1277] = 256'he6fbb0fb7dfb49fb24fb18fb1afb34fb68fba0fbe1fb25fc52fc72fc88fc8bfc;
    inBuf[1278] = 256'h98fcbbfcecfc4efde4fd92fe66ff4d001e01e50194020f037b03dd0329049004;
    inBuf[1279] = 256'h13059a054b061807dd07b9089a095b0a230be50b820c270dc90d4c0ee40e850f;
    inBuf[1280] = 256'h1410c61086113012f512ba135a140715a7151c16a0161f17811703188818f118;
    inBuf[1281] = 256'h7819f719501abc1a1a1b551bb11b101c611ce01c621dc81d451ea31eca1ef51e;
    inBuf[1282] = 256'hff1ee91e001f231f521fcb1f5920e32092211f227822cf22f322ea22fc22fe22;
    inBuf[1283] = 256'hf82225234b2363239423992372235123fc2283221d229521fa207a20dc1f2f1f;
    inBuf[1284] = 256'h9d1eef1d391da61cfa1b491bb21af51923195c1866176216771578148913cc12;
    inBuf[1285] = 256'h0c126211db1038108c0fe20e040e160d2f0c2b0b360a68099808e9075c07c306;
    inBuf[1286] = 256'h3706b3050a055d04aa03d202f7011c0126003aff59fe6efd9dfcdffb20fb7bfa;
    inBuf[1287] = 256'hdef931f98bf8d8f708f738f65ff578f4abf3ebf238f2abf12df1b9f05ff001f0;
    inBuf[1288] = 256'ha0ef4feff2ee93ee47eef2ed9bed53edfbeca1ec53ecf6eb9deb5aeb11ebd9ea;
    inBuf[1289] = 256'hc0eaa5ea9feab6eac4eaddea02eb0aeb0deb0cebe9eac6eaadea8aea86eaabea;
    inBuf[1290] = 256'hd8ea2deba1eb08ec77ece3ec22ed59ed87ed98edbdedfded40eeb1ee49efdeef;
    inBuf[1291] = 256'h8ff04bf1e7f185f21cf38df302f476f4c8f420f574f5a4f5d8f50ef62bf65ef6;
    inBuf[1292] = 256'ha7f6edf654f7d1f73bf8abf80ff942f964f977f965f960f971f981f9b4f904fa;
    inBuf[1293] = 256'h49fa96fadefafdfa11fb1efb0cfb03fb08fb01fb07fb1dfb1dfb22fb2cfb1ffb;
    inBuf[1294] = 256'h14fb12fbfbfae7fad9faaffa83fa5cfa1cfae0f9b5f97ef951f938f90bf9d8f8;
    inBuf[1295] = 256'ha4f849f8ddf770f7eaf66df610f6b8f57cf563f541f51df5fbf4b2f456f4f9f3;
    inBuf[1296] = 256'h82f30cf3b3f259f210f2e0f19ff15bf120f1cef07ef046f00cf0e9efe7efe0ef;
    inBuf[1297] = 256'he0efe5efcaefa3ef7eef45ef1eef1fef30ef6aefd0ef36f0a6f014f15cf18ff1;
    inBuf[1298] = 256'hb0f1adf1a6f1a6f19df1a9f1cff1f6f135f286f2ccf218f360f38bf3aff3c7f3;
    inBuf[1299] = 256'hc4f3caf3daf3e9f319f463f4b0f414f579f5c6f50af638f644f64ff65bf668f6;
    inBuf[1300] = 256'h9bf6eef653f7ddf770f8f4f871f9d4f911fa44fa69fa85fab8fafbfa46fbaafb;
    inBuf[1301] = 256'h10fc68fcbffc02fd2cfd52fd6dfd7ffd9bfdb7fdcdfdecfd03fe10fe23fe33fe;
    inBuf[1302] = 256'h44fe67fe95fec8fe09ff46ff77ff9fffb4ffb5ffb1ffa5ff97ff96ff99ffa1ff;
    inBuf[1303] = 256'hb3ffc4ffd3ffe5fff6ff080021003a0053006a00760077006e0058003f002c00;
    inBuf[1304] = 256'h200025003a0056007800930099008c006b003300faffc7ff9eff90ff9bffb1ff;
    inBuf[1305] = 256'hd9ff04002300440062007a00a400de001f017701da0130028b02de021f036b03;
    inBuf[1306] = 256'hc3031d049b042d05b8055206dd063f079607d807fb0732087c08cc084b09e309;
    inBuf[1307] = 256'h720a160baf0b1e0c920cfa0c430da70d150e6f0ee90e630fbb0f28109110e010;
    inBuf[1308] = 256'h5a11e81170122e13f7139d145315eb153f169616d916f9164e17c0173918fe18;
    inBuf[1309] = 256'hdd19a81a961b6a1cfc1c931d051e3f1e971eea1e251f991f142079201121a221;
    inBuf[1310] = 256'h1222ac22332391230b2464248324af24b0247a2463243a240024072415241c24;
    inBuf[1311] = 256'h5b2483247e2485245024dc237123dd223022b4213321b52076202c20d81faa1f;
    inBuf[1312] = 256'h5d1ff81eac1e3a1eaf1d3d1da21cf21b5a1ba11ae3195019b1182118c4175717;
    inBuf[1313] = 256'he6168216e71525155514461323121411f40ff30e280e600db10c1a0c590b830a;
    inBuf[1314] = 256'h990972083a070606c0049b039f02ac01e0002e006dffb8fe03fe32fd6afca6fb;
    inBuf[1315] = 256'hd1fa12fa59f997f8ecf746f799f607f67df5f1f481f413f49cf335f3c2f23df2;
    inBuf[1316] = 256'hc3f139f1a5f028f0a5ef27efc7ee65ee09eec7ed7eed3aed0cedd1ec96ec67ec;
    inBuf[1317] = 256'h1deccaeb7ceb12ebabea5dea0eeadfe9dfe9e8e910ea52ea81eaafeadbeadfea;
    inBuf[1318] = 256'hdceae0eaceead5eaffea2eeb86eb03ec7bec06ed98ed06ee70eed1ee0bef47ef;
    inBuf[1319] = 256'h87efafefe9ef34f072f0c9f035f196f10bf28bf2f2f25ef3c4f303f43ff476f4;
    inBuf[1320] = 256'h8ff4b3f4e4f408f543f58ef5ccf519f66bf6a5f6e5f625f74af777f7aaf7c9f7;
    inBuf[1321] = 256'hf5f72cf856f88ef8d5f812f95ef9b9f906fa5dfab9fafafa38fb70fb8afb9efb;
    inBuf[1322] = 256'hb3fbb2fbb6fbc3fbc2fbc7fbd5fbd1fbd1fbd7fbcbfbc2fbc0fbacfb99fb88fb;
    inBuf[1323] = 256'h60fb2ffbfafaacfa5bfa14fac9f993f97ef974f97ef997f99af989f961f90af9;
    inBuf[1324] = 256'h99f826f8adf74ef71ff70df724f75ef793f7c1f7e2f7d9f7b6f788f745f70af7;
    inBuf[1325] = 256'he5f6c8f6c4f6d7f6e8f6fef617f71df720f725f71af710f70af7f5f6ddf6c5f6;
    inBuf[1326] = 256'h9bf673f651f62cf615f60ef607f60af614f611f60df609f6f9f5eff5edf5eaf5;
    inBuf[1327] = 256'hf4f508f616f62df649f65bf677f69cf6c1f6f4f631f765f798f7c1f7d2f7d9f7;
    inBuf[1328] = 256'hdaf7d3f7dff701f832f87bf8cdf80df93cf94bf92ff9fcf8bff882f865f870f8;
    inBuf[1329] = 256'h9df8f1f857f9b2f9fbf923fa1cfafcf9cef9a1f991f9a9f9e7f94ffacffa4efb;
    inBuf[1330] = 256'hc6fb22fc55fc6efc6efc5efc56fc61fc82fcc2fc19fd7dfdecfd55feacfef8fe;
    inBuf[1331] = 256'h31ff56ff77ff94ffb1ffdcff120051009c00e7002c0169019201a601af01aa01;
    inBuf[1332] = 256'ha001a001a901c001e5010d023502570267026e02730275028c02c1020d037603;
    inBuf[1333] = 256'hf3036b04dd0438056f059605b605d3050e066e06e5067d072408b3082f098709;
    inBuf[1334] = 256'haa09b909bd09ba09d9091c0a700ae50a610bbe0b0b0c340c2a0c170c010ce60b;
    inBuf[1335] = 256'hf30b220c5b0cb60c140d530d8e0dae0da40da10d9f0d970dba0df90d400eb00e;
    inBuf[1336] = 256'h2c0f960f12108010cd1027117811b51117128612f61295134114e01492152b16;
    inBuf[1337] = 256'h9116ed161f172117301739173e177a17ca1718188618db18f9180219cd185b18;
    inBuf[1338] = 256'hf0177e171717fa16051728177a17b517bb17a5174717ac1616167915f614c314;
    inBuf[1339] = 256'hb914d01414153f153a151915af1412147513ce124112f911d211cd11f111fa11;
    inBuf[1340] = 256'hde11a61126117810c10ff30e350ea80d2d0dd20c9b0c540c000c9c0b010b470a;
    inBuf[1341] = 256'h7c098e08a607d70611066f05f20478040a049a0305035f02a801d4000b0056ff;
    inBuf[1342] = 256'haefe33fed8fd83fd41fdf6fc89fc0dfc76fbc5fa21fa8af903f9aef875f847f8;
    inBuf[1343] = 256'h2cf8fcf7a1f72ef78ef6cdf517f567f4d4f37ff349f329f322f300f3b8f256f2;
    inBuf[1344] = 256'hbff108f15cf0b2ef2aefe3eebfeec3eef1ee10ef1eef1befdeee7bee0fee8ded;
    inBuf[1345] = 256'h1dede0ecc2ecdbec30ed8aedeeed4bee6cee61ee38eedced7ded3eed14ed29ed;
    inBuf[1346] = 256'h85edf8ed8dee2def9aefe1efffefd7ef97ef5eef20ef0def31ef67efbdef22f0;
    inBuf[1347] = 256'h5ef080f084f04af003f0c3ef7eef62ef77ef9defe3ef38f06ef09bf0b6f0a8f0;
    inBuf[1348] = 256'h9ff0abf0bcf0fdf06ff1eff18cf234f3baf333f495f4c9f4f7f429f550f591f5;
    inBuf[1349] = 256'hedf547f6b5f62cf788f7e0f72ef856f875f88cf885f87df877f85ef852f855f8;
    inBuf[1350] = 256'h51f85ff87cf88cf8a0f8b2f8a7f896f883f85ef844f83bf832f83ef85df873f8;
    inBuf[1351] = 256'h90f8b1f8bef8cef8e5f8f4f812f942f96ff9a8f9e7f911fa32fa47fa3dfa2bfa;
    inBuf[1352] = 256'h19fafbf9eaf9e9f9e5f9e9f9f2f9e5f9d0f9b6f983f94ff91ef9dbf898f855f8;
    inBuf[1353] = 256'hf8f795f732f7c3f662f61bf6e2f5c7f5c6f5bef5b4f59cf559f5fdf494f41af4;
    inBuf[1354] = 256'hb3f374f359f375f3c4f329f49ff414f567f59ef5baf5aff59af58cf583f595f5;
    inBuf[1355] = 256'hc5f506f663f6cdf62bf786f7d4f702f81ff82df824f81bf816f811f81ef838f8;
    inBuf[1356] = 256'h52f879f8a2f8bef8dcf8f4f801f916f931f94bf973f9a0f9c6f9edf90afa14fa;
    inBuf[1357] = 256'h1cfa1cfa18fa28fa4afa7efacffa31fb99fb05fc5efc9dfccbfcddfcddfce2fc;
    inBuf[1358] = 256'hedfc0efd51fdaafd16fe91fefefe5bffa6ffd2ffecff0500170039007300b300;
    inBuf[1359] = 256'h02015c01a601e8012102410262028a02b102f0024803a2030a047604c7040f05;
    inBuf[1360] = 256'h490568059005c70506066f06fd06980750080c09ab09410aba0a030b430b790b;
    inBuf[1361] = 256'ha00be50b420ca60c320dcb0d500edc0e4e0f890fb40fbc0f970f7e0f660f490f;
    inBuf[1362] = 256'h5f0f910fc90f2c109310dc102a11571151114b113011fe10f61004111b116f11;
    inBuf[1363] = 256'hda114012c6123d138c13e51324143e147414a714ce1423158015d1154616b016;
    inBuf[1364] = 256'hfb165b17a317ca170818391852188b18b618c418e918f118cf18bc188e184018;
    inBuf[1365] = 256'h1218da1796177f176117321727170617c4169c165d160716d915aa157c158915;
    inBuf[1366] = 256'h9e15b415fc153b166616ac16d416dc16f516ef16cf16cb16bc16a616bd16d316;
    inBuf[1367] = 256'he7161f173f173e1740171217b5165a16da154a15dc146d140914d513a0136913;
    inBuf[1368] = 256'h471303139c122d128b11c9100c10390f690ec60d2f0db40c6c0c2a0cf20bcc0b;
    inBuf[1369] = 256'h890b2e0bcf0a460aa90916097808ea0788073707080708071007260748075007;
    inBuf[1370] = 256'h46072d07e9068c062306a1051c05a3042904c403790333030003d50297024e02;
    inBuf[1371] = 256'hea015a01ae00e7ff05ff29fe59fd9bfc09fc9bfb47fb15fbecfab9fa84fa38fa;
    inBuf[1372] = 256'hd1f961f9e4f860f8eef785f727f7e4f6acf680f66cf65ef658f666f670f676f6;
    inBuf[1373] = 256'h80f670f64af61cf6d5f588f546f508f5e3f4e2f4ebf407f536f552f563f56af5;
    inBuf[1374] = 256'h52f52bf503f5c9f496f472f446f423f410f4f0f3dbf3d6f3cbf3cff3e9f3fdf3;
    inBuf[1375] = 256'h1af43df445f443f439f410f4e8f3d0f3bbf3caf306f454f4bff43bf5a3f5fef5;
    inBuf[1376] = 256'h4cf672f685f691f686f681f68bf68ef6a2f6c3f6daf6fcf628f745f767f78cf7;
    inBuf[1377] = 256'h9af7a0f79bf775f745f711f7c9f690f674f665f67cf6b8f6fbf651f7abf7e5f7;
    inBuf[1378] = 256'h0ff829f820f814f811f80cf822f855f88bf8d5f82bf96ff9b0f9f1f91cfa46fa;
    inBuf[1379] = 256'h72fa8efaa9fac3fac3fabefab5fa96fa79fa6cfa5cfa59fa68fa6dfa71fa6dfa;
    inBuf[1380] = 256'h46fa0afabef954f9eaf88df82df8e5f7b7f788f761f73ff709f7d2f69ff65ff6;
    inBuf[1381] = 256'h31f619f601f6fcf509f609f60ef619f615f618f625f629f638f64ff655f65cf6;
    inBuf[1382] = 256'h65f65af651f652f64cf655f66ff680f699f6b1f6aaf694f66ef628f6e1f5a4f5;
    inBuf[1383] = 256'h6af551f55cf573f5a1f5d6f5f2f5fef5f2f5bdf57af531f5ddf4a1f482f473f4;
    inBuf[1384] = 256'h8df4c5f40af568f5cdf524f67df6c9f6f7f61ef73af744f75df784f7b5f70bf8;
    inBuf[1385] = 256'h7af8f4f884f916fa92fa03fb59fb8afba9fbb5fbaefbaffbb7fbc4fbe7fb15fc;
    inBuf[1386] = 256'h44fc7efcb3fcdefc0dfd38fd5bfd85fdadfdccfde8fdf7fdfbfd00fe01fe09fe;
    inBuf[1387] = 256'h29fe5cfea7fe0eff80fff7ff6f00d400260165018c01a801c701e70118026102;
    inBuf[1388] = 256'hb50219038603ec034d04a504ed0432057105a705e0051906460672069806b306;
    inBuf[1389] = 256'hcf06eb06060731076707a207f10747089708ea082d0957097409730954092d09;
    inBuf[1390] = 256'hfb08c808ad08a508b508ee0839098709df091f0a390a3a0a100abf096a091209;
    inBuf[1391] = 256'hc408a508ab08d3082a098a09e0092d0a530a490a270ae5098f0948090709d008;
    inBuf[1392] = 256'hb808aa089e08a308a108950895088f088208860885087f0885087f086a085908;
    inBuf[1393] = 256'h3e081e08130810081b084a088508c1080d094c0973099309990989097a095f09;
    inBuf[1394] = 256'h400934092a09230936094a095b0977098b09900995098709680948091809dd08;
    inBuf[1395] = 256'hab08730836080908db07ac0787075f0735071007e406b6068f0660062e060006;
    inBuf[1396] = 256'hca058c054f050a05c5048a0452042a0417040d0411042004280427041b04f703;
    inBuf[1397] = 256'hc60388033c03f302af027002430222020602f701ea01d201b30183013b01e500;
    inBuf[1398] = 256'h7900f7ff73ffe5fe51feccfd50fddffc87fc3bfcf9fbc6fb8afb42fbf5fa8efa;
    inBuf[1399] = 256'h13fa99f914f992f82af8cef78af76bf758f756f76bf776f778f779f759f724f7;
    inBuf[1400] = 256'he8f68ff62df6daf583f53bf515f5f7f4eef401f50bf513f51ff50bf5e5f4b9f4;
    inBuf[1401] = 256'h71f423f4e4f39df367f34df332f329f335f336f340f355f356f358f361f351f3;
    inBuf[1402] = 256'h3ef32df302f3daf2bdf293f27cf27df279f28cf2b4f2ccf2ecf215f328f33ff3;
    inBuf[1403] = 256'h5af35ff36af37cf377f379f384f37ef387f3a1f3b3f3dcf31df455f49bf4e9f4;
    inBuf[1404] = 256'h1cf549f569f564f559f54cf52cf520f52af535f55af597f5ccf50df655f689f6;
    inBuf[1405] = 256'hbff6f1f604f712f71af701f7e7f6d0f6adf69df6a6f6b4f6e3f62cf771f7c4f7;
    inBuf[1406] = 256'h16f849f86ff882f870f856f83df81af810f823f83df873f8c1f808f956f9a5f9;
    inBuf[1407] = 256'hdbf90bfa36fa45fa4bfa4bfa32fa17fa01fae1f9d4f9e3f9fef936fa89fadefa;
    inBuf[1408] = 256'h38fb8cfbc1fbe0fbeafbcefba6fb7efb50fb36fb39fb4bfb79fbbbfbf8fb38fc;
    inBuf[1409] = 256'h6efc85fc89fc80fc5cfc30fc02fccafb9cfb7afb58fb46fb47fb4afb57fb69fb;
    inBuf[1410] = 256'h6dfb6bfb62fb43fb20fbfffad9fabffab2faa6faa2faa3fa9afa8ffa83fa72fa;
    inBuf[1411] = 256'h6afa72fa87fab2faf0fa35fb7dfbbbfbe2fbf6fbf6fbe7fbdafbd9fbf1fb28fc;
    inBuf[1412] = 256'h7bfce5fc60fdd9fd45fea1fee3fe0eff26ff2cff2aff29ff27ff2fff45ff63ff;
    inBuf[1413] = 256'h90ffcdff0e0052009600ca00f10007010201ec00cc00a1007d00680062007900;
    inBuf[1414] = 256'hac00ee004701ac0108026002ad02e3020e032c03370347035c036f039a03da03;
    inBuf[1415] = 256'h23048b0405057d05fc057006c306070732073a07450751075a078307c2070608;
    inBuf[1416] = 256'h6708d1082d099109ee09340a820aca0afe0a420b830bac0be00b0d0c210c400c;
    inBuf[1417] = 256'h5f0c700c9e0cd90c100d670dc50d120e6e0ebb0ee40e0f0f260f1a0f1c0f1a0f;
    inBuf[1418] = 256'h0b0f210f460f710fcd0f37109c1022119b11ed113f126e1267125d123b120112;
    inBuf[1419] = 256'heb11e311e2111f127312c7124213b4130014501479146f1467144214fc13d513;
    inBuf[1420] = 256'hb11388139513b513dc133a149e14f2145e15a915bc15c21594152c15cc145f14;
    inBuf[1421] = 256'hec13b813a413a913ef133e148114d514ff14f114dc149c143414e01385132813;
    inBuf[1422] = 256'hfd12de12c712e112fa120b133b135913571362134c130f13d71281121612cc11;
    inBuf[1423] = 256'h821143113b1140114b1173118611781168113011d7108b103610e40fbb0f9c0f;
    inBuf[1424] = 256'h830f870f790f540f310fed0e900e400ee50d8d0d540d1d0dec0cce0ca00c640c;
    inBuf[1425] = 256'h2d0cdb0b750b160ba50a2f0ac8095909f208a90866083408230815080c080a08;
    inBuf[1426] = 256'hee07bb0776070d078f0616069a053305f304cd04cc04ec040f0532054b054105;
    inBuf[1427] = 256'h1705d0046604ec036e03ec027d022602df01b401a30199019c019c0187016201;
    inBuf[1428] = 256'h1d01ab001f0078ffbafe06fe5ffdcefc6afc25fcf8fbe5fbd2fbacfb7afb28fb;
    inBuf[1429] = 256'hb2fa2ffa9bf900f97af802f89df75df72ff711f70af702f7f9f6fbf6f0f6ddf6;
    inBuf[1430] = 256'hcdf6aef686f660f62af6eff5bef584f550f531f512f501f506f508f510f524f5;
    inBuf[1431] = 256'h20f50ff5f6f4b7f466f412f4a7f343f3fdf2c2f2acf2c3f2e1f212f354f377f3;
    inBuf[1432] = 256'h86f384f354f315f3d8f288f24bf231f21ef228f252f276f2a7f2e5f209f32ef3;
    inBuf[1433] = 256'h59f369f37af392f38ef38ef396f38bf38ff3aaf3c3f3fcf353f4a3f403f56bf5;
    inBuf[1434] = 256'hadf5ddf5fbf5e8f5cbf5a9f573f553f551f54ff570f5b0f5e5f529f674f69ff6;
    inBuf[1435] = 256'hc3f6daf6cbf6b5f69cf66bf64af643f63bf657f695f6d2f61ff774f7a7f7c8f7;
    inBuf[1436] = 256'hd4f7b1f782f74ef709f7dbf6cdf6c5f6d9f605f725f745f760f75ef756f74cf7;
    inBuf[1437] = 256'h2ff71cf714f7fff6f4f6f1f6dff6d3f6d3f6cdf6d6f6f1f607f728f74af753f7;
    inBuf[1438] = 256'h4ff73df70bf7d4f6a6f678f666f679f69cf6d5f61df752f777f787f76df73ef7;
    inBuf[1439] = 256'h0af7caf69bf68ff695f6b7f6f6f634f770f7a3f7b4f7acf792f75bf71bf7e4f6;
    inBuf[1440] = 256'hb0f692f694f6a6f6cdf606f737f75ff77bf778f760f73af702f7cdf6a8f68ef6;
    inBuf[1441] = 256'h91f6b4f6e9f633f789f7d6f71ef858f876f884f888f87df877f87ef88ff8baf8;
    inBuf[1442] = 256'h00f953f9b9f926fa86fadcfa20fb42fb50fb4ffb41fb38fb3efb51fb7dfbbffb;
    inBuf[1443] = 256'h09fc5bfcaafce6fc13fd2cfd2ffd27fd1afd0bfd07fd12fd2bfd58fd92fdd2fd;
    inBuf[1444] = 256'h1afe61fea2feddfe0bff2eff4eff68ff83ffa9ffdaff1d007500d5003a01a101;
    inBuf[1445] = 256'hf8013f0275029402a802bd02d302f7022f037103bf030f044e047c0497049504;
    inBuf[1446] = 256'h860473045f045b0467047e04a104c704e104f504fb04f004e504da04cd04cc04;
    inBuf[1447] = 256'hd104d604e204eb04ee04f604fc0404051a05360555057f05a405bc05d005d605;
    inBuf[1448] = 256'hd005ce05cd05d305f005170644067d06ad06cd06e306e306cb06ae0686065a06;
    inBuf[1449] = 256'h39061e06080603060006fe0508060b060506fd05e505b70580053805e804a204;
    inBuf[1450] = 256'h65043f043d0451047804af04dc04f204ef04c20472041404aa0348030403de02;
    inBuf[1451] = 256'hdd02ff022b0358037e03830367033403e5028a023202e0019f0177015d015501;
    inBuf[1452] = 256'h5e01640169016c015d0143011c01e400a60064001c00ddffabff82ff6dff66ff;
    inBuf[1453] = 256'h63ff67ff65ff52ff36ff0affd1fe9afe65fe35fe18fe07fef9fdf5fdedfddbfd;
    inBuf[1454] = 256'hc3fd9efd6dfd3efd0cfddbfcb6fc95fc76fc64fc4efc33fc1bfcf7fbcafb9dfb;
    inBuf[1455] = 256'h60fb1bfbd9fa91fa4dfa1dfaf6f9e1f9e7f9f2f9fff90efa05fae7f9bcf974f9;
    inBuf[1456] = 256'h22f9daf892f85df84cf84bf85ff88cf8b0f8ccf8e4f8daf8b7f88cf843f8f3f7;
    inBuf[1457] = 256'haff766f72bf70ff7fcf6fff620f73df761f78bf797f78cf76ff727f7ccf66ef6;
    inBuf[1458] = 256'h03f6abf579f559f55ef587f5aef5dbf505f608f6f6f5d2f58bf541f5fff4b8f4;
    inBuf[1459] = 256'h89f477f46bf479f4a0f4c2f4f3f42af54bf568f57df56df552f531f5f9f4ccf4;
    inBuf[1460] = 256'hb1f497f49bf4bdf4ddf407f533f53cf533f51bf5e2f4a9f47ef455f448f458f4;
    inBuf[1461] = 256'h66f47df496f492f482f46bf441f422f41bf41df43cf474f4a7f4dcf409f513f5;
    inBuf[1462] = 256'h0ef501f5e1f4cff4d4f4e1f40bf54bf584f5c3f500f624f647f66af67ff69ef6;
    inBuf[1463] = 256'hc7f6e5f607f729f738f74af760f770f792f7caf706f853f8a8f8e8f81bf93cf9;
    inBuf[1464] = 256'h38f925f90ff9f2f8e9f8f8f813f947f98ef9ccf90afa45fa6efa90faaefabffa;
    inBuf[1465] = 256'hd2fae8faf5fa08fb21fb38fb5efb96fbd8fb2efc91fcf2fc4cfd90fdaffdb3fd;
    inBuf[1466] = 256'h9bfd6ffd4bfd3cfd47fd7cfdd2fd38fea4fefdfe34ff4cff41ff1efffcfee6fe;
    inBuf[1467] = 256'he4fe06ff42ff91ffecff3e008400be00e300fd0017012e014b0172019901c601;
    inBuf[1468] = 256'hf701220252028702b902f3022f035e038903a803ae03ad03a903a303b603e003;
    inBuf[1469] = 256'h18046c04cb0417055a05820583057a056a0552055a058105b90515067e06da06;
    inBuf[1470] = 256'h3a078907b407dc07fc070b082a0855087d08bd0803093f098c09da091a0a6f0a;
    inBuf[1471] = 256'hc80a150b6e0bbe0bf20b240c430c460c570c6b0c7c0cb10cf60c380d8f0dde0d;
    inBuf[1472] = 256'h120e480e670e660e6d0e690e520e510e4d0e3f0e4b0e570e5e0e860eb20ed70e;
    inBuf[1473] = 256'h140f4a0f670f8a0f920f790f6d0f590f3d0f4b0f690f920fe40f36107510bc10;
    inBuf[1474] = 256'he810ed10f410e810ca10c810c510bb10d110e210e010f110f510e910f6100011;
    inBuf[1475] = 256'hfe1016111f110e110711e710ad1088105f103610351039103b105a1067105710;
    inBuf[1476] = 256'h50103010f70fd50fae0f860f830f7e0f6f0f780f6e0f4d0f400f290f090f0e0f;
    inBuf[1477] = 256'h170f1d0f3d0f4b0f410f420f290ffa0ee70ed30ec00ed40ee60eeb0eff0ef80e;
    inBuf[1478] = 256'hd00eb00e7d0e3f0e250e0f0efb0d060e050eeb0dd60da70d5b0d200de10ca40c;
    inBuf[1479] = 256'h910c870c7d0c8f0c930c7f0c730c530c1f0c040ce80bcb0bd10bd50bcf0bdc0b;
    inBuf[1480] = 256'hda0bca0bcf0bd10bd40bfb0b210c3d0c640c6e0c540c360cff0bbd0b9c0b8a0b;
    inBuf[1481] = 256'h8d0bbb0bed0b140c3b0c3a0c0e0cd80b880b2f0bf30ac60aac0ab60ac10ac20a;
    inBuf[1482] = 256'hc40aa90a750a440a0b0ad609be09ab099e09a009900969093d09fe08b6087f08;
    inBuf[1483] = 256'h51083608390840084808530846082208f907c0077e0746070b07d606aa067406;
    inBuf[1484] = 256'h3c060706c505840552052005f404d204a5046e042904c9035d03ed0276021002;
    inBuf[1485] = 256'hc401870164015501440137012101f700c400890042000400c8ff82ff43fffffe;
    inBuf[1486] = 256'haefe62fe16fecffda1fd84fd70fd6dfd60fd3bfd01fd9efc14fc7dfbd7fa38fa;
    inBuf[1487] = 256'hbdf95ef923f912f909f900f9f4f8c5f878f818f896f707f783f6fdf584f52af5;
    inBuf[1488] = 256'hd9f49cf47cf45af442f440f434f426f421f405f4ddf3b9f380f346f322f3fcf2;
    inBuf[1489] = 256'heaf2fef218f341f380f3aef3d5f3fbf302f4fdf3fbf3def3bcf3a6f37af34ff3;
    inBuf[1490] = 256'h32f309f3edf2ecf2e5f2eef20cf314f31af31df3f7f2c5f293f246f207f2e5f1;
    inBuf[1491] = 256'hc0f1b8f1d1f1e1f101f22af233f23ff250f243f240f24df247f252f269f268f2;
    inBuf[1492] = 256'h6ff27ef274f279f291f29cf2bef2f1f211f336f35af35df35ff360f347f339f3;
    inBuf[1493] = 256'h38f328f325f32cf323f321f323f313f30ef317f317f327f344f352f364f371f3;
    inBuf[1494] = 256'h64f353f341f321f313f321f33bf37bf3daf33cf4aef422f57bf5cdf512f639f6;
    inBuf[1495] = 256'h60f68cf6aef6e4f62cf773f7d1f73ff8a4f813f981f9d4f91dfa52fa5bfa50fa;
    inBuf[1496] = 256'h34fafef9d1f9b2f996f998f9b2f9d0f9f9f91bfa21fa17faf6f9b2f968f922f9;
    inBuf[1497] = 256'hddf8b1f8a3f8a6f8c2f8e8f805f91df929f91ef909f9f1f8d5f8c4f8c1f8c8f8;
    inBuf[1498] = 256'hdef801f926f955f98af9b8f9e3f909fa22fa31fa32fa26fa1dfa1bfa1efa37fa;
    inBuf[1499] = 256'h6afaa9faf5fa43fb7ffba6fbaefb8efb56fb11fbc6fa93fa82fa91faccfa2afb;
    inBuf[1500] = 256'h93fb00fc62fca5fcd0fce2fcddfcd7fcd9fce6fc10fd53fda4fd09fe7cfef0fe;
    inBuf[1501] = 256'h67ffdaff3e009600d900010113010e01f300cf00ac00900088009500b400e600;
    inBuf[1502] = 256'h1e014f0172017b0166013601f0009c004a000200cdffb1ffadffbbffd8fffcff;
    inBuf[1503] = 256'h23004a006e008a009f00ab00b000ae00a700a400aa00bd00e2001b016101b201;
    inBuf[1504] = 256'h07025902a402e40217034003610377038c039e03a703a803a30394037e036703;
    inBuf[1505] = 256'h510349034e035c0374038e039c03970378033b03e80287022202cd0195017b01;
    inBuf[1506] = 256'h8301a501d601100244026a0284028e02860276025f02420225020902f301ea01;
    inBuf[1507] = 256'hed01fd011e024b027b02aa02ca02d102c0028f023f02dd0172010801b0006f00;
    inBuf[1508] = 256'h490043004f0064007c008b00890076004c001200d2ff8dff48ff0cffe0fec7fe;
    inBuf[1509] = 256'hc8fee1fe0dff4bff91ffd3ff0c003100410042003500220018001d0032005b00;
    inBuf[1510] = 256'h9400d7001a0156018801ad01c301ce01d001ca01be01ad019601770149011001;
    inBuf[1511] = 256'hd000890042000200c7ff90ff5fff2bfff1feb1fe67fe16fec7fd77fd2dfdedfc;
    inBuf[1512] = 256'hb1fc7dfc52fc2afc07fcf3fbedfbf6fb15fc3ffc70fca4fccafcdffce2fccffc;
    inBuf[1513] = 256'haefc8dfc70fc63fc74fc9cfcdafc2cfd82fdd3fd15fe3cfe4bfe46fe2cfe05fe;
    inBuf[1514] = 256'hdffdb8fd9afd8efd8ffda2fdc8fdf8fd2ffe66fe8bfe9cfe96fe6cfe2afedefd;
    inBuf[1515] = 256'h89fd43fd1bfd0cfd20fd54fd90fdd1fd0afe25fe2cfe1ffef7fdccfda8fd88fd;
    inBuf[1516] = 256'h7bfd7ffd87fd97fdaafdadfdaafda0fd85fd65fd41fd12fde4fcb5fc7afc3efc;
    inBuf[1517] = 256'h05fcc8fb90fb62fb35fb11fbeffac4fa96fa67fa2ffafdf9d7f9bdf9b8f9c6f9;
    inBuf[1518] = 256'hdef9fef91ffa35fa40fa40fa34fa2bfa2cfa34fa4efa7dfabafa06fb59fba8fb;
    inBuf[1519] = 256'hfbfb49fc89fcc3fcf4fc15fd2efd3dfd3cfd3cfd3efd41fd58fd86fdc2fd13fe;
    inBuf[1520] = 256'h6cfeb4fee9fefefee1fe9efe3dfec5fd58fd04fdccfcc5fcebfc2dfd83fdd9fd;
    inBuf[1521] = 256'h19fe3ffe43fe1efedffd91fd39fdeefcbdfca9fcbafcecfc38fd96fdf9fd55fe;
    inBuf[1522] = 256'ha3fed9fef3fef2fed9feb3fe88fe61fe4bfe4afe5cfe81feb3feeafe23ff58ff;
    inBuf[1523] = 256'h83ffa6ffc1ffd0ffd4ffd1ffbfffa1ff7bff4eff26ff0eff09ff22ff5cffadff;
    inBuf[1524] = 256'h0d007400ca00040123011e01fc00cd009e0081008600ab00f3005f01d8015602;
    inBuf[1525] = 256'hd2023b039103d303fb03150425042b04300438043f04500469048304a804d504;
    inBuf[1526] = 256'h0305380568058805a305ab059705770548050805cd0494045f04450440044b04;
    inBuf[1527] = 256'h7904bc0406056205ba05fd05360654064e063e0622060006f705080634069106;
    inBuf[1528] = 256'h1107a2074c08f4088109f609410a570a4e0a290aed09bf09a2099a09c0090a0a;
    inBuf[1529] = 256'h6a0ae50a620bc70b160c380c1e0cda0b6e0be00a570adb0978094d094e096b09;
    inBuf[1530] = 256'had09f309200a3c0a2f0af509aa094909df0893085d083d084d087308a008e008;
    inBuf[1531] = 256'h150936095809660963096f0978097e099709ab09b309c309c009a90998097a09;
    inBuf[1532] = 256'h5409420932092509350949095a0977098309770965093909f208af0866082208;
    inBuf[1533] = 256'hfc07e907ec0715084a088008c408f908140923091809f408cd089d086c085308;
    inBuf[1534] = 256'h450846086c089f08d80826097009ab09de09f209e509c40982092709cf087108;
    inBuf[1535] = 256'h1c08eb07ce07c407da07f207ff070608e807a6074c07d0064206c1054605e104;
    inBuf[1536] = 256'ha804870480049704b004c604e004e404d704c804a904870471045c0454046304;
    inBuf[1537] = 256'h73048604a804c204d304e804f50403051805280538054e05570553054a052c05;
    inBuf[1538] = 256'hfc04c9048b0449041204e503c903c303c603ce03d903d303b8038c034703f102;
    inBuf[1539] = 256'h97023b02e701a70177015b015701600175019601b301ca01db01dc01d201bf01;
    inBuf[1540] = 256'h9f017c015c013c0125011e012201380160018f01c401f701170223021702e801;
    inBuf[1541] = 256'ha0014801e30082003000edffc6ffb9ffbfffd5fff1ff01000100eaffb1ff61ff;
    inBuf[1542] = 256'hfdfe90fe2bfed7fd9bfd7ffd84fd9efdc9fdfbfd28fe4bfe59fe51fe37fe0ffe;
    inBuf[1543] = 256'hddfdacfd82fd65fd59fd5afd65fd79fd8dfd9ffdaafda8fd99fd80fd58fd27fd;
    inBuf[1544] = 256'hf6fcc0fc8dfc62fc3bfc18fcfcfbdcfbbcfb9afb6dfb3efb12fbe4fabbfa9dfa;
    inBuf[1545] = 256'h83fa6efa61fa4ffa3bfa26fa0afaeaf9d0f9b8f9acf9b5f9cbf9f3f92ffa71fa;
    inBuf[1546] = 256'hb4faf8fa30fb59fb76fb7ffb7afb72fb66fb62fb6cfb85fbb1fbf0fb36fc7efc;
    inBuf[1547] = 256'hc6fcfdfc20fd2dfd20fd01fdd4fc9cfc6cfc49fc34fc37fc54fc80fcb9fcfbfc;
    inBuf[1548] = 256'h31fd5afd6ffd67fd48fd16fdcffc86fc46fc0cfcebfbedfb06fc3afc83fcc9fc;
    inBuf[1549] = 256'h05fd31fd35fd19fde6fc95fc39fce5fb97fb64fb57fb63fb8cfbcefb0ffc44fc;
    inBuf[1550] = 256'h6cfc71fc55fc22fcd4fb7bfb2cfbe5fab3faa3faadfad0fa0bfb4dfb8ffbcefb;
    inBuf[1551] = 256'hf8fb0dfc10fcfcfbdefbc5fbb1fbaefbc2fbe6fb19fc5bfc9afcd4fc09fd2cfd;
    inBuf[1552] = 256'h41fd50fd4efd47fd45fd40fd3ffd46fd46fd48fd4bfd41fd37fd34fd2afd27fd;
    inBuf[1553] = 256'h30fd33fd39fd40fd36fd22fd08fdd8fca1fc6afc26fcecfbc6fba3fb91fb98fb;
    inBuf[1554] = 256'ha2fbb4fbc9fbc8fbb9fb9cfb64fb1efbd7fa8bfa4cfa26fa0ffa12fa32fa58fa;
    inBuf[1555] = 256'h83faaffac8fad0fac8faaafa83fa5cfa33fa15fa0afa08fa17fa39fa60fa8efa;
    inBuf[1556] = 256'hc2faeffa1afb40fb57fb65fb68fb5bfb4cfb3ffb2ffb2ffb43fb65fb9dfbe8fb;
    inBuf[1557] = 256'h33fc82fccafcf7fc12fd18fd00fde1fcbffc99fc84fc86fc93fcb8fcedfc22fd;
    inBuf[1558] = 256'h5cfd94fdb6fdcffdd9fdcefdbcfda4fd82fd69fd59fd4efd55fd69fd84fdadfd;
    inBuf[1559] = 256'hdffd10fe45fe76fe9bfebafec8fec4feb5fe9cfe79fe58fe3dfe30fe3bfe5cfe;
    inBuf[1560] = 256'h92fedffe36ff88ffcaffedffedffcaff86ff30ffdcfe97fe70fe74fea2fef4fe;
    inBuf[1561] = 256'h63ffdbff4a00a200d600e200ca0094004d000700ccffa8ffa8ffc9ff06005d00;
    inBuf[1562] = 256'hc3002a018c01de01120228021c02f201b40167011b01e400c800ca00f1003601;
    inBuf[1563] = 256'h8b01e4013002650277025c021902b9014101c3004e00eeffabff8cff90ffafff;
    inBuf[1564] = 256'hdeff110040005d005b003e000400b3ff54fff6fea6fe70fe58fe62fe8dfed0fe;
    inBuf[1565] = 256'h22ff78ffc5ff06003600510058004e0037001a00fbffdfffd0ffd2ffe7ff1600;
    inBuf[1566] = 256'h5d00b40014017201c101f7010502eb01b0015b01fe00aa006d0053005e008600;
    inBuf[1567] = 256'hc40007013e015c0156012c01e6008b002900d1ff8fff67ff59ff60ff76ff92ff;
    inBuf[1568] = 256'ha8ffb1ffb1ffa6ff92ff7dff6bff5fff59ff59ff5aff57ff4dff38ff19fff2fe;
    inBuf[1569] = 256'hc6fe9dfe81fe73fe77fe8efeb2fedafefcfe0dff05ffe5feadfe65fe1cfedefd;
    inBuf[1570] = 256'hb4fdaafdbdfdedfd33fe80fec9fe06ff2cff3aff36ff23ff0bfff7feebfeecfe;
    inBuf[1571] = 256'hfafe10ff33ff5fff91ffcdff110057009e00e100150136013a012001f400b700;
    inBuf[1572] = 256'h73003c001b0014002d005f009e00e00014012b012401f4009f003500c0ff48ff;
    inBuf[1573] = 256'hdffe90fe5efe4dfe58fe78fea8fedafe00ff18ff1dff0affe0fea6fe62fe1efe;
    inBuf[1574] = 256'he4fdbafda6fdacfdcbfd00fe46fe90fed8fe17ff46ff60ff62ff4cff22ffecfe;
    inBuf[1575] = 256'haffe77fe4efe3dfe49fe74feb7fe0fff6fffc8ff0f00380040002800f3ffadff;
    inBuf[1576] = 256'h69ff30ff0bff07ff20ff54ff9ffff4ff48009600d100f50006010201e900c400;
    inBuf[1577] = 256'h9600630035001000f7fff9ff16004b009500ed0043018b01b501b80194014901;
    inBuf[1578] = 256'hdf006a00f8ff96ff51ff34ff3cff61ff97ffd2ff050020001900f2ffb2ff5dff;
    inBuf[1579] = 256'hfefea2fe55fe1ffe02fe00fe1afe48fe85fecbfe11ff50ff86ffaaffc1ffcbff;
    inBuf[1580] = 256'hc6ffb8ffa8ff97ff8aff87ff8effa6ffd2ff0f005f00c10029018f01e9012b02;
    inBuf[1581] = 256'h4e024e022802e8019d0152011a01060119015801be013902b70224036c038203;
    inBuf[1582] = 256'h6403110399020c027c010001a60077007a00a800f5005601b9010b0241024f02;
    inBuf[1583] = 256'h3102ec01890111019a003300ebffd2ffe6ff23008300f8006c01d10117023302;
    inBuf[1584] = 256'h2602f00199013701d10073003300180021005300ab001b01990113027c02cb02;
    inBuf[1585] = 256'hf202e902bf0278021a02bf017901510158019001ef016a02ed026103bf03f303;
    inBuf[1586] = 256'hf303cc0387032b03cf028102480232023f026802ac0201035c03ba030b044304;
    inBuf[1587] = 256'h690473045b042d04ee03a3035f032803030301031c034d039603e0031a044504;
    inBuf[1588] = 256'h50043304fe03b30359030403b8027c025f025d027002a102df021e0362039a03;
    inBuf[1589] = 256'hb803c403b6038e035c032103e702c302b002af02ca02f3021f034f0377039003;
    inBuf[1590] = 256'ha103a5039e039a0394038d038e038e038a038a03880386039103a303bf03ea03;
    inBuf[1591] = 256'h190444046d0485048604780457042704f703c8039f0387037b0375037c038603;
    inBuf[1592] = 256'h8d039b03a703ae03bb03c203be03b903a803870362033a031103f702e902eb02;
    inBuf[1593] = 256'h0b03370366039c03c803df03e503d103a4036c032703dc02a0026d0249024102;
    inBuf[1594] = 256'h4c0267029602c602f4021d03300327030a03d20289024002fa01c601b201b601;
    inBuf[1595] = 256'hd4010d024c028a02c202e502ef02e802cb029c0265022702eb01bd0199018801;
    inBuf[1596] = 256'h9401b501e80130027d02c002f5020d030203d7028e023402de0192015d014e01;
    inBuf[1597] = 256'h5c017f01b201e40104020f02fe01d5019d0159011301d5009a0066003f001f00;
    inBuf[1598] = 256'h0700feff02001500370063009500c900f00008010e01fd00da00af0080005a00;
    inBuf[1599] = 256'h47004b006a00a100e50031017a01b701de01ec01dc01b40177012d01df009c00;
    inBuf[1600] = 256'h6f005d0068008e00c300fd002d01460143012201e40091003600ddff8fff51ff;
    inBuf[1601] = 256'h24ff07fff8feedfee5fee0fed9fed4fed2fed2fed3fecdfebafe98fe68fe2afe;
    inBuf[1602] = 256'heafdb3fd8ffd89fda1fdd6fd20fe72febefef2fe06fff8fecefe8dfe44fe01fe;
    inBuf[1603] = 256'hd1fdbcfdc5fde6fd1cfe5afe99fed1fefafe11ff17ff0ffffcfee5feccfeb7fe;
    inBuf[1604] = 256'hacfeacfebafed3fef3fe1aff44ff6bff8dffa8ffb8ffc0ffc2ffbcffb5ffa9ff;
    inBuf[1605] = 256'h98ff88ff77ff67ff5fff5fff6aff83ffa6ffccfff2ff0a000e00ffffd7ff9bff;
    inBuf[1606] = 256'h57ff15ffe1fec2feb9fec7fee6fe08ff21ff2eff29ff0fffe5feb6fe8cfe6ffe;
    inBuf[1607] = 256'h61fe61fe6efe83fe9afeadfebdfec7fecdfed2fed4fed6fed9fedcfeddfedffe;
    inBuf[1608] = 256'he0fee2fee4fee5fee9fef0fef4fef7fefafefbfefbfefefe01ff0dff22ff3aff;
    inBuf[1609] = 256'h54ff6dff7dff85ff83ff76ff66ff59ff4dff48ff4cff55ff63ff70ff76ff79ff;
    inBuf[1610] = 256'h79ff70ff67ff63ff5dff59ff58ff55ff53ff4fff47ff41ff42ff46ff51ff64ff;
    inBuf[1611] = 256'h78ff8aff99ff9cff92ff7fff62ff3eff18fff0fecafeacfe90fe7bfe6ffe63fe;
    inBuf[1612] = 256'h5bfe59fe54fe50fe4bfe3efe29fe0bfee1fdb5fd8dfd68fd55fd59fd6dfd92fd;
    inBuf[1613] = 256'hc0fde6fd02fe0efe03fee5fdb9fd84fd57fd3afd27fd28fd3dfd5bfd7efd9ffd;
    inBuf[1614] = 256'hb6fdc6fdd0fdd0fdcefdd1fdd5fddffdeefdfdfd0ffe24fe36fe46fe57fe64fe;
    inBuf[1615] = 256'h72fe81fe8afe91fe98fe9afe99fe95fe89fe78fe62fe42fe1ffefefdddfdc3fd;
    inBuf[1616] = 256'hb9fdb9fdc5fddcfdf4fd08fe13fe0afef2fdcefda0fd74fd55fd42fd43fd5afd;
    inBuf[1617] = 256'h7cfda4fdcdfde9fdf6fdf3fddafdb9fd96fd6ffd51fd42fd3bfd41fd54fd68fd;
    inBuf[1618] = 256'h82fda1fdbbfdd4fdeffd00fe0ffe1afe1bfe19fe1afe18fe1bfe28fe35fe47fe;
    inBuf[1619] = 256'h5ffe6ffe79fe7dfe71fe5dfe44fe1efef5fdcffda5fd82fd6bfd55fd47fd44fd;
    inBuf[1620] = 256'h44fd4afd55fd5afd5dfd5cfd50fd3efd29fd0efdfbfcf3fcf3fcfefc14fd28fd;
    inBuf[1621] = 256'h3cfd46fd3dfd25fd03fdd6fcaafc86fc69fc60fc6bfc7dfc97fcb6fccbfcd9fc;
    inBuf[1622] = 256'he1fcdbfcd1fcc9fcc0fcc2fcd0fce0fcf8fc17fd2ffd41fd50fd4ffd44fd33fd;
    inBuf[1623] = 256'h18fdfcfce4fcc8fcb2fca6fc97fc8cfc89fc82fc7bfc7afc75fc70fc74fc77fc;
    inBuf[1624] = 256'h81fc94fca4fcb5fcc6fcc9fcc5fcbefcabfc98fc8cfc83fc85fc94fca2fcb2fc;
    inBuf[1625] = 256'hc1fcc0fcb4fc99fc6afc39fc0cfce3fbccfbcffbe5fb0ffc46fc79fcacfcd2fc;
    inBuf[1626] = 256'hdefcdafccafcaafc88fc6efc5afc58fc69fc84fcacfcdafc01fd21fd35fd34fd;
    inBuf[1627] = 256'h27fd12fdeffccdfcb3fca1fc9cfcabfcc6fceefc1dfd46fd6dfd8efd9efda3fd;
    inBuf[1628] = 256'ha4fd9dfd94fd8ffd8afd8dfd97fda3fdb5fdccfdddfdeefd01fe0efe1bfe28fe;
    inBuf[1629] = 256'h31fe3bfe46fe4cfe53fe5cfe64fe72fe84fe97feb1fed3fef3fe13ff34ff54ff;
    inBuf[1630] = 256'h71ff85ff90ff98ff9aff91ff86ff7dff74ff6fff6eff71ff7bff89ff95ffa2ff;
    inBuf[1631] = 256'hadffb1ffaeffa2ff8cff73ff59ff3eff28ff1eff1eff2bff40ff5bff7aff97ff;
    inBuf[1632] = 256'hadffbeffc6ffc2ffb8ffabff9fff97ff98ffa2ffb6ffd3fff9ff24004d007000;
    inBuf[1633] = 256'h8e00a300ae00b000ac00a700a500a800b300c600df00020129014a0168018101;
    inBuf[1634] = 256'h8e0191018c017e01710165015c015b015f01640170017d0185018c0190018e01;
    inBuf[1635] = 256'h8b0185017e017c017c017e018a019701a301b201c001c701d001d301d101d301;
    inBuf[1636] = 256'hd401d301db01e801f90111022602370247024e02490241023502290228022e02;
    inBuf[1637] = 256'h3b02550274029502b902d202e002e802e202d102c002ad029e029b02a102ac02;
    inBuf[1638] = 256'hc202d702e802fb0208030b030903fe02ec02e102d502c802c802d202de02f502;
    inBuf[1639] = 256'h0f0325033c034a034e0355035303460340033a033203340339033b0343034703;
    inBuf[1640] = 256'h45034803470342034a03570365037f039903ac03c403d403d603d603d003c303;
    inBuf[1641] = 256'hbf03be03c003d403ec03030421043a0445044a04400427040c04ec03c803b103;
    inBuf[1642] = 256'ha503a303b803d703fc032c0454046e04810482046e04550433040d04f403e203;
    inBuf[1643] = 256'hd803e403f8030f042c043d043d04390429040a04e903c603a3038f0382037803;
    inBuf[1644] = 256'h80039103a403c503e503ff031d0433043b043f043a042a041d040e04fd03f803;
    inBuf[1645] = 256'hfb0302041504270432043f04440439042e041f040a04fa03ed03e003e003e703;
    inBuf[1646] = 256'hed03fa0305040904120418041504160416041104110412040a040404f903e603;
    inBuf[1647] = 256'hd603c103a2038c0379036503600365036c0380039503a003a903a70395038103;
    inBuf[1648] = 256'h68034d0341033e0342035c037e039e03bf03d403d603cd03b3038b0366034503;
    inBuf[1649] = 256'h28031e031d03220332033e033e033b0330031d030c03fa02e902e602e902ef02;
    inBuf[1650] = 256'h000312031e032b0330032b03240319030b03070307030b031a032c033e035103;
    inBuf[1651] = 256'h5a03560349032f030c03e802c402a30295029802ab02ce02f7021e0341035303;
    inBuf[1652] = 256'h500340031f03f302ca02a6028c0286029102a702c902ec02070319031a030503;
    inBuf[1653] = 256'he302b10276023f021002eb01dc01e101f501190243026b028c029e029d029002;
    inBuf[1654] = 256'h76025102300219020b020d021a022f024b02620270027602700260024d023402;
    inBuf[1655] = 256'h19020202ec01d801cd01c301b801b401b301b501b901c001cc01de01eb01f201;
    inBuf[1656] = 256'hf501ef01df01ca01af0194017c0169015c01570156015c016501690169016601;
    inBuf[1657] = 256'h58013f011f01fa00d700b700a100970098009f00ae00c000cd00d400d300c800;
    inBuf[1658] = 256'hb3009700760057003b00230010000000f4ffecffe3ffd8ffceffc7ffbeffb5ff;
    inBuf[1659] = 256'haeffa5ff98ff87ff74ff63ff52ff43ff3dff3eff46ff54ff65ff75ff82ff87ff;
    inBuf[1660] = 256'h87ff81ff75ff66ff58ff4cff43ff3fff3eff3dff3fff40ff3eff3cff37ff32ff;
    inBuf[1661] = 256'h30ff2cff28ff25ff21ff18ff0dff00fff3fee7fedafed0fecdfecbfec9fecbfe;
    inBuf[1662] = 256'hcefecefecbfec3feb7fea9fe95fe7cfe66fe52fe41fe3afe38fe3bfe44fe4efe;
    inBuf[1663] = 256'h55fe58fe51fe41fe2ffe18fe01feeffde1fddcfde3fdebfdf1fdfafdfcfdf6fd;
    inBuf[1664] = 256'hecfddbfdc8fdbafdaffdaafdaffdb6fdbffdccfdcffdccfdc6fdb9fda7fd98fd;
    inBuf[1665] = 256'h8afd84fd88fd90fda0fdb4fdc1fdccfdd6fdd2fdc2fdaffd98fd82fd70fd5ffd;
    inBuf[1666] = 256'h5afd62fd6dfd7dfd91fd9cfd9efd98fd84fd68fd48fd24fd06fdf3fce6fce4fc;
    inBuf[1667] = 256'heefcf8fc05fd10fd10fd06fdf7fcdcfcbefca2fc87fc74fc6cfc67fc67fc6dfc;
    inBuf[1668] = 256'h6ffc71fc74fc70fc6bfc68fc5dfc54fc51fc4dfc4bfc4cfc4cfc4dfc50fc4bfc;
    inBuf[1669] = 256'h46fc44fc3cfc34fc2ffc27fc20fc1efc19fc16fc17fc13fc0efc0cfc03fcf9fb;
    inBuf[1670] = 256'hf4fbe9fbe3fbe5fbe6fbebfbf5fbfbfb02fc0bfc09fc04fc00fcf4fbe8fbdefb;
    inBuf[1671] = 256'hd0fbc6fbc2fbb8fbaffbadfba7fba3fba5fba3fba2fba5fb9ffb99fb93fb85fb;
    inBuf[1672] = 256'h79fb75fb6cfb68fb6bfb6ffb7dfb90fb9afba5fbb1fbb2fbaffba9fb99fb8afb;
    inBuf[1673] = 256'h80fb75fb6ffb70fb6efb74fb80fb88fb93fba1fba6fbaafbb1fbb0fbaffbb0fb;
    inBuf[1674] = 256'hadfbadfbb2fbb5fbc0fbd1fbdefbeffb04fc11fc19fc1dfc1bfc19fc14fc09fc;
    inBuf[1675] = 256'h01fcfefbf9fbf8fbfefb02fc0bfc1bfc28fc37fc49fc57fc65fc73fc7afc82fc;
    inBuf[1676] = 256'h8bfc8afc88fc8cfc8ffc96fca3fcb0fcc2fcdafcecfcfafc04fd03fdfffcf7fc;
    inBuf[1677] = 256'he3fccdfcbdfcabfc9ffc9dfc9efca9fcbdfcd2fce9fc00fd0efd17fd1bfd12fd;
    inBuf[1678] = 256'h04fdf7fce7fcdcfcddfce6fcfafc1bfd3efd64fd88fd9efdaafdadfda1fd8dfd;
    inBuf[1679] = 256'h79fd66fd59fd57fd5ffd74fd95fdb9fddffd07fe28fe41fe53fe58fe57fe53fe;
    inBuf[1680] = 256'h4cfe49fe4ffe5cfe72fe8efeadfecffeeffe03ff0cff0eff08fffcfeeefee2fe;
    inBuf[1681] = 256'hdafed8fedefeeafef9fe08ff15ff23ff2fff38ff3fff4bff5cff70ff84ff99ff;
    inBuf[1682] = 256'hacffbcffc4ffc7ffc6ffc1ffbeffbdffbcffc1ffcbffd4ffddffe6ffe9ffe7ff;
    inBuf[1683] = 256'he0ffd3ffc3ffb5ffa9ffa3ffa6ffafffc1ffdbfff8ff16003300490059006100;
    inBuf[1684] = 256'h60005d005a00570059006200710083009900ab00b900c200c400bf00b800b100;
    inBuf[1685] = 256'haf00b500c500dc00fa001a01380154016701710175017401740178017b017f01;
    inBuf[1686] = 256'h8c019e01b001c101cc01d201d001c301af019a0180016701580150014f015c01;
    inBuf[1687] = 256'h74019201b301cf01e601f601f601ea01dd01cd01c001be01c501d501f0010e02;
    inBuf[1688] = 256'h28023e02470246023f022c021302fd01ea01db01d701d801db01e401ec01f301;
    inBuf[1689] = 256'hfb01fe01fd01ff01fe01fd01020207020b0215021c021f0221021d0216021102;
    inBuf[1690] = 256'h0902000201020602100225023d0253026a0276027702710260024b023b023102;
    inBuf[1691] = 256'h330249026a029402c502f20217032f03330329031603f702d502bf02b302b302;
    inBuf[1692] = 256'hc302dc02fb021c033803490350034b033c0325030803ee02dd02d002cb02d602;
    inBuf[1693] = 256'hec02040320033b035203610363035c0355034b033b0330032a03250325032503;
    inBuf[1694] = 256'h21031f0319030f030803ff02f802f602f402ef02f102ee02e102d402c102a902;
    inBuf[1695] = 256'h97028a0284028d029d02b502d702f5020a031b031f0315030503ea02c902ad02;
    inBuf[1696] = 256'h9502870289029602b002d8020203270349035c035c034e0333031003f002d502;
    inBuf[1697] = 256'hc602cd02e10201032b03550377038f0391037f03620338030703d902b2029602;
    inBuf[1698] = 256'h880284028a029a02ab02b902c602ce02cf02c902b802a00288026e0254024102;
    inBuf[1699] = 256'h3702340238024302520263026f02740275026d025d0246022b020d02f201dd01;
    inBuf[1700] = 256'hce01c801c901d301e401fa010f0226023502390237022a021202f801de01c701;
    inBuf[1701] = 256'hbb01b601b801c401d501e401f001f301ee01e401d301bf01b001a3019b019e01;
    inBuf[1702] = 256'ha401ad01ba01c201c701cf01d201d101d301d101cd01cd01c901c201bc01b101;
    inBuf[1703] = 256'ha7019e0193018a018801850185018801890189018d0191019401970197019901;
    inBuf[1704] = 256'h990192018b0185017a017001680162015d01590154014f0148013c012e012101;
    inBuf[1705] = 256'h11010101f600ed00e500df00db00d800d500d200cd00ca00cb00ce00d200d300;
    inBuf[1706] = 256'hd300d600d500cf00c800c000b400a7009b009100890081007b007a007a007e00;
    inBuf[1707] = 256'h860090009d00ac00b700bc00ba00af009c008700710060005b00610072008e00;
    inBuf[1708] = 256'haa00c300d500d900cb00af00870056002400f7ffd7ffcbffd0ffe4ff02002500;
    inBuf[1709] = 256'h4900630068005e0047002200f5ffc7ff9eff82ff78ff7dff94ffb5ffd9fffaff;
    inBuf[1710] = 256'h110016000900ecffc4ff97ff6aff43ff2bff1eff1dff28ff36ff44ff53ff5eff;
    inBuf[1711] = 256'h62ff62ff60ff59ff52ff4aff40ff35ff2aff20ff17ff0fff0dff14ff21ff32ff;
    inBuf[1712] = 256'h4aff62ff73ff7cff7bff6dff52ff2eff09ffe7fec8feb3feaefeb4fec3fedcfe;
    inBuf[1713] = 256'hfbfe1bff36ff46ff4aff3eff22fffdfed7feb3fe95fe87fe88fe99feb4fed3fe;
    inBuf[1714] = 256'hf1fe08ff11ff0cfff6fed0fea4fe77fe4efe32fe28fe2afe38fe50fe6cfe88fe;
    inBuf[1715] = 256'ha2feb6fec5fed0fed7fedafed9fed3fecdfec7febdfeb6feb5feb6febafec5fe;
    inBuf[1716] = 256'hd1fedafee1fee3fedffed4febffea4fe8afe6dfe50fe39fe29fe22fe27fe37fe;
    inBuf[1717] = 256'h50fe70fe8ffeacfec2fecbfec9febcfea2fe7ffe60fe44fe31fe2efe39fe51fe;
    inBuf[1718] = 256'h72fe91fea9feb7feb6fea8fe91fe73fe5afe4dfe47fe4efe65fe83fea8feccfe;
    inBuf[1719] = 256'he8fe01ff14ff18ff18ff12ff04fff9fef2fee8fee5fee7fee4fee4fee5fee1fe;
    inBuf[1720] = 256'hddfed7fecbfec3febdfeb7feb9febffec5fed4fee3feeffefcfe02ff00fffffe;
    inBuf[1721] = 256'hfcfef6fef7fe00ff0cff1eff31ff3dff44ff46ff3dff2fff1eff0cfffefef3fe;
    inBuf[1722] = 256'heafee7fee6fee6fee9feecfeeffef4fefafefefe05ff0bff0eff13ff16ff12ff;
    inBuf[1723] = 256'h0cff08ff01fffbfef8fef7fefdfe09ff14ff20ff2cff30ff32ff31ff2bff27ff;
    inBuf[1724] = 256'h24ff1aff10ff08ff00ff00ff02ff07ff1bff38ff53ff6fff87ff94ff9aff96ff;
    inBuf[1725] = 256'h85ff72ff5cff45ff38ff31ff30ff3dff51ff68ff84ff9dffadffb6ffb6ffa9ff;
    inBuf[1726] = 256'h95ff78ff57ff39ff1fff0cff0bff1bff39ff65ff99ffcafff2ff0a000d00faff;
    inBuf[1727] = 256'hd5ffa8ff7aff53ff3dff3cff4cff6bff94ffbcffdcfff1fff6ffeeffd9ffb8ff;
    inBuf[1728] = 256'h92ff6fff53ff40ff36ff38ff42ff54ff6cff85ff9bffafffc0ffc8ffcaffc8ff;
    inBuf[1729] = 256'hbcffa6ff8fff7aff66ff58ff52ff54ff5dff6dff82ff9cffb7ffd2ffe7fff5ff;
    inBuf[1730] = 256'hf9ffeeffd7ffb8ff96ff77ff64ff60ff72ff9cffd2ff0d00470073008d008d00;
    inBuf[1731] = 256'h740048001400ddffb2ff9aff97ffacffd5ff07003a00680085008e0084006800;
    inBuf[1732] = 256'h46002100ffffe4ffd6ffd3ffdcffefff070020003600470050004c003f002b00;
    inBuf[1733] = 256'h1300fcffe9ffdcffd8ffdfffebfffaff0600100018001b001d00220026002b00;
    inBuf[1734] = 256'h320038003b003a003200260018000700f8fff1fff1fff9ff08001b002e003b00;
    inBuf[1735] = 256'h40003f00360028001a000e0009000b00100015001d00230028002f0034003700;
    inBuf[1736] = 256'h3900390035002c001f0012000500fafff3fff1fff3fffbff0700110019001f00;
    inBuf[1737] = 256'h240024002300230027002f0037003e00440046003f00310020000900f3ffe8ff;
    inBuf[1738] = 256'he4ffe7fff4ff02000f00180016000b00fbffe5ffcfffbdffaeffa5ffa4ffaaff;
    inBuf[1739] = 256'hb7ffc9ffdefff7ff0c00190020001f001000f7ffdbffbbff9fff89ff7bff78ff;
    inBuf[1740] = 256'h81ff92ffa6ffb9ffcaffd1ffc9ffb7ffa1ff88ff70ff60ff56ff53ff56ff5aff;
    inBuf[1741] = 256'h5eff63ff69ff70ff78ff82ff8eff96ff96ff8fff7eff61ff3fff1dfffefee7fe;
    inBuf[1742] = 256'hdffee3fef4fe0fff2dff47ff61ff73ff78ff71ff61ff4bff34ff1dff0bff01ff;
    inBuf[1743] = 256'h01ff0dff23ff3fff60ff85ffa6ffbfffcdffc9ffb2ff8dff5cff29fffffee3fe;
    inBuf[1744] = 256'hdafeeafe09ff32ff5dff7eff97ffa4ff9cff86ff6bff4aff2aff13ff01fffcfe;
    inBuf[1745] = 256'h06ff19ff35ff58ff7aff98ffadffb4ffafff9aff78ff55ff33ff12fffefef8fe;
    inBuf[1746] = 256'hfbfe0cff29ff45ff5dff6cff71ff6eff63ff55ff4eff4dff51ff5bff6aff77ff;
    inBuf[1747] = 256'h7fff7eff79ff76ff74ff74ff7cff88ff94ffa2ffadffb0ffabffa0ff8fff7aff;
    inBuf[1748] = 256'h68ff5bff59ff60ff70ff89ffaaffcdffedff08001c0028002d0029001e001200;
    inBuf[1749] = 256'h0600fdfffafffeff0d00260042005b0071007b0077006900510034001e000f00;
    inBuf[1750] = 256'h0c001a0031004d0069007e008c00940094009300960099009f00aa00b500bc00;
    inBuf[1751] = 256'hbf00bb00b000a100910083007b007c0086009500a500b100b700b700b300a800;
    inBuf[1752] = 256'h9a008f008a008d009500a100b200c200ce00da00e300e800ea00e600de00d600;
    inBuf[1753] = 256'hca00bc00b400b100b200b900c300cf00db00e000df00dd00d600d000d300da00;
    inBuf[1754] = 256'he600fb0010011f012b0130012b0123011501060100010501120125013b014f01;
    inBuf[1755] = 256'h5b015c0152013f0124010901f600ee00ef00fb000c011e01320143014a014c01;
    inBuf[1756] = 256'h4b0144013c01310124011a0112010c010e0115011d012a013a0144014a014a01;
    inBuf[1757] = 256'h43013701280117010d0106010101070113011e012801300132012f0127011c01;
    inBuf[1758] = 256'h160116011a0124012f0135013b013b0135012f012a01260128012b0131013a01;
    inBuf[1759] = 256'h4301490150015301510150014d01470143013b012f0125011f011b011e012201;
    inBuf[1760] = 256'h2c013d014e015c01670166015c014d0136011b010801fb00f600fd000b011f01;
    inBuf[1761] = 256'h3601430149014a01400132012601160107010001fa00f700fc0002010a011801;
    inBuf[1762] = 256'h2901390147014e0151014f014501330120010e01fc00f400f500f90005011301;
    inBuf[1763] = 256'h1d0125012801200116010e010101f700f100e800df00db00d300cc00c800c400;
    inBuf[1764] = 256'hc400c700cd00d600db00d900d600cc00b800a50093007d006f006a006a007000;
    inBuf[1765] = 256'h7a00850092009b00a000a1009d009400870077006500530045003c0036003600;
    inBuf[1766] = 256'h40004f005d00690070006f006600520037001e000a00fdfffbff040016002c00;
    inBuf[1767] = 256'h3f004d00540051004600360028001c0012000f00120016001a001d001e001c00;
    inBuf[1768] = 256'h140009000300fffffafffaff0000060011001d002200230021001b0013000700;
    inBuf[1769] = 256'hfbfff3ffefffeffff3fff9ff000009000c000700fbffe6ffcaffaeff96ff86ff;
    inBuf[1770] = 256'h82ff89ff9dffb7ffd1ffe6fff2fff0ffe4ffd0ffbaffa7ff97ff91ff97ffa4ff;
    inBuf[1771] = 256'hb4ffc6ffd1ffd3ffcdffbdffa9ff97ff84ff75ff6fff71ff77ff82ff8eff98ff;
    inBuf[1772] = 256'h9effa0ff9fff9bff97ff94ff93ff93ff96ffa0ffaaffb3ffbfffc8ffc9ffc7ff;
    inBuf[1773] = 256'hbeffabff9bff90ff88ff85ff8bff96ffa5ffb5ffc2ffc9ffcaffc4ffb9ffacff;
    inBuf[1774] = 256'ha2ff9eff9dffa3ffb3ffc4ffd2ffe2ffebffe8ffe4ffdaffcbffbdffb0ffa5ff;
    inBuf[1775] = 256'h9eff9aff98ff9aff9cff9dffa1ffa3ffa0ff9dff99ff94ff8eff88ff85ff84ff;
    inBuf[1776] = 256'h84ff89ff92ff9affa1ffa7ffa9ffa7ffa1ff99ff93ff8fff8cff8bff90ff99ff;
    inBuf[1777] = 256'ha1ffa5ffa6ffa2ff9cff95ff8aff7eff77ff78ff7dff84ff8fff9cffa9ffb4ff;
    inBuf[1778] = 256'hb9ffbcffbaffb4ffadffa3ff99ff94ff94ff98ffa1ffb0ffbeffcbffd7ffdaff;
    inBuf[1779] = 256'hd7ffceffbdffa9ff9aff8dff83ff85ff8fff9dffafffc4ffd5ffe1ffe2ffddff;
    inBuf[1780] = 256'hd6ffccffc2ffbbffb9ffbdffc5ffceffd6ffdeffe1ffdeffdbffd6ffcfffc9ff;
    inBuf[1781] = 256'hc5ffc1ffc1ffc3ffc3ffc4ffc6ffc5ffc2ffc0ffbbffb8ffbaffc0ffc9ffd6ff;
    inBuf[1782] = 256'he5fff5ff04000d000d000400f6ffe3ffceffbaffabffa5ffa9ffb4ffc6ffdaff;
    inBuf[1783] = 256'hebfff5fff8fff0ffe0ffccffb5ffa1ff95ff92ff9cffb1ffc9ffe5ff03001900;
    inBuf[1784] = 256'h25002a0021000f00faffe3ffcdffc0ffbaffbaffc2ffd0ffe2fff3ffffff0500;
    inBuf[1785] = 256'h0500fffff5ffe8ffdaffd0ffcaffc8ffceffd8ffe3fff1fffdff020003000100;
    inBuf[1786] = 256'hfbfff1ffe6ffdcffd2ffc5ffbdffb9ffb5ffb2ffb1ffafffacffacffaeffafff;
    inBuf[1787] = 256'hafffaeffadffabffa6ffa0ff9bff97ff93ff90ff8cff8bff8aff85ff80ff7eff;
    inBuf[1788] = 256'h76ff6bff63ff5aff50ff48ff41ff3cff3bff39ff35ff37ff37ff34ff30ff2dff;
    inBuf[1789] = 256'h2cff2bff2bff2dff30ff32ff36ff3aff3bff39ff36ff30ff28ff20ff17ff10ff;
    inBuf[1790] = 256'h0dff0cff0fff15ff19ff1eff22ff1eff1aff17ff0eff04fffefef9fef5fef5fe;
    inBuf[1791] = 256'hf8fefbfefbfefcfefdfefbfef5feeefee8fee1fed9fed4fed2fed0fecafec5fe;
    inBuf[1792] = 256'hc3fec0febbfeb9febbfebbfebbfebefec2fec3fec3fec2fec1febcfeb3feabfe;
    inBuf[1793] = 256'ha8fea3fea0fea2fea6feaefeb8febdfebffec1febcfeb4feadfea4fe9dfe97fe;
    inBuf[1794] = 256'h92fe91fe96fe9bfea2feabfeb4febcfec1febffebefebcfeb6feb0feacfea7fe;
    inBuf[1795] = 256'ha7feaafeabfeb1febafec3fecefed7fedefee4fee8fee5fedffedafed4fecdfe;
    inBuf[1796] = 256'hc7fec5fecbfed7fee4fef2fe03ff13ff1eff21ff1dff17ff10ff05fffafef5fe;
    inBuf[1797] = 256'hf5fefbfe07ff12ff1eff2cff34ff35ff32ff28ff1cff11ff07ff01ff03ff0bff;
    inBuf[1798] = 256'h18ff29ff37ff44ff4eff4fff4cff48ff40ff3cff3aff39ff42ff52ff5eff6cff;
    inBuf[1799] = 256'h78ff7dff7eff78ff6dff61ff55ff4eff4fff55ff5fff70ff83ff93ffa0ffa9ff;
    inBuf[1800] = 256'habffa9ffa2ff9aff96ff95ff9affa3ffafffc1ffd6ffe6ffeffff5fff7fff2ff;
    inBuf[1801] = 256'hebffe2ffdaffd8ffd9ffdaffe0ffecfff6ff01000b00110016001c0021002600;
    inBuf[1802] = 256'h2d00370042004900500056005500510051004e00470049004d00510059006400;
    inBuf[1803] = 256'h6f00780079007500710069005c0053004c004b005500640078009300ad00c000;
    inBuf[1804] = 256'hd100d900d700cd00be00ad009f00950090009400a200b600ca00dd00ef00fb00;
    inBuf[1805] = 256'hfe00fa00f300e700d700cb00c600c800d000e000f4000c012401390147014f01;
    inBuf[1806] = 256'h51014b01420139012e0123011f01210125012f013f015001610171017c018401;
    inBuf[1807] = 256'h850181017d0176016e016d017001740182019401a401b801c801d101d901da01;
    inBuf[1808] = 256'hd101c901c101b801b201af01b001ba01c501d001e001ea01ee01f101ee01e801;
    inBuf[1809] = 256'he501e001db01de01e301e901f60102020b02140218021902180214020f020c02;
    inBuf[1810] = 256'h0a020b02110216021d0227022b022e02320231022c022b022702220224022802;
    inBuf[1811] = 256'h2a023002360238023e0242024102440246024202430244024402470248024702;
    inBuf[1812] = 256'h4b024d024a024f025202510259025d025b02600263025f025f025c0253025302;
    inBuf[1813] = 256'h53024e02520255025702600267026b02740275026f026f026c0261025c025802;
    inBuf[1814] = 256'h53025302530254025c026002620268026a02680266025f0255024d0242023802;
    inBuf[1815] = 256'h33022c0227022a02300236023f02440247024b0247023e02330221020d02ff01;
    inBuf[1816] = 256'hf301e901ea01ef01f9010c021a0223022a02260217020602f101da01c601b601;
    inBuf[1817] = 256'hb001b701c001cf01e401f401fe010302fb01ea01d701be01a301910186018101;
    inBuf[1818] = 256'h89019701a701b801c101c101c201b901a50191017c0168015c01550152015801;
    inBuf[1819] = 256'h5e0164016b016c0166015c014d013b012e012201160112011101120117011801;
    inBuf[1820] = 256'h1801190114010c010401fc00f400ed00e600e200df00d900d300cb00be00b400;
    inBuf[1821] = 256'haa009a008c0083007a0073006f006b0066006000580051004b00420037002f00;
    inBuf[1822] = 256'h290024001f001a0016000f000300f8ffecffdcffcbffbeffb2ffa8ffa4ffa3ff;
    inBuf[1823] = 256'h9eff97ff91ff8bff82ff76ff6bff5fff55ff4eff4fff54ff59ff60ff65ff69ff;
    inBuf[1824] = 256'h69ff63ff57ff48ff37ff27ff1aff0dff04ff01ff01ff04ff05ff04ff00fffafe;
    inBuf[1825] = 256'hf0fee4fed6fecafec0feb8feb4feb3feb3feb7febcfebdfebcfebefebbfeb3fe;
    inBuf[1826] = 256'haafe9efe91fe86fe79fe69fe5dfe52fe46fe3afe32fe2cfe28fe24fe23fe23fe;
    inBuf[1827] = 256'h20fe1cfe15fe0dfe05fefdfdf2fde7fde1fddffddffde3fde8fdecfdf0fdf0fd;
    inBuf[1828] = 256'hecfde6fddafdc9fdbbfdacfd9ffd97fd91fd91fd97fd9dfda3fdacfdb1fdb2fd;
    inBuf[1829] = 256'hb3fdadfda7fda1fd9afd95fd95fd91fd91fd97fd9afd9dfda2fda1fda2fda6fd;
    inBuf[1830] = 256'ha2fd9afd95fd8cfd83fd7dfd72fd6bfd69fd65fd65fd69fd69fd6dfd76fd78fd;
    inBuf[1831] = 256'h79fd79fd73fd6cfd67fd5ffd58fd56fd56fd5bfd64fd6bfd74fd7cfd7dfd7bfd;
    inBuf[1832] = 256'h79fd70fd63fd5afd51fd4dfd4efd4cfd50fd5bfd60fd60fd63fd60fd57fd4ffd;
    inBuf[1833] = 256'h47fd3ffd3cfd3afd3ffd47fd4cfd53fd5afd58fd54fd50fd47fd3dfd34fd2cfd;
    inBuf[1834] = 256'h2bfd2efd2ffd34fd3afd3bfd3cfd3bfd32fd2afd26fd1ffd19fd18fd1bfd22fd;
    inBuf[1835] = 256'h2bfd34fd3ffd48fd4cfd4ffd4ffd4cfd4cfd4cfd49fd4afd4efd4ffd51fd52fd;
    inBuf[1836] = 256'h50fd52fd55fd52fd51fd54fd50fd4ffd53fd51fd4ffd50fd4efd4efd4ffd4efd;
    inBuf[1837] = 256'h53fd5cfd63fd6cfd76fd7afd80fd82fd7afd75fd71fd65fd5dfd5afd57fd5cfd;
    inBuf[1838] = 256'h62fd67fd71fd78fd77fd78fd75fd68fd5ffd59fd52fd51fd56fd5cfd68fd79fd;
    inBuf[1839] = 256'h84fd8dfd93fd92fd8cfd84fd7bfd72fd6dfd6dfd73fd7efd89fd94fd9ffda7fd;
    inBuf[1840] = 256'ha8fda6fda1fd98fd93fd8efd8bfd92fd9cfdaafdbdfdcbfdd2fdd9fdd8fdd0fd;
    inBuf[1841] = 256'hc9fdc0fdb9fdb9fdbafdc0fdd0fdddfdeafdf9fdfffd01fe02fefafdf0fdeafd;
    inBuf[1842] = 256'he3fde2fde9fdf1fd01fe14fe1ffe29fe2ffe2cfe27fe20fe16fe10fe0ffe11fe;
    inBuf[1843] = 256'h1bfe27fe34fe46fe54fe5bfe60fe64fe62fe5efe5cfe5dfe64fe6dfe79fe88fe;
    inBuf[1844] = 256'h95fe9efea5fea8fea3fe9afe92fe8afe87fe8afe8efe97fea5feb0feb8fec2fe;
    inBuf[1845] = 256'hc7fec4febffebafeb5feb3feb3feb8fec7fed7fee7fef7fe03ff07ff06fffdfe;
    inBuf[1846] = 256'heefee2fed6feccfecafeccfed4fee3fef4fe02ff0fff16ff18ff18ff14ff0fff;
    inBuf[1847] = 256'h0bff0aff11ff1dff2cff41ff57ff69ff79ff84ff86ff84ff81ff7aff71ff6cff;
    inBuf[1848] = 256'h6eff72ff78ff83ff90ff9cffa5ffadffb2ffb2ffafffadffabffaeffb7ffc1ff;
    inBuf[1849] = 256'hcdffdbffebfff7fffeff02000200fffff9fff2ffebffe7ffe8ffeaffeffff6ff;
    inBuf[1850] = 256'hfbfffdfffdfff8fff0ffe8ffe0ffdaffdaffe1ffedfffdff0c001e002f003900;
    inBuf[1851] = 256'h400042003c0033002c00250025002b0034004200530063007000780076006f00;
    inBuf[1852] = 256'h640055004a00430043004c005d0073008e00a900bc00c800cc00c900c000b600;
    inBuf[1853] = 256'hac00a500a700b100c100d600eb00ff000f01160114010a01fb00ec00e100d800;
    inBuf[1854] = 256'hd800e300f30005011d01340144014d014d0147013f0136013101330139014801;
    inBuf[1855] = 256'h5f0177019001a401b001b801b601ac01a4019b01920192019a01a601bc01d301;
    inBuf[1856] = 256'he401f501000201020002fa01ee01ec01ef01f401020216022a0243025b026902;
    inBuf[1857] = 256'h76027b02770274026e02650266026b026f027e0290029c02aa02b502b802bc02;
    inBuf[1858] = 256'hbb02b602b702ba02b902c202d102df02f4020803160329033c03460353035d03;
    inBuf[1859] = 256'h62036d037803810391039d03a203ae03bc03c203ca03d403da03e503ee03f403;
    inBuf[1860] = 256'hff0308040a0416042204280437044704530465047704830493049e04a404ac04;
    inBuf[1861] = 256'hb004af04b304b404b504bd04c004c304d004d704d504da04dd04db04de04e004;
    inBuf[1862] = 256'he004eb04f8040305190530053f0556056a0574057f0588058905900598059b05;
    inBuf[1863] = 256'ha805b805c205d505e605ed05f905010601060406050602060b0615061c063006;
    inBuf[1864] = 256'h440655067006830689069806a1069e06a406a606a006a906b406b906c706d306;
    inBuf[1865] = 256'hd606e106e606e006e206dd06d106d206d306d106df06eb06f306080717071a07;
    inBuf[1866] = 256'h240728072007230724071f07280733073a074d075e0766077407790772077107;
    inBuf[1867] = 256'h69075a075a075b07580769077d0789079e07ad07b007b707b207a10799078d07;
    inBuf[1868] = 256'h7b077a077e0781079407a407a907ba07c007b007a40792077507630753074307;
    inBuf[1869] = 256'h4807510754076707770778077c0776076107500739071c070f070607ff060b07;
    inBuf[1870] = 256'h17071e073107380730072e0722070a07ff06f106e006e406ea06ec06fd060807;
    inBuf[1871] = 256'h0a0712070e07fc06f306e006c506bb06b106a606ab06ad06ab06b106a9069506;
    inBuf[1872] = 256'h87067006520641062f061e061f0620061f0629062a06200617060306e305c705;
    inBuf[1873] = 256'ha6058405730567055f0567056d056e056d056005460528050205d704b5049904;
    inBuf[1874] = 256'h860485048c049704ad04be04c104be04ac04890464043a041104f703e703e003;
    inBuf[1875] = 256'heb03fe030c04170416040404e803bf038a0358032a030403f302f002f7020903;
    inBuf[1876] = 256'h1b03250328031b03fa02cd029a0267023b0217020302ff0103020c0217021b02;
    inBuf[1877] = 256'h1302fe01d801a80174013f011001ec00d500ce00d100d900e200e500de00cc00;
    inBuf[1878] = 256'hae0086005c0034001000f4ffe2ffdcffdeffddffddffd9ffccffb5ff96ff6eff;
    inBuf[1879] = 256'h45ff1efff8fedbfec7feb6feabfea1fe90fe7dfe66fe44fe1dfef7fdd1fdadfd;
    inBuf[1880] = 256'h90fd76fd62fd54fd43fd31fd20fd04fde2fcbefc95fc6bfc4afc2bfc11fc00fc;
    inBuf[1881] = 256'hf0fbe3fbd6fbbffba4fb88fb5efb33fb0bfbe1fabffaa9fa94fa87fa86fa7cfa;
    inBuf[1882] = 256'h73fa6cfa53fa33fa15faebf9c2f9a5f986f971f96af95ff95bf95df950f940f9;
    inBuf[1883] = 256'h2ef907f9dbf8b5f883f855f834f811f8f8f7eef7ddf7d0f7c8f7aff795f77df7;
    inBuf[1884] = 256'h52f729f70df7e7f6c7f6b7f69ef68cf687f678f668f65cf63df61ff609f6e1f5;
    inBuf[1885] = 256'hbaf5a0f578f557f545f524f509f5fdf4dff4c4f4bbf4a2f48ff48bf476f467f4;
    inBuf[1886] = 256'h66f451f43df437f41ef407f4fff3e5f3d1f3d0f3bef3b2f3b3f39ff38cf383f3;
    inBuf[1887] = 256'h5ff33bf321f3f2f2cdf2baf29af28cf293f28af28df29ef292f287f285f264f2;
    inBuf[1888] = 256'h46f234f20bf2f0f1edf1dbf1d8f1ecf1eaf1ecf1f6f1dff1c5f1b2f17ff151f1;
    inBuf[1889] = 256'h35f10bf1f4f0f9f0f0f0f9f017f11cf124f135f125f112f106f1ddf0c1f0bdf0;
    inBuf[1890] = 256'ha8f0a5f0bcf0c2f0d5f0f4f0f2f0eff0eef0caf0a8f094f066f047f041f02df0;
    inBuf[1891] = 256'h2ff049f050f061f07af074f06ff06ff04df034f02bf00ef005f015f013f021f0;
    inBuf[1892] = 256'h3ff042f04bf05df04bf038f02ff00ef0f7eff6efe4efe4effbef01f013f033f0;
    inBuf[1893] = 256'h33f036f042f033f02af030f023f025f03bf041f057f07cf085f095f0aef0a6f0;
    inBuf[1894] = 256'ha2f0abf09af096f0a6f0a5f0b4f0d8f0e6f0fbf01bf11ef123f131f122f11cf1;
    inBuf[1895] = 256'h26f11ef128f148f154f16df195f1a4f1b8f1d0f1caf1caf1d1f1c3f1c5f1dbf1;
    inBuf[1896] = 256'he1f1f7f11ff236f256f27df288f293f2a4f29ef29ff2acf2a9f2b3f2d0f2e3f2;
    inBuf[1897] = 256'h03f32ff347f365f389f394f3a0f3b3f3b2f3baf3d1f3dbf3f6f322f43ef464f4;
    inBuf[1898] = 256'h95f4b0f4cff4f4f4fef40df525f529f535f550f55ef579f5a3f5bef5e3f510f6;
    inBuf[1899] = 256'h28f643f664f672f685f69df6a9f6c1f6e3f6f9f61cf74af76cf797f7c6f7e4f7;
    inBuf[1900] = 256'h07f82bf83df855f872f882f89cf8bdf8d6f8fcf826f942f968f994f9b4f9d7f9;
    inBuf[1901] = 256'hfcf916fa38fa5dfa78fa9afac1fae2fa0cfb38fb5cfb85fbaffbd2fbfbfb24fc;
    inBuf[1902] = 256'h45fc6bfc91fcaefccffcf0fc0afd29fd48fd67fd8efdb5fdd8fd04fe32fe5afe;
    inBuf[1903] = 256'h85feaefed2fef6fe13ff2dff4dff6aff88ffb0ffdaff06003a0067009200c200;
    inBuf[1904] = 256'he700060125013d01550171018b01ac01d801030236026e02a202d7020a033003;
    inBuf[1905] = 256'h540374038a03a503c103da0300042d0456048d04c904fb04310563058705ad05;
    inBuf[1906] = 256'hcc05db05f4050f06240649067806a506e206210755078f07c007dd07fd071508;
    inBuf[1907] = 256'h1a082b0840084e0871089f08cb080a0948097709af09d909e909020a120a100a;
    inBuf[1908] = 256'h220a3d0a560a890ac10af10a350b750b9d0bcb0be60be80bf50bfa0bf30b0c0c;
    inBuf[1909] = 256'h2a0c440c7f0cbc0cec0c2d0d5d0d720d920da30d9c0dab0db70dbd0de60d130e;
    inBuf[1910] = 256'h3a0e800ec00eea0e1e0f410f480f580f590f4b0f5a0f690f720f9e0fce0ff30f;
    inBuf[1911] = 256'h2f105f107a10a310b610ae10bb10c010b610cd10e510f7102d1160118311be11;
    inBuf[1912] = 256'he811f31110121b120a1212121212031218122e123c126c129612ac12db12fa12;
    inBuf[1913] = 256'hfb120c130b13f412fb12fa12ee120c1328133c1373139e13b113d813ea13df13;
    inBuf[1914] = 256'he613d813b713b513ae13a113bf13db13eb131b143c1440145714551438142f14;
    inBuf[1915] = 256'h1714f413f913fc13f9131f14411452147b148f1485148c147a144b143b142414;
    inBuf[1916] = 256'h02140a141414141437144e144e1464146214421437141b14ee13e513d713c013;
    inBuf[1917] = 256'hd213de13dd13fa130414f413f913e813c013b4139a137513781371135f137013;
    inBuf[1918] = 256'h7313611369135e133c1334131b13f212e812d412b412b612ab12931299128f12;
    inBuf[1919] = 256'h6e12671252122c1222120d12ec11e911d911bb11ba11a81184117b1165113d11;
    inBuf[1920] = 256'h32111c11f810f010dd10ba10b3109f1079106c1052102a101d100310e00fdd0f;
    inBuf[1921] = 256'hcc0fad0faa0f970f720f650f470f1d0f0d0fef0eca0ec30eb00e930e920e830e;
    inBuf[1922] = 256'h620e540e330e010ee40dba0d850d6d0d500d320d310d290d170d180d060de10c;
    inBuf[1923] = 256'hc70c9a0c600c380c080cd80bc80bb70ba60bb00baf0ba10b9b0b7c0b480b1a0b;
    inBuf[1924] = 256'hd50a870a540a230af609ec09e809e609f809f809e409d309a80964092609dd08;
    inBuf[1925] = 256'h920862083c0823082b0835083b084b0843082208f807b4075d071007c0067b06;
    inBuf[1926] = 256'h56063b0630063e064b06500653063c060d06d40587053105e804a40472045d04;
    inBuf[1927] = 256'h5504580467046f04680456042b04ee03a90356030303c1028902620255025302;
    inBuf[1928] = 256'h570261026202520236020502c3017b012f01e800b00085006900610063006900;
    inBuf[1929] = 256'h6d00660050002d00f6ffb0ff63ff16ffd4fe9efe76fe65fe64fe68fe70fe74fe;
    inBuf[1930] = 256'h68fe4cfe1cfedafd90fd40fdf0fcb0fc80fc63fc5dfc62fc6dfc7afc77fc63fc;
    inBuf[1931] = 256'h3efc01fcb4fb65fb14fbcffaa0fa7efa73fa7efa87fa91fa99fa88fa62fa2efa;
    inBuf[1932] = 256'he2f98ff943f9f9f8c2f8a5f894f896f8a7f8adf8adf8a8f883f84ff818f8cff7;
    inBuf[1933] = 256'h88f751f71df7fcf6f4f6ecf6eef6faf6f0f6dcf6c4f691f654f61ef6daf59df5;
    inBuf[1934] = 256'h79f553f53af536f527f51bf516f5f9f4d9f4bff48bf459f437f405f4def3cdf3;
    inBuf[1935] = 256'haff39af394f377f35df34cf31ef3f1f2d3f29ef273f25af22ff20ff204f2e1f1;
    inBuf[1936] = 256'hc4f1b6f18ff16bf156f128f1fff0eaf0c1f0a6f0a1f086f073f071f053f036f0;
    inBuf[1937] = 256'h21f0eeefc1efa4ef6def41ef2fef0beff5eef7eee1eed4eed6eeb5ee95ee80ee;
    inBuf[1938] = 256'h49ee17eefaedc6eda7eda8ed95ed91eda8eda0ed9ceda2ed7eed5aed40ed02ed;
    inBuf[1939] = 256'hcfecb6ec88ec72ec7eec74ec7bec9aec92ec8aec8dec63ec3aec22eceaebc3eb;
    inBuf[1940] = 256'hbbeb9feb9cebb6ebb3ebbcebd6ebc9ebbbebb7eb8ceb69eb5aeb31eb1eeb27eb;
    inBuf[1941] = 256'h19eb1deb39eb34eb37eb47eb2feb1eeb1feb00ebf2eafdeaeaeae9ea00ebf4ea;
    inBuf[1942] = 256'hf0ea00ebebeaddeae3eac7eabceacdeac4eaceeaf2eaf5ea02eb1eeb0feb05eb;
    inBuf[1943] = 256'h0aebe9ead6eae0ead4eae1ea0aeb17eb38eb69eb6feb77eb86eb64eb47eb3beb;
    inBuf[1944] = 256'h10ebfdea0feb12eb33eb75eb9debd2eb0eec19ec22ec2eec0aeceeebe7ebc9eb;
    inBuf[1945] = 256'hc6ebe9ebffeb30ec7beca4ecd2ec02ed00edf7ecefecbeec9aec94ec7eec87ec;
    inBuf[1946] = 256'hb7ecd9ec12ed64ed93edc0edf0edf3edf1edf5edd7edcbedd8edd3edeaed20ee;
    inBuf[1947] = 256'h41ee73eeb2eecbeee4eeffeef3eeefeef5eedeeedbeef1eef5ee10ef41ef5aef;
    inBuf[1948] = 256'h84efbdefd6eff8ef25f033f04bf070f07bf093f0b8f0c2f0d6f0f6f0fdf011f1;
    inBuf[1949] = 256'h31f13af154f182f19bf1bef1eaf1fdf118f237f23cf249f261f265f27cf2a8f2;
    inBuf[1950] = 256'hcaf201f34af380f3bff302f424f442f45df457f457f462f461f474f49df4bff4;
    inBuf[1951] = 256'hf7f43df570f5aaf5e3f5fcf513f62af62bf637f64ff661f68cf6caf602f74af7;
    inBuf[1952] = 256'h98f7cff704f834f849f85cf86ff876f88af8a6f8c2f8f1f829f958f990f9c7f9;
    inBuf[1953] = 256'hedf913fa33fa47fa62fa81faa0fad3fa0dfb43fb86fbc4fbf2fb1ffc42fc53fc;
    inBuf[1954] = 256'h64fc74fc85fca6fcd1fc02fd44fd8dfdcffd10fe41fe5efe6ffe71fe69fe69fe;
    inBuf[1955] = 256'h75fe91fec8fe14ff6fffd7ff37008900c700e300e300d200ae00880077007d00;
    inBuf[1956] = 256'ha600f4005c01d8015702c0020f033b0338031503e102a4027c0277029602e802;
    inBuf[1957] = 256'h6503f4038f041c057e05b705b90583053605dc04850459045f0494040805a405;
    inBuf[1958] = 256'h4706ea066c07b707d307b40761070707af0668065f068f06ed0685073308d708;
    inBuf[1959] = 256'h6f09d109ed09d9098f091a09ae0855081c0829087008e0088409310ac40a410b;
    inBuf[1960] = 256'h8b0b8f0b6c0b210bbb0a6b0a370a250a5a0abe0a3b0bda0b700cdb0c2d0d470d;
    inBuf[1961] = 256'h230de90c920c2c0cef0bd10bd20b180c810cf50c840dff0d4e0e8a0e950e6c0e;
    inBuf[1962] = 256'h420e080ec90db90dc30de00d340e960eef0e570fa10fc20fd90fc80f920f6d0f;
    inBuf[1963] = 256'h460f200f2a0f480f6f0fc00f11104d109510c010c610d110c710a810a410a110;
    inBuf[1964] = 256'h9b10bf10e81006113f116a117811921196117e117a116f115b116d1181118e11;
    inBuf[1965] = 256'hbf11e411f2111712281219121d121412f91100120412ff11231240124c127312;
    inBuf[1966] = 256'h89127f12831274124d1240122c121212221234123f1270129712a912d012df12;
    inBuf[1967] = 256'hcf12cd12b512871278126112431250125c1260128912a512a912c012bf129f12;
    inBuf[1968] = 256'h9512771247123a122b1218122f12471258128d12b312bf12de12e312c312b412;
    inBuf[1969] = 256'h92125a12421224120012081210120f1231124512421257125412321225120812;
    inBuf[1970] = 256'hd811cc11be11ac11c611e011f11120123f1246125c1254122d121612ea11aa11;
    inBuf[1971] = 256'h8b1167113e113e1140113f115e1170116c117c11751150113f111d11ec10de10;
    inBuf[1972] = 256'hcd10b910cd10e410f2101a1136113a11461134110211dc10a11055102910fd0f;
    inBuf[1973] = 256'hd00fcf0fd30fd40ff40f0710061011100110d60fbb0f8b0f4c0f2f0f150fff0e;
    inBuf[1974] = 256'h130f290f390f630f790f730f730f520f0e0fd40e880e320efd0dcc0da40dab0d;
    inBuf[1975] = 256'hb70dc10de70dfe0dfa0df70dd60d970d600d1b0dcf0ca50c860c710c870ca20c;
    inBuf[1976] = 256'hb80cdd0cee0cde0cc60c8d0c330cdd0b7e0b1f0be50abd0aa70abc0ada0af50a;
    inBuf[1977] = 256'h1a0b230b0c0be90aa40a460af1099809480921090f0912093a0960097c099909;
    inBuf[1978] = 256'h930964092409c6085708f6079b0754073b073707470772079607a907b3079907;
    inBuf[1979] = 256'h5e071407b3064c06fa05b6058b0585059005a905d005e605e605d605a7056005;
    inBuf[1980] = 256'h1105b90463042404f603dd03df03eb03fc030e041104ff03e003aa0363031b03;
    inBuf[1981] = 256'hd202910261023e02290221021e021b0217020502e901c30192015b012501f100;
    inBuf[1982] = 256'hc2009b007e006b005c004c003d0028000a00e8ffbdff8cff5aff23ffedfebffe;
    inBuf[1983] = 256'h91fe65fe45fe25fe07fef0fdd3fdb3fd96fd72fd4afd27fdfefcd5fcb4fc90fc;
    inBuf[1984] = 256'h6bfc4cfc2afc07fce9fbc1fb98fb72fb42fb11fbe6fab3fa83fa5cfa30fa08fa;
    inBuf[1985] = 256'he7f9bef995f976f94df924f903f9dbf8b7f89df87bf85cf846f825f804f8ecf7;
    inBuf[1986] = 256'hc6f79af773f73ff70cf7e3f6aef67ff65ef635f614f602f6e2f5c3f5aff58cf5;
    inBuf[1987] = 256'h67f54bf51cf5f0f4d1f4a4f47ef46cf450f43cf43af428f418f412f4f1f3ccf3;
    inBuf[1988] = 256'haef374f33bf311f3d7f2a7f290f271f263f26cf265f265f270f25bf241f22cf2;
    inBuf[1989] = 256'hf4f1bbf195f15df134f129f118f118f131f136f140f151f13cf11df101f1c2f0;
    inBuf[1990] = 256'h80f051f016f0f0efecefe4eff2ef1cf030f047f062f054f03df027f0edefb5ef;
    inBuf[1991] = 256'h8fef58ef39ef3def38ef4aef75ef85ef9aefb4efa1ef88ef73ef38ef06efebee;
    inBuf[1992] = 256'hbeeeaaeebaeebeeedaee0def23ef3fef5fef51ef40ef31effbeecceeb3ee88ee;
    inBuf[1993] = 256'h75ee80ee7dee92eebbeec7eedaeef4eee4eed4eecdeea3ee85ee7cee61ee5eee;
    inBuf[1994] = 256'h76ee7cee95eec1eecfeee1eef8eee8eeddeedceebbeea6eea4ee8dee87ee98ee;
    inBuf[1995] = 256'h93ee9ceeb5eeb3eebaeed0eec8eecbeedeeed6eedceef5eef6ee00ef18ef15ef;
    inBuf[1996] = 256'h1aef2def27ef2def44ef46ef56ef76ef7fef91efabefa8efabefb6efa4ef9bef;
    inBuf[1997] = 256'ha1ef95ef9defbcefcfeff5ef2bf04bf073f0a0f0a8f0b1f0bdf0acf0a3f0abf0;
    inBuf[1998] = 256'ha1f0adf0d2f0ebf015f152f176f19ff1cbf1d1f1d4f1d9f1bff1b0f1b4f1a7f1;
    inBuf[1999] = 256'hb2f1dcf1fdf132f27af2acf2e1f218f32af338f344f32ef31ef31ff311f31af3;
    inBuf[2000] = 256'h41f362f398f3e2f317f44ef484f495f49ef4a4f489f473f46cf45af462f487f4;
    inBuf[2001] = 256'haaf4e4f431f56cf5abf5e6f5fcf509f610f6f9f5eaf5e6f5daf5e5f50cf632f6;
    inBuf[2002] = 256'h6df6b6f6f0f62bf761f775f782f786f771f762f75cf751f75df77ff7a3f7dbf7;
    inBuf[2003] = 256'h1ef854f88ff8c4f8dcf8f2f801f9f8f8f5f8f8f8f5f807f92bf94bf97ff9bdf9;
    inBuf[2004] = 256'hedf923fa53fa6afa7dfa8afa84fa83fa88fa85fa94fab1facefafbfa30fb5bfb;
    inBuf[2005] = 256'h8bfbb6fbd1fbebfbfefb04fc11fc22fc31fc4cfc6ffc90fcb9fce4fc08fd2cfd;
    inBuf[2006] = 256'h4afd5efd74fd86fd95fda8fdbffdd7fdf7fd17fe35fe56fe72fe89fea2feb8fe;
    inBuf[2007] = 256'hccfee7fe05ff28ff50ff78ffa0ffcaffecff07001f002f003a00470055006800;
    inBuf[2008] = 256'h8600aa00d6000801370165019001ab01bd01c901cd01d101d801e201f9011e02;
    inBuf[2009] = 256'h48027c02b802ee022003490362037103760370036d036f0373038703ab03d603;
    inBuf[2010] = 256'h0c0447047e04b104d904ef04fd04fc04f004e704e104de04ee040c0533056905;
    inBuf[2011] = 256'ha205d7050b06300642064d064a063b06310626062206330650067406a906e206;
    inBuf[2012] = 256'h13074407660774077c0775075f07530749073f074d0765078007af07e1070708;
    inBuf[2013] = 256'h310850085b08660865085608520850084c085d0878089208bc08e70806092c09;
    inBuf[2014] = 256'h480951095c0960095409530952094b095809690976099609b709cc09ec09060a;
    inBuf[2015] = 256'h100a230a300a2f0a3b0a460a490a5c0a6f0a7a0a960aaf0abc0ad50ae90aef0a;
    inBuf[2016] = 256'h010b0e0b0f0b1e0b2c0b2f0b410b4f0b500b610b6d0b6e0b7f0b8e0b940bb00b;
    inBuf[2017] = 256'hca0bda0bfc0b190c250c3f0c4c0c470c4f0c4d0c3d0c440c4c0c4e0c6b0c890c;
    inBuf[2018] = 256'h9d0cc60ce60cef0c030d070df40cf10ce70cd00cd90ce70cf00c190d450d650d;
    inBuf[2019] = 256'h980dbb0dc30dd40dd30db70dac0d9b0d810d870d920d9a0dc20dea0d030e2d0e;
    inBuf[2020] = 256'h4a0e4e0e5c0e590e410e3d0e330e200e2b0e390e400e640e850e960ebb0ed20e;
    inBuf[2021] = 256'hd20ee00ee10ecf0ed00ec60eb10eb80ebb0eb40ec90edb0ee00efd0e110f150f;
    inBuf[2022] = 256'h2d0f370f2e0f3a0f390f270f2c0f270f160f1f0f220f1c0f310f3d0f3d0f550f;
    inBuf[2023] = 256'h600f570f630f5f0f480f460f3a0f1f0f200f1a0f0d0f200f2d0f2f0f4d0f620f;
    inBuf[2024] = 256'h640f780f7b0f690f670f550f320f270f150ffa0eff0e010ffc0e170f2b0f300f;
    inBuf[2025] = 256'h480f500f410f400f2c0f050ff30edb0ebb0ebc0ebe0ebf0edf0efa0e070f260f;
    inBuf[2026] = 256'h320f250f200f050fd50eb70e910e680e600e5b0e590e780e930ea40ec50ed20e;
    inBuf[2027] = 256'hc70ec20ea60e780e5b0e350e0c0e040eff0dfc0d190e300e3b0e560e5b0e490e;
    inBuf[2028] = 256'h3c0e190ee40dc10d950d660d570d4c0d410d550d650d6a0d7e0d820d710d680d;
    inBuf[2029] = 256'h4c0d1d0d000dda0cac0c9b0c890c730c780c790c6f0c750c6f0c580c4e0c340c;
    inBuf[2030] = 256'h0b0cf20bd10ba50b900b790b5c0b540b480b350b350b2d0b180b110bff0ae00a;
    inBuf[2031] = 256'hce0aaf0a820a640a3f0a110af609d609b409a709970983098109760961095709;
    inBuf[2032] = 256'h40091c09ff08d508a4088108590831081e080808f307ef07e107ce07c207a407;
    inBuf[2033] = 256'h7a0757072407eb06bd0689065a063e0621060a060506fb05ee05ea05d705b905;
    inBuf[2034] = 256'h9e0573053f051105d804a10478044c04290416040104ef03e703d403bb03a103;
    inBuf[2035] = 256'h760341030b03ca028c0257022402fe01eb01dd01db01e001de01d801c801a301;
    inBuf[2036] = 256'h71013101e100930049000200ceffabff95ff90ff91ff8eff8cff7aff53ff22ff;
    inBuf[2037] = 256'hdffe8efe41fef5fdb1fd86fd68fd59fd60fd67fd6bfd70fd5efd37fd06fdbcfc;
    inBuf[2038] = 256'h65fc12fcbafb6cfb38fb0dfbf5faf6faf5faf6fafcfaecfacbfaa2fa5ffa10fa;
    inBuf[2039] = 256'hc7f975f92bf9fbf8d1f8b9f8baf8b7f8b9f8c0f8aef88df866f820f8cff782f7;
    inBuf[2040] = 256'h28f7daf6a5f673f656f654f64ef651f65cf64cf634f618f6ddf59bf55ef511f5;
    inBuf[2041] = 256'hd0f4a7f479f460f45ef450f449f44cf431f411f4f1f3b3f376f343f3fef2c8f2;
    inBuf[2042] = 256'haaf280f268f267f253f248f247f22af20ff2fbf1ccf1a1f183f150f129f114f1;
    inBuf[2043] = 256'heaf0c9f0bbf095f076f067f03ff01ff010f0e9efccefc2ef9eef81ef75ef4def;
    inBuf[2044] = 256'h29ef15efe7eec2eeb2ee8cee74ee73ee5dee51ee58ee41ee2cee23eef7edcded;
    inBuf[2045] = 256'hb2ed7bed50ed3eed19ed09ed15ed0ded10ed27ed1eed16ed17edf1ecccecb7ec;
    inBuf[2046] = 256'h83ec5eec53ec34ec2cec41ec3eec48ec65ec5cec55ec57ec2fec0becf7ebc2eb;
    inBuf[2047] = 256'h9deb96eb79eb72eb8aeb86eb93ebb3ebacebaaebb4eb91eb74eb68eb38eb15eb;
    inBuf[2048] = 256'h0eebeeeae3eaf4eae7eaeaea07ebfeeaffea12ebfceaedeaf1eaceeab7eab7ea;
    inBuf[2049] = 256'h95ea87ea94ea84ea88eaa8eaa8eab6ead8ead4ead7eae6eacbeab8eab6ea8fea;
    inBuf[2050] = 256'h7aea80ea6eea74ea9aeaa7eac7eafbea0beb20eb3deb2deb20eb1febfaeae6ea;
    inBuf[2051] = 256'hedeadfeaecea1beb33eb60eb9febb7ebd4ebf5ebe7ebdbebdaebb5eba3ebaceb;
    inBuf[2052] = 256'ha2ebb8ebedeb0cec41ec88eca8ecccecf3ececece8ecedeccfecc2eccfecc9ec;
    inBuf[2053] = 256'hdfec12ed2fed60eda0edbceddcedffedf8edf4edf9ede0edd9edeaedeaed06ee;
    inBuf[2054] = 256'h3dee61ee96eed9eefcee21ef48ef49ef4def59ef49ef48ef5eef65ef83efb9ef;
    inBuf[2055] = 256'hddef11f052f076f09df0c9f0d6f0eaf008f110f127f153f172f1a3f1e4f113f2;
    inBuf[2056] = 256'h4df28ef2b4f2e0f210f327f347f371f38bf3b3f3e7f30ef442f47ef4a8f4daf4;
    inBuf[2057] = 256'h11f533f55ef58ff5b2f5dff516f640f674f6aff6dbf60bf73ef75ef784f7aff7;
    inBuf[2058] = 256'hcaf7eff71cf841f870f8a5f8cef8fdf82df94bf96df98ff9a3f9bdf9dff9fbf9;
    inBuf[2059] = 256'h24fa58fa86fabffafcfa2dfb5ffb8dfbaafbc7fbe2fbf4fb0dfc2bfc4afc76fc;
    inBuf[2060] = 256'haafcddfc17fd50fd7ffdadfdd5fdf0fd0bfe25fe3dfe5ffe89feb6fef1fe31ff;
    inBuf[2061] = 256'h71ffb4fff0ff2300510073008e00a900c100dd0003012f016401a001dd011a02;
    inBuf[2062] = 256'h54028302ac02d002e80200031d03390360039003c203fc0339046c049d04c704;
    inBuf[2063] = 256'he104f8040c0519052d05490567059405c705f4052806560674069006a306a706;
    inBuf[2064] = 256'hb006bd06c606e206080730076807a107cf070008280839084c08580857086608;
    inBuf[2065] = 256'h7b088e08ba08ef0820096209a109ce09010a2a0a3c0a580a700a7d0aa10acb0a;
    inBuf[2066] = 256'hf00a2f0b720bab0bf60b390c670ca10cd00cea0c130d380d4f0d7e0dad0dd10d;
    inBuf[2067] = 256'h0f0e4c0e790ebb0ef70e1e0f580f8a0fa40fd20ff80f0b103210521060108610;
    inBuf[2068] = 256'ha710b510dc10fd100c1132114f115711741187118211921199118a1194119911;
    inBuf[2069] = 256'h8d119e11ab11a811c011d111cd11e011e711d411d811cf11b211b011a8119011;
    inBuf[2070] = 256'h9911a2119b11b511c811c511dc11e811da11e211dd11c311c911ca11bc11d511;
    inBuf[2071] = 256'hed11f711241249125912811298129312a612a81293129f12a6129f12c212e412;
    inBuf[2072] = 256'hf7122e135a136d139a13b213ab13bd13be13a813b613bf13bc13e21304141514;
    inBuf[2073] = 256'h48146a146e148b1490147414731461143b143a14341423143c144d144d146c14;
    inBuf[2074] = 256'h79146a147214621438142b141214e813e713e213d213eb13fa13f5130c140f14;
    inBuf[2075] = 256'hf613f813e513bb13b413a5138c13a013b013b413de13fd13041424142d141b14;
    inBuf[2076] = 256'h24141e14061417142914331469149d14c2140615361548156e15781565157015;
    inBuf[2077] = 256'h6d155e157e15a115bd15051645166f16b016d416d016db16c9169b168b167516;
    inBuf[2078] = 256'h561668167e168a16bc16df16e316f416e216a71678163016d115951557151615;
    inBuf[2079] = 256'h0415f414da14df14cf14a0147d143914d31380131a13a61257120812ba119711;
    inBuf[2080] = 256'h711140112c110511c51096104e10f00fac0f5b0f010fcd0e980e610e500e390e;
    inBuf[2081] = 256'h180e150e020edf0dd20db40d850d6f0d4c0d200d130dfe0ce30ce90ce90ce10c;
    inBuf[2082] = 256'hf60c010d010d160d1b0d120d1b0d130dfd0cfb0cef0cdb0ce20ce30ce00cf70c;
    inBuf[2083] = 256'h050d0a0d220d270d1b0d1b0d080de30cca0ca40c780c610c420c220c1a0c050c;
    inBuf[2084] = 256'hea0be00bc70b9f0b820b500b110be10aa30a600a310af809bf099e0973094409;
    inBuf[2085] = 256'h2709fe08ce08a908750838080708ca07880757071c07e206be0695066c065806;
    inBuf[2086] = 256'h410629061d060706ee05de05c205a0058a056b054c053c052b05200525052805;
    inBuf[2087] = 256'h30053f0548054d0553054b053d0530051705fe04eb04d604c704c004ba04bc04;
    inBuf[2088] = 256'hc004bb04b604ad049804790450041b04e403aa036b033203fb02c50297026702;
    inBuf[2089] = 256'h33020202c7017c012f01d5006c00040094ff1fffb4fe4cfee7fd91fd3dfde8fc;
    inBuf[2090] = 256'h9ffc4efcf5fb9efb3cfbcefa64faf3f982f91cf9b6f858f80ff8c8f789f75bf7;
    inBuf[2091] = 256'h29f7f4f6c8f691f654f61df6d9f597f565f52ef502f5eef4dbf4d6f4e6f4f0f4;
    inBuf[2092] = 256'hfbf411f517f518f51cf50cf5fcf4f7f4e6f4e1f4f1f4fbf413f53ff55ff583f5;
    inBuf[2093] = 256'haff5c2f5cef5dbf5cef5bef5b5f59af589f58af57df57cf58cf588f588f591f5;
    inBuf[2094] = 256'h7df564f551f520f5ecf4c4f485f44bf423f4e8f3b2f38ff357f323f300f3c7f2;
    inBuf[2095] = 256'h8ef262f21ff2def1abf160f116f1dbf089f03df006f0bdef7def58ef24effcee;
    inBuf[2096] = 256'hebeec6eea7ee97ee6cee41ee23eeededbceda3ed7ced69ed73ed71ed82edabed;
    inBuf[2097] = 256'hbdedd3edf3edefedeaedeeedd1edbeedc1edb1edbbede4edfced29ee6bee8dee;
    inBuf[2098] = 256'hb3eee1eee1eedeeee4eec2eea8eea6ee88ee80ee98ee94eea0eec2eebaeeb2ee;
    inBuf[2099] = 256'hb2ee7fee46ee18eebded68ed2cedd2ec8dec69ec27ecf7ebe1eba4eb6beb40eb;
    inBuf[2100] = 256'he4ea86ea38eac0e953e901e994e83de80be8bde785e76ae72ce7f9e6d8e689e6;
    inBuf[2101] = 256'h41e60de6b5e56ce541e5fee4d6e4d2e4b7e4b6e4d4e4d3e4e2e407e507e515e5;
    inBuf[2102] = 256'h37e538e54be578e589e5b1e5f4e51ae656e6a9e6dbe61fe779e7ade7f2e74de8;
    inBuf[2103] = 256'h81e8c6e81de94ce989e9d9e901ea38ea83eaaaeae5ea37eb66eba6ebf7eb1dec;
    inBuf[2104] = 256'h50ec8eec97eca2ecb8eca0ec94ec9bec7fec79ec90ec87ec90ecafeca7eca3ec;
    inBuf[2105] = 256'ha7ec7aec4dec27ecd7eb94eb69eb23ebf6eae9eac7eabaeac6eab2eaa4ea9cea;
    inBuf[2106] = 256'h69ea39ea12eacbe993e973e942e92ee93de93fe95ae98ee9a7e9cce9fae901ea;
    inBuf[2107] = 256'h0bea20ea18ea20ea3fea4dea79eac6ea04eb5bebc8eb1aec77ecdbec18ed5bed;
    inBuf[2108] = 256'ha7edcfed06ee53ee8aeed9ee44ef98ef03f07ef0d8f03af19ff1d9f117f25bf2;
    inBuf[2109] = 256'h79f2a0f2d7f2f2f220f35ef382f3b5f3f2f310f435f45ff467f477f48af482f4;
    inBuf[2110] = 256'h88f495f487f489f495f48af489f490f47ff478f479f468f463f463f451f44df4;
    inBuf[2111] = 256'h4ef43bf433f430f41df416f41af418f426f444f461f48ef4c8f4fbf436f573f5;
    inBuf[2112] = 256'ha0f5d0f502f629f659f692f6ccf61bf778f7d7f748f8bff82bf99af903fa57fa;
    inBuf[2113] = 256'ha9faf8fa37fb80fbd5fb2bfc94fc09fd7efd01fe85fef8fe66ffc5ff0a004a00;
    inBuf[2114] = 256'h8100a600d100030133017001b401f40139027702a102c202d202cd02c102aa02;
    inBuf[2115] = 256'h8c02770265025502540257025a025f025a024a0231020a02d901a5016b013201;
    inBuf[2116] = 256'h0101d500b000940079006500510036001d000100dfffc3ffa8ff8dff80ff79ff;
    inBuf[2117] = 256'h73ff7aff87ff94ffaaffc0ffd3ffefff0f002b0054008400b200ed002b016201;
    inBuf[2118] = 256'ha401e90128027302c00208035e03bb0312047704e2044005a30507065a06b106;
    inBuf[2119] = 256'h06074f07a307f80742089c08ff085509b309130a5f0aae0af70a290b600b960b;
    inBuf[2120] = 256'hbc0beb0b1b0c410c790cb20cdd0c130d430d5e0d820d9d0da10db10dbb0db50d;
    inBuf[2121] = 256'hc30dcf0dcd0de40dfa0d010e1d0e330e380e530e640e640e7e0e900e950eba0e;
    inBuf[2122] = 256'hd90eea0e1e0f4d0f690fa30fd40ff10f2a1058107110a810d710f61039117411;
    inBuf[2123] = 256'h9d11ec1134126a12be12051335138013bf13ea1332146e149814e31421154915;
    inBuf[2124] = 256'h8f15c615e1150f16281625163516341622162a16241612161e161b1604160116;
    inBuf[2125] = 256'he815b21587154415eb14a5144e14f013af1365131613e2129d124a1201129b11;
    inBuf[2126] = 256'h1f11ac101d10850f040f770eef0d8b0d200db70c6b0c100cab0b560be30a640a;
    inBuf[2127] = 256'hfc097e090109a8084b08f707ce079f076f075f073d070d07f306c50688066906;
    inBuf[2128] = 256'h4206180618061906190642066a068806c206f306150750078207a707e9072908;
    inBuf[2129] = 256'h5e08b5080c095209b1090c0a530ab20a0e0b570bb60b150c660ccf0c380d8c0d;
    inBuf[2130] = 256'hf40d550e9a0eee0e3e0f760fbf0f0a1048109c10ef1035118f11df1112125412;
    inBuf[2131] = 256'h86129712b612cd12cf12ee121113291362139a13c413081439144a146e147a14;
    inBuf[2132] = 256'h65146a1467145314681480148f14cc14051528156a1596159f15bf15c515a915;
    inBuf[2133] = 256'hb015ae159d15be15e015f91545168a16bb160d1745175a178a179d179217a717;
    inBuf[2134] = 256'had17a317c517de17eb171e1841184e1875187f186a18681848180f18ed17ba17;
    inBuf[2135] = 256'h7b1758172c17f916e016b81683165e161e16ca157c1513159b142d14a2130d13;
    inBuf[2136] = 256'h8b12f9116611e4105210c10f3e0fa40e060e730dc50c0f0c640ba40ae5093309;
    inBuf[2137] = 256'h7208b90715076506c0052d058b04f1036703cb023102a40105016800dbff44ff;
    inBuf[2138] = 256'hb7fe3cfebafd46fdedfc91fc3ffc04fcc6fb8ffb69fb3bfb0dfbeefacbfaabfa;
    inBuf[2139] = 256'h9bfa8ffa8bfaa0fac0faeafa29fb71fbb8fb06fc4ffc8bfccafc06fd35fd6bfd;
    inBuf[2140] = 256'hacfdeffd4bfec0fe39ffc5ff6300f2007e010a027c02df023c038503d0032804;
    inBuf[2141] = 256'h7d04e5046605e805730606078607fd076708af08ed08240947097209a809e109;
    inBuf[2142] = 256'h310a8f0aec0a560bba0b040c4c0c810c970cab0cb40cb00cc10cd60ceb0c1c0d;
    inBuf[2143] = 256'h520d810dc30dfb0d1d0e470e5d0e5c0e6b0e700e650e720e7e0e840ea30ec00e;
    inBuf[2144] = 256'hd20ef80e130f1f0f390f470f440f4f0f4c0f3c0f370f240f080ffd0ee70ecb0e;
    inBuf[2145] = 256'hc00ead0e960e8f0e7d0e640e4e0e250ef20dbb0d6f0d1f0dce0c6c0c140cc40b;
    inBuf[2146] = 256'h670b150bc90a6c0a110aad092d09ac081c086e07c6061c066105b90417046e03;
    inBuf[2147] = 256'hdf025302b80129019200e0ff30ff71fe9afdccfcf6fb18fb50fa86f9bdf80ff8;
    inBuf[2148] = 256'h60f7abf60cf662f5aaf4fff346f381f2cdf115f15ef0bfef22ef90ee1aeea8ed;
    inBuf[2149] = 256'h3aeddfec81ec25ecd6eb7ceb29ebe5ea99ea5aea31ea09eaf3e9f1e9eee9fae9;
    inBuf[2150] = 256'h17ea2dea4fea7bea9fead3ea11eb46eb91ebeeeb45ecb0ec29ed98ed19eea4ee;
    inBuf[2151] = 256'h1defa6ef36f0b7f047f1daf15bf2eef288f30ff4a3f43af5bbf546f6d3f64af7;
    inBuf[2152] = 256'hcef755f8c8f848f9cbf93cfab9fa35fb99fb05fc6afcb1fcfefc48fd7afdb3fd;
    inBuf[2153] = 256'heefd1dfe57fe93febffef3fe23ff3fff5bff71ff72ff73ff72ff69ff6aff72ff;
    inBuf[2154] = 256'h77ff86ff98ffa3ffb1ffbaffafff9cff85ff63ff43ff27ff0cff00ff03ff08ff;
    inBuf[2155] = 256'h1aff32ff3dff41ff41ff2eff0effedfec0fe92fe72fe57fe48fe4efe50fe53fe;
    inBuf[2156] = 256'h5cfe53fe39fe1afedffd98fd57fd04fdb6fc80fc3ffc05fce7fbb6fb78fb47fb;
    inBuf[2157] = 256'hf9fa96fa38fabbf934f9c2f839f8b1f749f7d0f654f6f2f572f5e4f467f4c2f3;
    inBuf[2158] = 256'h10f373f2b5f1f1f04cf08fefd5ee3fee8fede1ec51ec9eebe6ea4cea95e9dde8;
    inBuf[2159] = 256'h47e898e7f0e669e6cce538e5c2e431e4a8e33ae3b0e22fe2cbe152e1ebe0a6e0;
    inBuf[2160] = 256'h52e014e0f5dfc4dfa8dfa7df8edf87df9adf97dfa9dfd6dff4df2ce081e0c9e0;
    inBuf[2161] = 256'h2fe1ace112e294e22be3a3e32ce4c6e448e5dee584e613e7c1e783e82ee9f5e9;
    inBuf[2162] = 256'hccea82eb48ec15edb9ed6aee1fefaaef48f0f5f07ff121f2d6f269f30ff4bcf4;
    inBuf[2163] = 256'h39f5bff541f68af6d5f623f743f770f7abf7c2f7eef72bf843f865f88ef888f8;
    inBuf[2164] = 256'h7df871f836f8fbf7cbf77ff73ff716f7dff6b5f69af66cf643f61af6d2f588f5;
    inBuf[2165] = 256'h3ef5e0f489f443f4fbf3caf3b0f394f387f38af381f378f372f35cf345f336f3;
    inBuf[2166] = 256'h21f319f326f339f361f39cf3d4f319f463f498f4d2f40ff534f560f598f5c3f5;
    inBuf[2167] = 256'h00f654f69bf6f0f655f7a2f7eff73ef866f88cf8b4f8b4f8b9f8cef8c5f8c8f8;
    inBuf[2168] = 256'he4f8e4f8eaf801f9f1f8daf8c6f882f836f8f2f785f716f7bbf645f6d7f580f5;
    inBuf[2169] = 256'h11f5a8f44ff4d3f355f3e1f246f2a4f10ff15df0abef10ef68eecded4bedbfec;
    inBuf[2170] = 256'h44ecddeb65ebf4ea8eea14eaa1e93ae9c4e85ee80fe8bfe788e76de755e758e7;
    inBuf[2171] = 256'h72e788e7afe7e3e70ce841e87fe8b5e8fee853e9a8e91deaa4ea2bebd2eb8aec;
    inBuf[2172] = 256'h38edfaedbeee71ef37f0f9f0a7f16bf232f3e5f3b3f48ff559f636f715f8ddf8;
    inBuf[2173] = 256'hb3f981fa2cfbdffb8bfc14fda7fd37fea9fe2affacff10007b00e20024016701;
    inBuf[2174] = 256'ha101b401c601d401c001ad019a016c0142011a01db009d0060000e00b8ff61ff;
    inBuf[2175] = 256'hfcfe94fe29feb3fd3efdcbfc53fce0fb6efbfdfa96fa36fad9f981f930f9e9f8;
    inBuf[2176] = 256'ha8f869f837f80bf8e2f7caf7bbf7b4f7c6f7e9f714f854f8a3f8f5f857f9c2f9;
    inBuf[2177] = 256'h2afa9ffa18fb8dfb13fca6fc36fdd8fd8dfe41ff0300d00096015e022903e503;
    inBuf[2178] = 256'h9b045405ff05a1064907ea0786082709c109500ade0a620bda0b480ca50cf30c;
    inBuf[2179] = 256'h3a0d6e0d920dad0db50dac0d9c0d830d5b0d280def0cb10c6a0c1d0ccc0b6d0b;
    inBuf[2180] = 256'h040b990a1b0a92090c097908dd074f07c0063306bc054505d004700407049803;
    inBuf[2181] = 256'h3b03d1025d0201029f013e010701da00b400ba00c700d5000701350157019401;
    inBuf[2182] = 256'hce01f9013f028d02da024c03ca034804eb0497053606e80699073808e2088a09;
    inBuf[2183] = 256'h230aca0a740b160cc70c7c0d250ed40e7e0f1510a8102b119b1108126412b012;
    inBuf[2184] = 256'hff1246137d13b513e413051420142b1424141614f413c2138e134a13f712a812;
    inBuf[2185] = 256'h4e12e911891119119e102a10a70f1b0f9d0e100e780df30c640cce0b500bc80a;
    inBuf[2186] = 256'h350abe094009ba085508e90773072607da0686065d0635060306ff05fd05ee05;
    inBuf[2187] = 256'h0d062b0637067306b106db0634079307e1075e08dc084509df097e0a030bb20b;
    inBuf[2188] = 256'h640cfc0cba0d790e1f0fe80fb31067113c121013cb13a21473152716f216b217;
    inBuf[2189] = 256'h5118ff18a019211aaf1a321b9c1b141c7c1cce1c351d8e1dcb1d141e491e611e;
    inBuf[2190] = 256'h811e891e721e641e401e031ed51d941d421d071db91c571c101cb41b411be41a;
    inBuf[2191] = 256'h6f1adf196719d9183518b31720177c1602167f15ef148e142014a5135513f212;
    inBuf[2192] = 256'h7b123112d41165112511db1087106c104b10221031103810301056106c106d10;
    inBuf[2193] = 256'h9110a1109f10c410de10f21038117d11bc1127128c12e1125113ac13e9132b14;
    inBuf[2194] = 256'h5414671488149a14a214c714e7140115311558156b1582157c1554152615dd14;
    inBuf[2195] = 256'h7a141b14b1134213e8128a122912d611761105119110fb0f4a0f980ec80de80c;
    inBuf[2196] = 256'h1b0c490b7b0ad2092c098c080f088a07ff068806f8055705cc042b048103fc02;
    inBuf[2197] = 256'h7502f201a4015d011d010d01fe00ee0002010a0107012301340137015d018001;
    inBuf[2198] = 256'h9f01e80137028602000384030404a7044b05e1058f063707c5076308f9087709;
    inBuf[2199] = 256'h080a9a0a1e0bbb0b610cfb0caa0d5d0efa0e9c0f3110a61017117411af11eb11;
    inBuf[2200] = 256'h24124e128712ca120c136013b81303144b147d14921493146c142514d5137213;
    inBuf[2201] = 256'h0713ab124f120112cd11951161113711f110911023108e0fe20e2e0e600d990c;
    inBuf[2202] = 256'heb0b3f0bab0a3d0acd09690913099f081a088e07d7060b06420567049603ea02;
    inBuf[2203] = 256'h4902c70171012501eb00bc0076002200c6ff43ffb2fe24fe8cfd03fd9bfc4afc;
    inBuf[2204] = 256'h1bfc10fc15fc2afc43fc4dfc4afc2cfcf3fbb2fb60fb04fbbafa7bfa4cfa3ffa;
    inBuf[2205] = 256'h40fa4dfa6dfa7ffa86fa8bfa6efa3bfa04fab1f956f90cf9b3f863f82df8edf7;
    inBuf[2206] = 256'hb4f78ef74df705f7c2f65df6e8f575f5e4f451f4cdf335f3a5f22ef2acf139f1;
    inBuf[2207] = 256'hdef074f010f0beef57efefee90ee19eea0ed2ceda6ec28ecc0eb56eb02ebccea;
    inBuf[2208] = 256'h99ea80ea84ea86ea95eaafeabceaceeae3eae6eaf3ea0feb25eb54eb9febf3eb;
    inBuf[2209] = 256'h64eceeec76ed0deeaaee2eefb3ef33f096f0fbf065f1c2f135f2bbf240f3e4f3;
    inBuf[2210] = 256'h99f43df5f1f5a3f62ef7b7f731f87cf8c9f816f945f985f9d8f91dfa7dfaf0fa;
    inBuf[2211] = 256'h49fba8fb05fc33fc52fc64fc44fc1afcedfba2fb62fb3dfb0dfbf4faf7faedfa;
    inBuf[2212] = 256'hecfaf5fadafab0fa80fa24fab9f953f9d2f850f8e8f77bf71ff7dff697f653f6;
    inBuf[2213] = 256'h1cf6c8f56af510f594f40cf48df3fcf273f20af29af13af102f1c2f084f05cf0;
    inBuf[2214] = 256'h21f0deefa4ef4defebee94ee29eec5ed78ed22eddcecb5ec81ec5dec54ec37ec;
    inBuf[2215] = 256'h1fec1becfbebddebd1ebaaeb88eb78eb4feb36eb39eb28eb29eb49eb54eb72eb;
    inBuf[2216] = 256'habebc4ebe4eb14ec1bec23ec38ec25ec18ec1dec06ec05ec22ec2cec4eec87ec;
    inBuf[2217] = 256'ha2ecccecffec02ed0aed16edf5ecddecd6ecb1eca4ecb3ecacecbdece3eceaec;
    inBuf[2218] = 256'hf8ec0bedf5ecddecc2ec86ec59ec3dec13ec05ec13ec1dec46ec82ecaaecdeec;
    inBuf[2219] = 256'h13ed2aed45ed5eed60ed71ed8eeda3edd5ed1cee63eec6ee37ef9bef0ef084f0;
    inBuf[2220] = 256'he7f056f1c5f124f293f20cf37bf302f497f423f5c5f56ef603f7a4f746f8cbf8;
    inBuf[2221] = 256'h55f9ddf948fab8fa28fb84fbedfb5afcb3fc1afd86fddafd38fe95fed4fe13ff;
    inBuf[2222] = 256'h49ff5eff73ff86ff7dff75ff70ff5eff56ff54ff41ff35ff2cff0dffe8fec0fe;
    inBuf[2223] = 256'h80fe36fee7fd89fd2cfdd6fc7bfc2dfcf0fbb3fb7bfb52fb29fbfdfad4faa8fa;
    inBuf[2224] = 256'h7afa4ffa20faf4f9d2f9b4f99bf98ff986f980f981f980f980f985f988f98af9;
    inBuf[2225] = 256'h92f999f9a6f9b9f9ccf9e9f90efa33fa5ffa90fabffaf3fa27fb53fb83fbb0fb;
    inBuf[2226] = 256'hcffbeffb0dfc1afc29fc3bfc42fc4dfc5dfc67fc79fc8efc98fca6fcb6fcb6fc;
    inBuf[2227] = 256'hb3fcaffca0fc8efc82fc71fc64fc5efc5afc5dfc63fc64fc66fc65fc59fc49fc;
    inBuf[2228] = 256'h38fc1ffc07fcf5fbe5fbddfbddfbe2fbeefbfafb07fc19fc28fc33fc44fc53fc;
    inBuf[2229] = 256'h63fc7efc9cfcc0fcf3fc27fd5efd9ffddbfd17fe59fe95fecdfe0bff44ff80ff;
    inBuf[2230] = 256'hc2fffdff40008f00d70025018101d90133029902fa025f03c80329048b04ef04;
    inBuf[2231] = 256'h44059905ef053a068606d80623077407ca071a086e08c208070946098109b009;
    inBuf[2232] = 256'hda09fe09190a390a5a0a760a960ab60ace0ae40af20aed0adc0ac10a990a680a;
    inBuf[2233] = 256'h2e0aee09b20974093409fa08ba0872082c08d8077c072507c0065506fa059b05;
    inBuf[2234] = 256'h3c05f004a0044c040b04c50377033603ec02980259021902d601ae0189016401;
    inBuf[2235] = 256'h5a01510144014c01530155016b0181019701c601f9012d027d02d10223038603;
    inBuf[2236] = 256'he40337049704ef0437058905da0520066d06bc06050752079907d50715085108;
    inBuf[2237] = 256'h7f08ad08d808f80818093109410950095a0955094d093c091b09fa08d4089f08;
    inBuf[2238] = 256'h6b083608f607b90779072e07e40694063b06e40589052a05da048b043a040104;
    inBuf[2239] = 256'hcf039c037c035b03370326031003ef02e202d502bf02c002c602ca02e6020403;
    inBuf[2240] = 256'h1f0353038b03b803f8033a047004b904060549059d05f6054506a10601075807;
    inBuf[2241] = 256'hbb071e087508d3082e097b09cc09170a510a8d0ac30ae90a110b360b500b6f0b;
    inBuf[2242] = 256'h8a0b9d0bb20bbd0bbc0bbc0bb30b9a0b800b5c0b2f0b080bdf0ab20a8c0a620a;
    inBuf[2243] = 256'h300a030ace098c094809fa08a1084b08ed078f074007f206a90672063906fe05;
    inBuf[2244] = 256'hce0592054e051205cc047c043904f803bc03950370034f0341032e0314030603;
    inBuf[2245] = 256'heb02c102a2027b024b022e02170204020b021b022e0258028302a402ce02f102;
    inBuf[2246] = 256'h070325033a0343035a0372038403a803d60302043b047404a804e70423055205;
    inBuf[2247] = 256'h8505b505d705fc052106450670069b06c406f506260753078307ac07cc07e907;
    inBuf[2248] = 256'hf807f807f407e707cf07b907a2078a07780768075607470733071807fc06d106;
    inBuf[2249] = 256'h9b0669063006f305c505960567054f053d05280521051605ff04f204db04b504;
    inBuf[2250] = 256'h99047a0454044304380430043f04530468049104ba04dc040c0539055d058f05;
    inBuf[2251] = 256'hbe05e705230662069e06e5062b076d07b407f10723085b088608a108be08d508;
    inBuf[2252] = 256'he308f308fe08060914091f0924092509200915090109df08b60883083f08f507;
    inBuf[2253] = 256'ha7074f07f4069d064006eb059b054205e80496043904d2036903f3027a020702;
    inBuf[2254] = 256'h8e011901b5005500fdffbdff81ff48ff21fffbfed1feaffe8afe63fe48fe2cfe;
    inBuf[2255] = 256'h14fe11fe14fe1bfe38fe5afe7ffeb3fee8fe17ff4eff83ffb1ffe5ff1c005300;
    inBuf[2256] = 256'h9400d7001c016b01bc0109025902a502e90227035d038803ad03c703d903ee03;
    inBuf[2257] = 256'h00040e041f042f043f0451045e04620461045b044b042f040c04e303b3037d03;
    inBuf[2258] = 256'h48031503e202b20285025a022d02fe01cb01920157011a01dd00a10067003500;
    inBuf[2259] = 256'h0f00edffcdffb9ffabff9aff8aff7bff69ff57ff42ff2eff24ff1dff1bff26ff;
    inBuf[2260] = 256'h37ff4dff6bff8affa7ffc7ffe3fff7ff0a001b002b0042005a0075009a00c500;
    inBuf[2261] = 256'hf5002c0163019901cf0101022d0251026c02830295029e02a602ae02b302b802;
    inBuf[2262] = 256'hbb02be02c402c202ba02b302a4028d02740250022702ff01ce019a016b013601;
    inBuf[2263] = 256'hff00cc008d0048000700bbff64ff0effaffe4afeedfd89fd22fdc7fc6dfc10fc;
    inBuf[2264] = 256'hbbfb61fb03fbadfa54faf4f99bf93ff9e3f897f84bf802f8c8f792f75ff73cf7;
    inBuf[2265] = 256'h1bf7f7f6def6c9f6b3f6a6f69bf690f68cf68cf691f69ff6adf6bff6d8f6f0f6;
    inBuf[2266] = 256'h10f73cf764f793f7cff70cf84df895f8d7f81df966f9a4f9e6f928fa5cfa95fa;
    inBuf[2267] = 256'hd4fa01fb32fb69fb8ffbb7fbe3fb01fc23fc47fc5afc73fc8efc93fc9bfca8fc;
    inBuf[2268] = 256'ha0fc99fc8ffc6cfc49fc28fceefbb7fb8bfb50fb16fbe8fab0fa7ffa54fa1afa;
    inBuf[2269] = 256'he2f9aff96df92bf9eef8a5f85ff81ff8d7f798f762f728f7f9f6d2f6a3f67ff6;
    inBuf[2270] = 256'h67f649f633f627f61bf61af620f622f631f643f64cf661f67df68ff6aaf6cef6;
    inBuf[2271] = 256'he9f60ff73ff769f79bf7d7f709f842f880f8b2f8e7f823f950f97ff9b2f9d6f9;
    inBuf[2272] = 256'hfaf924fa3cfa4ffa68fa73fa7dfa8bfa89fa8cfa98fa95fa94fa99fa8bfa7dfa;
    inBuf[2273] = 256'h75fa5afa39fa1cfaecf9b8f98cf94ef90ef9d7f892f84ef815f8ccf784f746f7;
    inBuf[2274] = 256'hfff6bef68df651f618f6ecf5baf58cf564f52df5f9f4c9f48df455f425f4f2f3;
    inBuf[2275] = 256'hccf3b6f3a0f39df3a9f3b0f3c2f3def3edf3fff312f416f420f42ef432f441f4;
    inBuf[2276] = 256'h5af46df48df4bbf4e4f416f54ff57ff5b9f5f6f528f662f6a1f6d4f612f754f7;
    inBuf[2277] = 256'h88f7c3f7fff729f859f889f8a6f8c6f8e8f8f8f812f932f947f968f990f9a9f9;
    inBuf[2278] = 256'hcff9fff91dfa40fa65fa78fa8bfa9afa94fa94fa95fa82fa76fa72fa67fa67fa;
    inBuf[2279] = 256'h70fa72fa81fa98faa2fab1fabefabbfabafab6faa1fa91fa81fa68fa56fa4cfa;
    inBuf[2280] = 256'h3efa3cfa40fa3dfa43fa4dfa4bfa50fa5dfa64fa73fa89fa9cfab9faddfafcfa;
    inBuf[2281] = 256'h1cfb39fb4bfb5dfb6cfb70fb75fb7afb7dfb8bfba3fbc1fbf0fb29fc62fca7fc;
    inBuf[2282] = 256'heffc2ffd70fdaafdd1fdf7fd18fe2afe39fe47fe4ffe62fe7cfe90feadfed4fe;
    inBuf[2283] = 256'hf6fe1dff4bff6cff87ffa3ffb8ffc2ffc4ffbeffb5ffa6ff90ff7dff6cff56ff;
    inBuf[2284] = 256'h42ff32ff1fff0cfffafee8fed7fec7feb6fea7fe9afe8dfe83fe7bfe71fe64fe;
    inBuf[2285] = 256'h52fe40fe2cfe12fef6fddbfdc1fdaefda3fda1fdb0fdcbfdedfd1bfe50fe84fe;
    inBuf[2286] = 256'hbbfef0fe1cff43ff65ff81ff9dffb5ffccffeeff180045007e00c3000d015d01;
    inBuf[2287] = 256'hb10106025c02ae02f8023f038303c003f503270457048104a504c604e7040105;
    inBuf[2288] = 256'h17052d0543055405680581059a05b805db05fa051b063b065406670671066b06;
    inBuf[2289] = 256'h5b063f061806f005c40593056f0553053c0539053e05420555056b0577058705;
    inBuf[2290] = 256'h8d05810578056805480530051805fd04f604f404f0040405200538055f058805;
    inBuf[2291] = 256'haa05d405fa0516063c065b066e068e06a806b706d106e606f00608071e072a07;
    inBuf[2292] = 256'h43075d0773079b07c607ee0726085f089208cf0805092c09520969096e097209;
    inBuf[2293] = 256'h68094f093c0925090909fc08f308ed08fc080e091d093e09570964097a098709;
    inBuf[2294] = 256'h81097e096f09500939091709e908ca08a60879085f08460827081d0812080208;
    inBuf[2295] = 256'h08080b0805081008120808080c080308e907dd07c807a4079307810769076807;
    inBuf[2296] = 256'h69076a078607a507c007f40727084e088608b608d60802092309330953096909;
    inBuf[2297] = 256'h71098b09a409b809e609150a400a870ad20a120b660bb60bf30b3a0c780ca30c;
    inBuf[2298] = 256'hd20cf00cfb0c100d1c0d190d240d290d230d2f0d3a0d3c0d4d0d5a0d600d760d;
    inBuf[2299] = 256'h820d830d8e0d890d720d650d450d100de10ca40c580c190cd00b800b470b0a0b;
    inBuf[2300] = 256'hc90aa20a7b0a4f0a380a1e0afa09e709cb09a3098b09670935091209e308a808;
    inBuf[2301] = 256'h800851081c080208e807cd07d307da07df0703082808450876089f08b608d808;
    inBuf[2302] = 256'hee08f508070910091109250939094c097709a109c709030a3b0a6b0aa80adb0a;
    inBuf[2303] = 256'h020b320b530b630b770b7b0b6e0b680b560b380b240b080be80ad60ac00aab0a;
    inBuf[2304] = 256'ha70a9d0a8f0a8d0a820a6b0a560a310afd09cc098c094109fb08a6084b08fe07;
    inBuf[2305] = 256'ha7074e070907c0067a064c061c06ef05da05c205a6059b058705680554053305;
    inBuf[2306] = 256'h0305df04b1047e045e043f041f04190419041a0431044c0465048e04b504d404;
    inBuf[2307] = 256'hfd04200539055b0578058e05ab05c105d305ec05000610062906450663068c06;
    inBuf[2308] = 256'hb906e6061a074a0773079b07b807c907d307cd07b907a30782075b0734070807;
    inBuf[2309] = 256'hdd06bb069b067c06630647062d061706f905d405ad057b053c05f504a1044304;
    inBuf[2310] = 256'hdd036c03fd0291022202be0163010d01c500840042000800d0ff8eff4eff0eff;
    inBuf[2311] = 256'hc4fe7bfe32fee0fd95fd4ffd04fdc1fc87fc4bfc13fce7fbbffb9ffb88fb7bfb;
    inBuf[2312] = 256'h77fb79fb83fb95fba8fbbafbcbfbd5fbddfbe1fbdcfbd8fbd9fbd9fbdefbeffb;
    inBuf[2313] = 256'h05fc21fc47fc70fc9dfccefcf9fc26fd50fd6bfd84fd9bfda4fda9fdacfda0fd;
    inBuf[2314] = 256'h93fd89fd74fd62fd56fd42fd33fd2efd20fd13fd0afdf4fcd9fcbbfc8dfc5afc;
    inBuf[2315] = 256'h22fcd6fb86fb38fbdafa7afa21fabbf95af905f9a8f852f80cf8c1f77ff74df7;
    inBuf[2316] = 256'h15f7dff6b6f680f643f609f6bff56cf51df5bff462f415f4c8f385f35af335f3;
    inBuf[2317] = 256'h21f324f322f327f33cf348f352f362f365f36bf37af37df389f3a2f3aef3c3f3;
    inBuf[2318] = 256'heaf300f41bf444f45af478f4a7f4c0f4e3f419f539f55ef591f5a8f5c4f5e8f5;
    inBuf[2319] = 256'hecf5eef5f8f5e3f5d2f5cff5aff596f592f574f55ef55df545f533f530f513f5;
    inBuf[2320] = 256'hf7f4e6f4b2f47cf44df4fcf3a8f35ff3f9f297f248f2e8f191f154f109f1cdf0;
    inBuf[2321] = 256'ha6f06ef03ef01ff0e6efaeef80ef3aeff8eec5ee7bee3bee0eeeceed98ed78ed;
    inBuf[2322] = 256'h45ed18ed00edd8ecbbecb6eca0ec96eca8ecacecbcece0ecefec02ed20ed24ed;
    inBuf[2323] = 256'h2aed3eed38ed3bed4fed52ed64ed8deda9edd8ed1cee4dee8aeed2eefdee2eef;
    inBuf[2324] = 256'h6aef87efaaefd6efe1eff6ef1bf027f03ff06bf07ef0a0f0d6f0f3f01bf153f1;
    inBuf[2325] = 256'h6df18af1b2f1b9f1c1f1d5f1caf1c4f1cef1c2f1c0f1ccf1bff1bff1cff1c4f1;
    inBuf[2326] = 256'hbff1c6f1b1f1a2f19df184f179f181f171f16ef17af16df165f166f14af12ef1;
    inBuf[2327] = 256'h17f1e4f0bbf0a3f07df06cf073f070f07ff0a6f0c0f0e0f009f11ef131f145f1;
    inBuf[2328] = 256'h3ff13ff147f13ef141f152f157f170f19cf1baf1e4f11df248f27df2bcf2e7f2;
    inBuf[2329] = 256'h1bf358f37ff3adf3e4f308f434f469f48af4b5f4eaf410f540f578f59af5c8f5;
    inBuf[2330] = 256'h02f624f651f688f6a9f6d5f60af728f74cf77af790f7a8f7c1f7c1f7c5f7cdf7;
    inBuf[2331] = 256'hc3f7c5f7d4f7d8f7ecf70ff829f854f887f8a5f8c5f8e5f8ecf8f1f8f1f8def8;
    inBuf[2332] = 256'hd0f8c8f8b7f8b5f8bff8c3f8d3f8eff802f91bf937f94bf966f982f996f9b2f9;
    inBuf[2333] = 256'hd2f9ecf910fa38fa55fa76fa97faaffaccfaeafafffa1cfb3ffb62fb8ffbc2fb;
    inBuf[2334] = 256'hf4fb2efc6bfca3fcdffc18fd4afd7ffdaffddbfd08fe2ffe53fe7efea5fec8fe;
    inBuf[2335] = 256'hf4fe24ff56ff90ffcdff10005c00a500ec00300169019a01c401e101fa011002;
    inBuf[2336] = 256'h1f0233024f026c029102bf02ee0224035d038d03be03ee031204360459047204;
    inBuf[2337] = 256'h8e04a704b604cb04dd04e304ef04fa04fc040605140520053d055d057905a405;
    inBuf[2338] = 256'hcf05ed05120630063b064d0659065206510651064a06510658065c0674068c06;
    inBuf[2339] = 256'h9c06bf06e60603072d07550774079f07c607df0700081808220835083f083f08;
    inBuf[2340] = 256'h5208650873089608bc08e1081a094e097709b109e4090a0a3d0a660a810aab0a;
    inBuf[2341] = 256'hcd0ae20a080b250b310b4c0b600b660b830b9e0bad0bd60b080c2f0c680ca10c;
    inBuf[2342] = 256'hcb0c030d2e0d400d560d5d0d4c0d470d390d1d0d180d170d110d240d350d3e0d;
    inBuf[2343] = 256'h640d850d970dbd0dd80de40d060e1e0e220e3a0e440e390e3e0e370e1d0e1b0e;
    inBuf[2344] = 256'h120efc0d050e110e150e3c0e670e860ebf0ef30e140f460f6a0f770f950fa70f;
    inBuf[2345] = 256'ha20fb50fc40fc30fdc0ff10ffc0f241047105c109010c110e1101b114a116111;
    inBuf[2346] = 256'h9011af11af11c311cb11b911bb11b511a011a611a8119e11b111be11bb11d011;
    inBuf[2347] = 256'hda11cf11da11d711c011c011b0118f1186116f1142112811fb10bd1093105810;
    inBuf[2348] = 256'h0e10e10fb00f7d0f6e0f5c0f460f4f0f500f400f430f320f090fee0ec10e7f0e;
    inBuf[2349] = 256'h530e1f0ee20dc20da00d7b0d780d730d650d750d800d7f0d960da50da70dba0d;
    inBuf[2350] = 256'hbf0db50dbd0db60d9b0d960d870d6b0d6a0d670d5a0d6d0d800d8b0db20dd40d;
    inBuf[2351] = 256'he50d070e1e0e200e300e320e1f0e180e050ee60dd70dbb0d940d830d660d410d;
    inBuf[2352] = 256'h370d2a0d140d190d190d0f0d190d170d060dff0ce30cb10c8c0c520c050cce0b;
    inBuf[2353] = 256'h8f0b480b1e0bf40ac90abc0aac0a930a930a880a6f0a6b0a5d0a3d0a2f0a180a;
    inBuf[2354] = 256'hf309da09b90991097809510922090909eb08ca08c108b808b208c608d508e208;
    inBuf[2355] = 256'h05091f0930094b09570957095f0955093f09370925090b09ff08ec08d608d608;
    inBuf[2356] = 256'hd608d508e708f90809092809430950095d095f094f0939091109de08aa086e08;
    inBuf[2357] = 256'h33080408d207a7079007790761075707440725070907e306ad0675063206e705;
    inBuf[2358] = 256'h9c054905f404a60452040004b7036d032503e802a90274024b021d02f401d301;
    inBuf[2359] = 256'haa0180015b012801f000bc007c003d000500c5ff8aff5dff2eff08fff4fee2fe;
    inBuf[2360] = 256'hd9fedefee2feedfe02ff12ff23ff39ff45ff4cff55ff54ff4cff44ff3aff32ff;
    inBuf[2361] = 256'h31ff33ff3cff4dff64ff82ffa3ffc2ffdffff7ff090016001800170013000500;
    inBuf[2362] = 256'hf5ffe8ffd3ffbcffa9ff8fff73ff5bff3dff20ff06ffe7fecbfeb8fe9dfe7ffe;
    inBuf[2363] = 256'h66fe43fe19feedfdb5fd75fd33fdeafc9dfc57fc12fcd2fb9ffb75fb53fb3efb;
    inBuf[2364] = 256'h2efb22fb1afb0ffb03fbf4fadcfabcfa9afa72fa48fa22fafef9dff9cbf9c1f9;
    inBuf[2365] = 256'hc2f9d0f9e5f901fa28fa4ffa77fa9dfab9fad3faecfaf8fa00fb0cfb0ffb15fb;
    inBuf[2366] = 256'h24fb29fb33fb48fb51fb5ffb77fb81fb8afba0fba7fbb0fbc6fbc9fbcafbd5fb;
    inBuf[2367] = 256'hcbfbbcfbb1fb8dfb64fb41fb07fbc9fa97fa56fa1afaeef9bbf98ff971f945f9;
    inBuf[2368] = 256'h1ef900f9cff89bf86ef82bf8e0f79bf744f7edf6a1f64cf600f6c4f581f547f5;
    inBuf[2369] = 256'h21f5f7f4d3f4bdf49ef481f46ff453f435f41ef4fdf3dff3c6f3a1f382f370f3;
    inBuf[2370] = 256'h55f341f33ff335f335f347f352f36af395f3b5f3dff318f446f476f4acf4cef4;
    inBuf[2371] = 256'hf1f416f522f530f545f545f54ff568f573f58af5b2f5d2f503f642f66df6a1f6;
    inBuf[2372] = 256'hdcf6fef620f740f741f743f747f730f71ef715f7f8f6e4f6dcf6c4f6baf6bdf6;
    inBuf[2373] = 256'hacf6a0f69cf683f66cf65bf632f60df6eff5baf58af566f531f503f5e1f4acf4;
    inBuf[2374] = 256'h7ff460f42ff404f4e9f3c1f3a1f390f376f363f35ef34df343f344f336f329f3;
    inBuf[2375] = 256'h26f316f308f304f3f6f2f2f2faf200f314f334f351f382f3bef3ecf322f462f4;
    inBuf[2376] = 256'h91f4c4f4fbf41ef544f570f58af5a7f5cff5ecf510f63ef663f68ef6c3f6eef6;
    inBuf[2377] = 256'h1ff758f780f7a8f7d3f7e7f7fbf712f812f812f816f806f8f8f7f2f7d7f7c2f7;
    inBuf[2378] = 256'hb9f79ef788f77cf75ef746f736f711f7f2f6dcf6aef681f65ff628f6f0f5c1f5;
    inBuf[2379] = 256'h82f547f517f5daf4a5f481f456f437f426f40bf4fdf3f9f3e4f3d5f3cdf3b3f3;
    inBuf[2380] = 256'h9ff393f375f35ef355f347f344f34ef352f369f38ef3acf3d7f30ef439f470f4;
    inBuf[2381] = 256'hadf4d9f40df546f56bf597f5c9f5e8f511f642f665f693f6cdf6faf631f775f7;
    inBuf[2382] = 256'habf7ecf733f869f8a6f8ebf81af94ef988f9abf9cff9f8f90cfa22fa39fa3cfa;
    inBuf[2383] = 256'h44fa4ffa49fa49fa53fa53fa5efa72fa7bfa8dfaa1faa7fab3fabdfaaefa9efa;
    inBuf[2384] = 256'h8dfa68fa44fa23faf5f9cff9b2f98ff979f971f962f95af95af950f94bf94af9;
    inBuf[2385] = 256'h3cf931f926f90ef9faf8e8f8cbf8b5f8a7f893f887f88bf88ef89bf8b0f8c6f8;
    inBuf[2386] = 256'he8f811f933f959f983f9a7f9ccf9eef906fa24fa44fa5cfa78fa96fab2fad8fa;
    inBuf[2387] = 256'h00fb25fb55fb8bfbbefbfcfb3efc79fcbdfc03fd3dfd79fdb1fdd9fdfefd1ffe;
    inBuf[2388] = 256'h2ffe3efe4cfe52fe5cfe6dfe7afe8bfea5febafed4fef1fe05ff18ff28ff2cff;
    inBuf[2389] = 256'h2cff29ff17ff04fff0fed2feb4fe98fe77fe5bfe43fe27fe0ffefcfde6fdd5fd;
    inBuf[2390] = 256'hc4fdaffd9efd8ffd7afd64fd4efd33fd18fdfdfce4fccdfcb6fca6fc9cfc93fc;
    inBuf[2391] = 256'h90fc93fc98fca9fcc2fcdafcf6fc18fd3bfd5cfd7dfd9afdb6fdd3fde9fdf9fd;
    inBuf[2392] = 256'h0cfe21fe39fe56fe7dfeaffee9fe28ff6cffbbff090051009900da000b013801;
    inBuf[2393] = 256'h5f0177018c01a301b501c901e001f9011a023c025c028402ac02cc02ef021103;
    inBuf[2394] = 256'h2a0341035403600369036a0365035f03520340032d031403fd02ea02d502c802;
    inBuf[2395] = 256'hbf02b402b302ba02bc02c002c502c502c502bf02b002a00287026a0254023b02;
    inBuf[2396] = 256'h200211020502fd0104020f0220023e025a0274029702b202c702e002ee02f402;
    inBuf[2397] = 256'hff02030302030c03170322033c035a037703a103d203ff03330468049904cd04;
    inBuf[2398] = 256'hfe042705520576059005ab05c005ce05df05ed05f105fe05100621063b065906;
    inBuf[2399] = 256'h7a06a606d006f606280752076c078a07a007a507aa07a4079007820772075a07;
    inBuf[2400] = 256'h4b073f07340738073b073e0750076007690779078207830785077b0768075d07;
    inBuf[2401] = 256'h460726071007f706db06cf06c106b306b706ba06b906c806d206d406e406f106;
    inBuf[2402] = 256'hef06f506fa06f806fd06f906ed06f206f306ee06f906000703071b0732074507;
    inBuf[2403] = 256'h6c079207af07db0701081d0844085f086c088408930893089f08a708a808bb08;
    inBuf[2404] = 256'hcd08db08fe08220941096b098f09ad09d609f609080a1f0a2e0a2e0a330a310a;
    inBuf[2405] = 256'h270a280a220a160a190a170a100a1d0a280a2d0a410a510a590a6c0a760a730a;
    inBuf[2406] = 256'h7b0a780a670a600a500a370a2a0a180a010afd09f409e709f009f309f109030a;
    inBuf[2407] = 256'h100a130a250a2f0a2e0a3b0a3d0a320a370a320a230a240a1c0a0d0a140a170a;
    inBuf[2408] = 256'h130a230a330a3d0a580a6d0a7b0a960aa60aaa0abb0ac00aba0ac10abe0ab10a;
    inBuf[2409] = 256'hb50ab40aab0aba0ac40ac90ae70a010b110b350b530b660b870b9e0ba40bb70b;
    inBuf[2410] = 256'hbf0bb90bbf0bba0bac0bb10bb00ba80bb70bc50bca0be40bfc0b0c0c2d0c460c;
    inBuf[2411] = 256'h530c700c840c8b0ca10ca90ca10caa0caa0c970c920c890c740c6e0c610c4b0c;
    inBuf[2412] = 256'h4d0c4b0c420c4c0c510c4c0c590c5b0c4f0c500c400c1c0c0b0cef0bc00ba30b;
    inBuf[2413] = 256'h800b530b3c0b200bfc0af00ae10ac70ac30ab80a9e0a950a800a5f0a500a320a;
    inBuf[2414] = 256'h060aee09d009a7099309790959094e093d092a092e092b0922092e0933093009;
    inBuf[2415] = 256'h410945093d0947094a0943094c094b094009440945093e094409480949095709;
    inBuf[2416] = 256'h62096d098909a109b309d109e809f6090a0a130a100a140a0b0af809ef09db09;
    inBuf[2417] = 256'hc309bc09b209a309a509a509a109a809a4099609940984096609510932090709;
    inBuf[2418] = 256'he308b9088808610832080108dd07b00781075f0731070107e006b7068c066c06;
    inBuf[2419] = 256'h44061b06fd05d405aa058c05620532051005e404b40492046c0444042b041304;
    inBuf[2420] = 256'hfa03ef03e703dd03dd03da03d403d403ce03bf03b703ae039e0394038f038b03;
    inBuf[2421] = 256'h91039903a403ba03d203ea0306041e04310442044f0457045e045c0457045804;
    inBuf[2422] = 256'h54044e044f044a0442043d0433042804230416040604f903e803d603c303ab03;
    inBuf[2423] = 256'h9203760350032903f902be0283024502fc01b50170012501dd00990055001800;
    inBuf[2424] = 256'hddffa1ff6aff30fff1feb3fe70fe26fedefd95fd48fdfffcb7fc6efc2bfceefb;
    inBuf[2425] = 256'hb6fb85fb57fb2dfb0afbe8fac8faaefa94fa77fa5ffa47fa2efa1cfa09faf5f9;
    inBuf[2426] = 256'heaf9e3f9dcf9dcf9def9e1f9ebf9f5f905fa1bfa2bfa3efa5bfa6ffa82fa9dfa;
    inBuf[2427] = 256'haefabbfad0fadafae0faeafaeafae7faebfae5fae2fae9fae6fae4faedfaebfa;
    inBuf[2428] = 256'he8faecfae0fad2fac8faabfa8bfa6efa3cfa09fae1f9a8f96df93df902f9ccf8;
    inBuf[2429] = 256'ha1f868f835f80ef8d9f7a7f77ff744f70cf7e2f6a4f663f630f6eff5aff57af5;
    inBuf[2430] = 256'h3bf500f5d5f4a0f46ff44df422f400f4edf3d1f3bff3b9f3a5f39af3a0f395f3;
    inBuf[2431] = 256'h8ef397f38ff38bf397f393f395f3a8f3abf3b6f3d1f3e1f3faf324f440f463f4;
    inBuf[2432] = 256'h92f4aef4cef4fcf414f52bf54bf557f568f582f587f595f5aef5b3f5c2f5dff5;
    inBuf[2433] = 256'he4f5f2f50cf60bf60ff620f616f60ef610f6f3f5d7f5c8f59ef576f55bf526f5;
    inBuf[2434] = 256'hf6f4d5f4a0f470f44ef419f4ecf3cff39bf36ff351f31bf3eaf2c8f28ff25af2;
    inBuf[2435] = 256'h31f2f2f1b9f191f155f11ef1f8f0c4f099f07ef056f03bf032f019f00bf00ff0;
    inBuf[2436] = 256'h05f000f00af004f006f013f011f015f025f027f035f051f05ef077f09ef0baf0;
    inBuf[2437] = 256'he2f019f13df16cf1a8f1cff1fcf134f257f282f2b6f2d2f2f6f225f33ff366f3;
    inBuf[2438] = 256'h98f3b1f3d8f30bf423f446f477f48df4adf4d9f4e7f4faf41bf521f52af53cf5;
    inBuf[2439] = 256'h35f534f53bf52bf523f523f50df504f507f5f2f4e9f4eef4dff4d7f4d9f4c9f4;
    inBuf[2440] = 256'hc0f4bef4a7f494f489f46ef45bf44df430f41df414f400f4fdf304f4fef307f4;
    inBuf[2441] = 256'h1cf421f431f44ef45cf472f48ff49ff4b5f4d5f4e8f405f52cf547f56cf599f5;
    inBuf[2442] = 256'hbdf5edf524f64df683f6c2f6f3f62ef771f7a7f7e7f72cf85ff899f8d8f809f9;
    inBuf[2443] = 256'h44f97ff9a9f9dcf914fa39fa68fa9cfac3faf1fa24fb48fb71fb9bfbb7fbd7fb;
    inBuf[2444] = 256'hf4fb02fc14fc26fc28fc2dfc36fc34fc37fc3efc3cfc3efc44fc43fc48fc4ffc;
    inBuf[2445] = 256'h4dfc4bfc4afc43fc3cfc34fc26fc1cfc11fcfffbf4fbeafbdbfbd2fbcefbc8fb;
    inBuf[2446] = 256'hc9fbcefbd1fbdcfbecfbfbfb0ffc23fc36fc51fc6bfc82fc9dfcb7fccefceafc;
    inBuf[2447] = 256'h06fd21fd41fd64fd87fdb4fde0fd0cfe40fe74fea7fedffe14ff47ff7cffadff;
    inBuf[2448] = 256'hd9ff080033005c008700ae00d400fd0026014e017a01a601d001f8011d024402;
    inBuf[2449] = 256'h69028802a902c802dd02f3020a031b032b033d03490356036603700379038503;
    inBuf[2450] = 256'h8d039903a803b203be03ce03d903e403f003f503fd030604030405040c040704;
    inBuf[2451] = 256'h06040d040f04150420042a043d045304610478049104a104b704cd04dc04f004;
    inBuf[2452] = 256'h01050a051e0530053d0557056e057c059805b805cd05ec050e0628064c067006;
    inBuf[2453] = 256'h8d06b306d706f30619073a0750076f078b079e07b607c807d307e907fc070808;
    inBuf[2454] = 256'h1f08340843085b086f087c089308a208a808b908c208c208cc08ce08c808d108;
    inBuf[2455] = 256'hd408cc08d408d808d008d408d408c808c908c608b308ab08a208900887087c08;
    inBuf[2456] = 256'h6b0867085d084d084a084208340835082e082108250821081708220823081c08;
    inBuf[2457] = 256'h2c083708360846084f084c08590861085c0867086d086a087708800881089408;
    inBuf[2458] = 256'ha408ad08c608d908e208fa080b091209260934093a094c0959095e0970097a09;
    inBuf[2459] = 256'h7d0990099a099909a409a7099e09a309a1099309950990097e097b0975096809;
    inBuf[2460] = 256'h66095f094e0948093e09290920091309fd08f108df08c708bf08b408a1089908;
    inBuf[2461] = 256'h8d087908710864084e0844083608210818080a08f807f307e907dd07e007da07;
    inBuf[2462] = 256'hce07d307d007c507c807c407b807be07bd07b707c307c907c707d607de07df07;
    inBuf[2463] = 256'hf007f807f80707080a080608100810080808120814080e08150814080d081208;
    inBuf[2464] = 256'h0d0800080008f707e807e207d407c407c007b1079f079c079107800778076607;
    inBuf[2465] = 256'h50074707350718070207e806c806b30695066f06550637061006f105cf05a905;
    inBuf[2466] = 256'h8c056a05440529050905e604d004b7049a04890476045f0451043e042a041e04;
    inBuf[2467] = 256'h0b04f403e903d903c403b903aa0398038f038303750371036a0361035f035903;
    inBuf[2468] = 256'h5303550353035003560359035a03620367036c0377037e0383038c038f039303;
    inBuf[2469] = 256'h9b039e039f03a403a2039d039c0395038a037f037203610350033a0323030e03;
    inBuf[2470] = 256'hf402dc02c702b002990284026c02510238021d020102e301c1019f017b015201;
    inBuf[2471] = 256'h2a010101d300a8007e0050002400faffcdffa3ff7bff50ff2aff08ffe3fec0fe;
    inBuf[2472] = 256'ha1fe82fe66fe4dfe32fe1afe06feeefddbfdccfdbefdb5fdadfda6fda5fda6fd;
    inBuf[2473] = 256'ha6fdabfdb4fdbafdc2fdcafdd0fdd8fde1fde5fde9fdeffdf4fdfcfd04fe0efe;
    inBuf[2474] = 256'h1bfe26fe31fe41fe4dfe56fe64fe70fe7bfe88fe8ffe93fe99fe9bfe9bfe9cfe;
    inBuf[2475] = 256'h97fe8ffe88fe79fe66fe54fe3bfe1ffe06fee6fdc5fdabfd89fd67fd4afd24fd;
    inBuf[2476] = 256'hfefcdefcb6fc8cfc67fc3afc0dfce8fbbbfb8dfb6afb43fb1efb02fbe5facafa;
    inBuf[2477] = 256'hb2fa94fa7afa63fa45fa28fa0ffaeff9d2f9bcf9a2f98ff980f96ef965f966f9;
    inBuf[2478] = 256'h60f960f96af970f97af98af996f9a9f9c0f9d3f9eff90efa26fa42fa60fa76fa;
    inBuf[2479] = 256'h92faaefabefad4faeefafbfa0afb1ffb2dfb3ffb53fb5dfb70fb85fb8afb95fb;
    inBuf[2480] = 256'ha7fba9fbacfbb4fbaefbacfbb0fba7fba2fba5fb99fb8ffb8ffb80fb70fb65fb;
    inBuf[2481] = 256'h4bfb30fb19fbf3faccfaabfa7efa52fa2cfafbf9ccf9a5f974f946f920f9f2f8;
    inBuf[2482] = 256'hc8f8a7f87ef859f83ef81df8fff7ecf7d5f7c2f7b3f79df78cf781f76df75bf7;
    inBuf[2483] = 256'h4ef73cf72cf725f71bf716f718f719f720f72df739f74cf761f771f789f7a3f7;
    inBuf[2484] = 256'hb5f7d0f7f0f709f82bf854f875f89df8ccf8f5f826f959f980f9adf9ddf900fa;
    inBuf[2485] = 256'h24fa4cfa68fa86faa4fab9fad3faecfaf9fa0afb1efb25fb30fb3efb3efb43fb;
    inBuf[2486] = 256'h4afb46fb47fb4dfb44fb40fb40fb37fb30fb2afb18fb09fbfafadffac7fab2fa;
    inBuf[2487] = 256'h92fa75fa5bfa38fa1bfa01fadff9c5f9aff98ff977f967f94df938f92bf919f9;
    inBuf[2488] = 256'h0df908f900f9fff803f906f912f922f932f94bf965f97cf99bf9bbf9d7f9fbf9;
    inBuf[2489] = 256'h1ffa3efa65fa8cfaacfad3fafbfa1cfb44fb6efb93fbc0fbedfb14fc44fc76fc;
    inBuf[2490] = 256'ha2fcd6fc0dfd3cfd6efda1fdccfdfafd26fe49fe70fe93fea9fec1fed9fee8fe;
    inBuf[2491] = 256'hf6fe02ff07ff0dff10ff0bff09ff04fff5fee9fedcfec8feb7fea5fe8dfe79fe;
    inBuf[2492] = 256'h67fe52fe40fe30fe1dfe0ffe01feeffde0fdd4fdc3fdb1fda0fd8efd7efd6afd;
    inBuf[2493] = 256'h55fd43fd32fd1ffd10fd01fdf3fce9fce0fcd9fcd8fcd9fcddfce6fcf0fcfffc;
    inBuf[2494] = 256'h14fd2bfd45fd62fd7ffd9efdc0fde2fd07fe2cfe4efe74fe9afebbfedefe05ff;
    inBuf[2495] = 256'h26ff48ff6eff91ffb5ffdbfffdff1f00430066008800ad00cd00ee0012013301;
    inBuf[2496] = 256'h520173019201b201d401f201120231024d026b0285029902ab02bb02c502cf02;
    inBuf[2497] = 256'hd502d402d402d402cd02c702c202bb02b502b002ab02aa02a802a402a302a002;
    inBuf[2498] = 256'h9c029f02a1029f02a402a702a602ad02b402b602be02c402c502cd02d302d302;
    inBuf[2499] = 256'hdd02e502e502ed02f802fd02070312031a032a033b0346035a03710382039c03;
    inBuf[2500] = 256'hb903d003f10314043004530476049504b804d804f1040d05280539054c055f05;
    inBuf[2501] = 256'h6a0573057c0583058a058e058e059005920591059105920590058e058c058805;
    inBuf[2502] = 256'h8705830580057e05790571056c05620556054c053d052a0519050305ea04d504;
    inBuf[2503] = 256'hbb04a0048a046f0453043c0421040304eb03d203b803a50392037f0372036503;
    inBuf[2504] = 256'h5b035a03560354035a035a0358035f035f0359035a0355034b0347033e033203;
    inBuf[2505] = 256'h2e0326031c031c031a03140317031803150319031c031d0327032d032e033a03;
    inBuf[2506] = 256'h45034b035a0367036f037f038b039203a103ab03ae03b803c003c203c803cd03;
    inBuf[2507] = 256'hcd03d303d403d203d803d803d403d903dc03dd03e603ed03f203020411041e04;
    inBuf[2508] = 256'h36044b045c0476048d049d04b504ca04d804ea04fa0402050f0519051e052705;
    inBuf[2509] = 256'h2e05300538053c053d054805500552055c0567056f057e058a059305a205ac05;
    inBuf[2510] = 256'hb305c005c805cc05d505da05db05e105e305e005e205e105dc05da05d205c505;
    inBuf[2511] = 256'hbb05ab05970585056d055405400527050f05fd04e804d404c804ba04ac04a304;
    inBuf[2512] = 256'h97048a048304770467045c044e043b0429041404ff03ea03cf03b20399037c03;
    inBuf[2513] = 256'h5d03410324030703ed02d102b602a1028c027702670257024602380228021b02;
    inBuf[2514] = 256'h0f02ff01f201e701da01cd01c101b301a50199018801760164014e0138012201;
    inBuf[2515] = 256'h0801ee00d400b8009f0087006d00580043002b0017000500f2ffe3ffd5ffc4ff;
    inBuf[2516] = 256'hb8ffaeffa0ff94ff88ff78ff69ff5aff45ff30ff19fffcfee0fec4fea3fe84fe;
    inBuf[2517] = 256'h69fe4cfe33fe1dfe08fef7fde9fdd9fdccfdc2fdb6fdaefda7fd9ffd98fd95fd;
    inBuf[2518] = 256'h93fd92fd96fd9cfda2fdadfdb8fdc3fdcefdd9fde1fdebfdf5fdfbfd02fe0bfe;
    inBuf[2519] = 256'h15fe1ffe2dfe3cfe4efe63fe78fe91feaffeccfeeafe0dff2eff50ff76ff9cff;
    inBuf[2520] = 256'hc1ffeaff120037005e008300a400c400e000f7000e01220130013f014e015901;
    inBuf[2521] = 256'h640171017c01870193019c01a601ae01b301b801bc01bb01b901b801b401af01;
    inBuf[2522] = 256'hab01a6019f0198018f01830176016701550141012a011101f700db00bd009f00;
    inBuf[2523] = 256'h81006200430025000600e8ffcbffaeff95ff7dff67ff54ff44ff36ff2bff22ff;
    inBuf[2524] = 256'h1bff14ff0cff02fff8feeafedbfecafeb7fea2fe8dfe77fe63fe50fe3dfe2dfe;
    inBuf[2525] = 256'h21fe12fe04fefbfdeefddffdd4fdc5fdb6fdaafd9afd8cfd82fd75fd67fd60fd;
    inBuf[2526] = 256'h53fd43fd3afd2afd15fd03fdeafccefcb4fc92fc6efc50fc2dfc06fce5fbbdfb;
    inBuf[2527] = 256'h94fb73fb4bfb1ffbf9facefaa1fa7dfa53fa29fa0afae8f9c5f9adf992f977f9;
    inBuf[2528] = 256'h62f94af92ef918f9fcf8ddf8c1f8a0f880f864f845f828f811f8f9f7e5f7d7f7;
    inBuf[2529] = 256'hc8f7c0f7bcf7b7f7b8f7bdf7bff7c9f7d7f7e4f7f9f711f828f848f868f886f8;
    inBuf[2530] = 256'haff8d8f8fbf828f957f980f9b1f9e3f911fa47fa7cfaaefae9fa23fb57fb95fb;
    inBuf[2531] = 256'hd2fb08fc47fc85fcbdfcfffc42fd80fdc6fd0bfe4cfe96feddfe1eff65ffa9ff;
    inBuf[2532] = 256'he4ff22005d009000c500f4001d0148016f019001b601d601f2010f0229023e02;
    inBuf[2533] = 256'h54026802780289029602a302b102bc02c702d402dd02e702f002f502fa02fd02;
    inBuf[2534] = 256'hfa02f902f602ed02e602de02d202c802bf02b202a8029d028f02830276026402;
    inBuf[2535] = 256'h550248023702270219020c020002f601ef01e901e301df01dd01d701d201ca01;
    inBuf[2536] = 256'hbf01b301a4018f017b01640147012c010e01ec00cd00ab00840061003a000f00;
    inBuf[2537] = 256'he9ffbdff8bff61ff31fffafecbfe97fe5dfe2bfef4fdb6fd81fd45fd02fdc9fc;
    inBuf[2538] = 256'h89fc41fc02fcbefb72fb30fbe9fa9bfa57fa0efac2f980f938f9eff8b1f86ef8;
    inBuf[2539] = 256'h2bf8f2f7b7f77cf74bf719f7ebf6c4f69cf67af660f643f62df61ef60df602f6;
    inBuf[2540] = 256'hfcf5f4f5f2f5f5f5f4f5fcf508f60ff622f638f64bf66af68df6aef6dcf60df7;
    inBuf[2541] = 256'h3cf77bf7b9f7f5f741f88cf8d2f827f97cf9cbf927fa80fad5fa36fb94fbebfb;
    inBuf[2542] = 256'h51fcb2fc0dfd74fdd7fd33fe9cfefffe5dffc6ff27008400ec004b01a5010a02;
    inBuf[2543] = 256'h6602be0220037b03d20331048704dd043a058c05de0534067e06c80615075507;
    inBuf[2544] = 256'h9507d6070b08410876089f08cc08f80818093c09600979099609b209c309db09;
    inBuf[2545] = 256'hf009fa090d0a1c0a210a2e0a380a390a420a460a420a430a3d0a300a290a180a;
    inBuf[2546] = 256'h000aed09d209b209960973094c092a090009d508ae087e084d082008e807af07;
    inBuf[2547] = 256'h78073607f506b6066c062506e10591054705fe04aa045c040f04b4035e030703;
    inBuf[2548] = 256'ha3024402e20174010d01a3002e00c3ff57ffe1fe76fe0afe96fd2cfdc1fc4ffc;
    inBuf[2549] = 256'he8fb7efb0efbabfa45fadaf97bf91af9b6f85ef802f8a5f753f7fcf6a5f659f6;
    inBuf[2550] = 256'h07f6b7f573f529f5e4f4abf46ef438f40df4dff3b9f39ef37ef367f35bf349f3;
    inBuf[2551] = 256'h41f341f33df345f353f35df376f394f3adf3d6f303f42af461f49bf4d0f413f5;
    inBuf[2552] = 256'h57f597f5e6f534f67ef6d8f631f786f7ebf74df8adf81df989f9f4f970fae6fa;
    inBuf[2553] = 256'h5cfbe4fb65fce6fc78fd02fe8bfe23ffb0ff3c00d5005f01ea01810208039103;
    inBuf[2554] = 256'h2604ac043505cb055306de067407fa078508170998091c0aa60a1e0b980b170c;
    inBuf[2555] = 256'h840cf50c6a0dcd0d360ea10efa0e590fb70f04105410a210de101d1157118011;
    inBuf[2556] = 256'had11d311e911051217121b122512241216120c12f711d611ba1191115e113311;
    inBuf[2557] = 256'hf810b7107e103610e80fa20f4b0fef0e980e300ec30d5b0ddf0c610ce80b5d0b;
    inBuf[2558] = 256'hd20a4e0abb092a09a1080a087807ed065406c1053405980401047103d2023902;
    inBuf[2559] = 256'ha60107016f00ddff40ffaefe20fe8afdfefc77fce7fb63fbe1fa59fadcf95ff9;
    inBuf[2560] = 256'hdcf865f8ebf770f700f78ff61df6b7f550f5eaf492f437f4e0f398f34bf304f3;
    inBuf[2561] = 256'hccf28ef256f22bf2faf1cff1aef186f165f14ef12ef117f109f1f4f0e9f0e9f0;
    inBuf[2562] = 256'he3f0e7f0f6f000f117f135f14ff177f1a4f1ccf103f23ef275f2b9f202f348f3;
    inBuf[2563] = 256'h9cf3f1f346f4aaf40df570f5e3f553f6c4f644f7c1f740f8cef856f9e1f97bfa;
    inBuf[2564] = 256'h0dfba2fb47fce0fc7dfd29fec9fe6dff1f00c4006f012902d40287034804fa04;
    inBuf[2565] = 256'hb20577062a07e207a3085109020ab80a590bfe0ba70c3a0dd20d6e0ef60e830f;
    inBuf[2566] = 256'h131091101311961106127a12ea124613a613fd1340148614c214eb1416153715;
    inBuf[2567] = 256'h47155b1562155b155a1549152b151215e914b41483144014f213a9134c13e612;
    inBuf[2568] = 256'h87121212961123119a100d10890ff20e580ec90d270d860cf00b460ba00a060a;
    inBuf[2569] = 256'h5909af0810085f07b2060f065905a90403044c039c02f80143019900faff4fff;
    inBuf[2570] = 256'haffe1afe7bfde9fc60fccdfb49fbcbfa43fac9f954f9d6f866f8f9f786f71ff7;
    inBuf[2571] = 256'hbbf653f6f9f5a0f544f5f9f4adf45ff421f4e1f3a1f36ef337f300f3d4f2a3f2;
    inBuf[2572] = 256'h72f24ef221f2f6f1daf1b5f194f182f16af158f154f14bf14af155f159f165f1;
    inBuf[2573] = 256'h7bf189f19ef1bbf1d0f1ebf10df228f24df277f29cf2ccf203f335f375f3bbf3;
    inBuf[2574] = 256'hfdf34df4a0f4f1f44ff5aef50bf676f6def645f7baf72cf89ef81df997f913fa;
    inBuf[2575] = 256'h9efa21fba6fb3afcc5fc52fdeefd80fe14ffb6ff4b00e30087011d02b5025803;
    inBuf[2576] = 256'hec0381042005af053f06d8066207ef07830807098f091c0a990a190b9d0b0f0c;
    inBuf[2577] = 256'h830cf60c580db90d170e640eb20efa0e310f6a0f9d0fc20fe90f0a101e103710;
    inBuf[2578] = 256'h47104b105410511043103a1023100110e30fb60f7f0f4c0f090fc00e7c0e290e;
    inBuf[2579] = 256'hd00d7f0d200dbe0c620cf70b8b0b270bb20a3b0acb094a09c9084e08c3073807;
    inBuf[2580] = 256'hb506230695050f057c04ee036a03db025302d2014601c2004400baff3affbefe;
    inBuf[2581] = 256'h36feb7fd3cfdb7fc3bfcc2fb41fbcbfa57fadcf96ef901f98ef828f8c3f75af7;
    inBuf[2582] = 256'hfff6a2f643f6f1f59bf543f5f9f4aaf458f414f4caf37ef341f3fcf2b8f283f2;
    inBuf[2583] = 256'h49f211f2e7f1b7f18bf16ff14cf12bf118f1fcf0e6f0daf0c4f0b4f0aef09ef0;
    inBuf[2584] = 256'h96f099f092f094f0a3f0abf0bef0dcf0f2f016f142f166f198f1d2f101f23bf2;
    inBuf[2585] = 256'h7bf2b2f2f5f23af377f3c1f30df451f4a5f4faf447f5a7f508f663f6cef639f7;
    inBuf[2586] = 256'h9df711f882f8edf867f9daf946fabffa33fb9efb17fc8afcf7fc71fde5fd54fe;
    inBuf[2587] = 256'hcffe43ffb4ff3100a50014018d01fc016702d8024003a3030b046a04c6042605;
    inBuf[2588] = 256'h7b05cf0527067606c30614075d07a507ef0730087208b508ef08280960098f09;
    inBuf[2589] = 256'hbd09e709080a290a460a5a0a6d0a7a0a810a890a8d0a8c0a8c0a870a7e0a780a;
    inBuf[2590] = 256'h6b0a5b0a4c0a330a170afc09d409aa0980094a091209db08990857081608cc07;
    inBuf[2591] = 256'h83073d07ed069f065206fa05a7055105f00492043304c8036203f80283021602;
    inBuf[2592] = 256'ha6012d01bc004900ceff5effeafe6ffefffd8cfd12fda4fc31fcb5fb46fbd5fa;
    inBuf[2593] = 256'h5afaebf97af903f998f828f8b6f752f7e9f67ef623f6c5f565f512f5bef46bf4;
    inBuf[2594] = 256'h24f4d8f390f354f312f3d3f2a1f269f234f20cf2ddf1b4f198f176f15cf14ef1;
    inBuf[2595] = 256'h39f12ef12ff129f12cf13af140f151f16bf17af194f1b5f1ccf1eff119f238f2;
    inBuf[2596] = 256'h62f294f2bcf2f0f22cf35ef39cf3e1f31df466f4b3f4f5f444f597f5dcf52ef6;
    inBuf[2597] = 256'h82f6c9f61bf770f7b9f70cf862f8aef805f95df9aff90afa66fabbfa19fb76fb;
    inBuf[2598] = 256'hcefb2dfc88fcdefc3bfd93fde8fd43fe98feebfe46ff9cfff1ff4c00a300fc00;
    inBuf[2599] = 256'h5a01b3010d026c02c4021e037c03cf0324047f04d00421057405c0050e065d06;
    inBuf[2600] = 256'ha406ee0639077d07c307080847088a08ca08040940097909aa09dd090d0a340a;
    inBuf[2601] = 256'h5e0a820a9e0aba0acf0ade0aef0af90afd0a030b020bfc0af60ae90adb0acc0a;
    inBuf[2602] = 256'hb20a960a7a0a500a250af909be0983094809fe08b6086f081a08c80779071d07;
    inBuf[2603] = 256'hc60670060e06b3055805ef048b042904b8034c03e2026d02fd018d0111019d00;
    inBuf[2604] = 256'h2d00b5ff43ffd5fe5efef1fd88fd19fdb2fc4efce5fb86fb2dfbcdfa74fa21fa;
    inBuf[2605] = 256'hc9f979f92df9e1f89cf859f818f8e0f7a9f775f74af724f701f7e4f6c8f6b2f6;
    inBuf[2606] = 256'ha4f695f68af686f680f67ff686f68af693f6a3f6b1f6c7f6e3f6fcf61df745f7;
    inBuf[2607] = 256'h6af797f7c8f7f7f72df867f89df8d9f817f951f991f9d1f90cfa4efa8ffacafa;
    inBuf[2608] = 256'h0dfb50fb8efbd3fb18fc5bfca5fcedfc36fd86fdd3fd1efe6ffebefe0dff5eff;
    inBuf[2609] = 256'habfff9ff48009100de002f017801c60117026002b00204034f03a103f5033e04;
    inBuf[2610] = 256'h8d04df0425057305c00501064c069906d7061d076607a507ed0736087408ba08;
    inBuf[2611] = 256'h00093c098109c509fe093d0a7c0ab00aea0a1f0b4a0b7b0ba70bc70bef0b120c;
    inBuf[2612] = 256'h2b0c490c610c700c870c970ca00cb00cb90cba0cc20cc10cb90cb60ca80c960c;
    inBuf[2613] = 256'h8a0c6e0c4c0c300c080cdc0bb30b7b0b430b120bd20a900a540a090abf097c09;
    inBuf[2614] = 256'h2809d40885082708c80770070a07a5064506d9056f050c059d043104ce036303;
    inBuf[2615] = 256'hfc029a023102cc016c010601a2004600e5ff83ff27ffc8fe6afe10feb7fd63fd;
    inBuf[2616] = 256'h12fdbffc73fc2dfce8fba9fb71fb3dfb0cfbe1fabafa99fa7dfa65fa50fa3efa;
    inBuf[2617] = 256'h30fa25fa1ffa1efa1efa22fa2bfa36fa45fa5bfa70fa89faabfaccfaedfa19fb;
    inBuf[2618] = 256'h43fb6bfb9cfbcdfbfcfb33fc67fc9cfcd8fc11fd4bfd8efdccfd0cfe55fe96fe;
    inBuf[2619] = 256'hd9fe27ff6dffb2ff000047008c00d8001b015c01a101df011b025b029302c902;
    inBuf[2620] = 256'h020334036903a103d10306043f046d04a104da0408053a056f059805c705f705;
    inBuf[2621] = 256'h1a0642066c068b06ab06cd06e806070725073c07590775078907a207ba07cc07;
    inBuf[2622] = 256'he307f6070208140822082a0838084308470852085b085e0867086c086d087408;
    inBuf[2623] = 256'h7608720874087108680865085a0849083d0829081008fb07de07bb079d077607;
    inBuf[2624] = 256'h4d072807fa06cb06a20670063e061106db05a50573053805fc04c2047e043904;
    inBuf[2625] = 256'hf403a60359030c03b4025f020c02b1015601fe00a0004500e9ff89ff2dffd0fe;
    inBuf[2626] = 256'h6ffe14feb6fd54fdf8fc9cfc3efce7fb8dfb36fbe6fa93fa40faf9f9b3f96bf9;
    inBuf[2627] = 256'h2cf9eef8b2f87df847f815f8eaf7bef796f773f750f732f71af701f7eff6e4f6;
    inBuf[2628] = 256'hd6f6d3f6d8f6ddf6ecf602f717f736f75cf782f7aef7e0f711f847f881f8bbf8;
    inBuf[2629] = 256'hfaf838f978f9c0f907fa4cfa9afae6fa30fb83fbd3fb22fc7afccefc1ffd76fd;
    inBuf[2630] = 256'hcbfd1efe76fec9fe1bff73ffc1ff10006500b100fa004b019401d90127026a02;
    inBuf[2631] = 256'ha802ed022b036603a403d90309043a0462048704ae04cc04e504000514052405;
    inBuf[2632] = 256'h36054805570562056a0576057f0584058c05920592058f058b0584057b056d05;
    inBuf[2633] = 256'h5e0550053c0522050a05ef04d304b704970478045b0438041504f403cf03ab03;
    inBuf[2634] = 256'h8903660341031b03f202cc02a7027e0256022e020002d701b101830155012a01;
    inBuf[2635] = 256'hfd00d200a4006f003f000e00d5ffa1ff6bff2ffff5febafe7afe3dfefdfdbafd;
    inBuf[2636] = 256'h7dfd3efdfbfcbffc7efc3cfc02fcc4fb82fb49fb0cfbcafa8ffa4efa0cfad0f9;
    inBuf[2637] = 256'h8cf945f909f9c7f883f847f806f8c2f788f74cf713f7e0f6a7f674f64bf61cf6;
    inBuf[2638] = 256'hf0f5cdf5a7f586f56df54ff537f526f50ff502f5fdf4f2f4eff4f2f4f0f4f8f4;
    inBuf[2639] = 256'h08f512f526f540f554f56ff592f5b2f5daf506f62ef660f696f6c7f603f744f7;
    inBuf[2640] = 256'h81f7c8f711f859f8abf8fdf84bf9a4f9fef952fab0fa0cfb62fbc3fb1efc73fc;
    inBuf[2641] = 256'hd4fc30fd82fdddfd36fe86fedffe32ff7dffd3ff24006b00ba00050147019101;
    inBuf[2642] = 256'hd701130253028f02c602ff0231035b038703af03d003f0030c04230439044904;
    inBuf[2643] = 256'h53045d04620463046404600456044704370424040e04f703db03bb039e038003;
    inBuf[2644] = 256'h5b0337031003e702c1029d02720247021c02ed01c1019301620135010701d100;
    inBuf[2645] = 256'h9e006e0038000500d2ff9fff6fff3eff0bffddfeaffe7efe54fe2afefffdd8fd;
    inBuf[2646] = 256'hb3fd8cfd6cfd4afd23fd04fde7fcc6fca9fc8dfc6efc52fc36fc17fcfefbe4fb;
    inBuf[2647] = 256'hc9fbb3fb9afb7efb68fb4ffb37fb24fb0cfbf4fae3facafab2faa2fa8dfa76fa;
    inBuf[2648] = 256'h69fa54fa3ffa35fa23fa0efa06fafaf9e7f9dbf9cdf9bff9b6f9a8f999f991f9;
    inBuf[2649] = 256'h83f976f96ef961f955f950f947f940f93df939f939f93df93ef944f94ff956f9;
    inBuf[2650] = 256'h63f975f983f995f9abf9bef9d7f9f3f90afa27fa49fa64fa85faadfad0faf7fa;
    inBuf[2651] = 256'h23fb4dfb7afbaafbdafb0cfc41fc75fcadfce6fc1bfd57fd94fdcffd0efe4cfe;
    inBuf[2652] = 256'h87fec9fe0cff49ff8bffcbff070047008900c800090145017e01bb01f5012a02;
    inBuf[2653] = 256'h62029502c402f50223034c0374039903bd03e103030422043f04590473048a04;
    inBuf[2654] = 256'h9c04b004c004c904d304dc04e004e104de04d804d304c804ba04af04a1048c04;
    inBuf[2655] = 256'h79046504500439041e040504ef03d203b4039703770359033e031b03f902dc02;
    inBuf[2656] = 256'hba0298027a02570237021e020002e001c601aa018f0179015e01460134011e01;
    inBuf[2657] = 256'h0501f400e200cc00bc00ae009f00920086007b0073006c006600630060006000;
    inBuf[2658] = 256'h62006400660069006c0073007c00820088008e0093009c00a800b000b700c000;
    inBuf[2659] = 256'hc900d400e000eb00f800060112011e012901340140014c0154015e0168016f01;
    inBuf[2660] = 256'h74017c01830188018d019101960199019c019e01a001a101a201a501a501a101;
    inBuf[2661] = 256'h9e019a01960192018d0185017f0176016d0167015e01550151014b0143013c01;
    inBuf[2662] = 256'h36012f012b01260122011f011901130112010f010a0109010801040106010a01;
    inBuf[2663] = 256'h0a010a010e0116011e0124012b01350140014a015801670173017f018d019b01;
    inBuf[2664] = 256'hab01bd01cc01dc01ee01ff0115022a023a0250026a0280029802b002c402dc02;
    inBuf[2665] = 256'hf8020f03230338034c036303780388039c03b003c003d303e403f10304041604;
    inBuf[2666] = 256'h2204340441044a045a0467046c047804820486048f04960496049b04a104a004;
    inBuf[2667] = 256'ha304a604a604a904a904a504a704a804a304a704a7049f049e049c0496049704;
    inBuf[2668] = 256'h94048c048e048e0488048c048d0488048f04970498049f04a404a704b904c404;
    inBuf[2669] = 256'hc404d304e304e804f60401050705180525052c053e054c055405660576058005;
    inBuf[2670] = 256'h9305a505b005c005cd05d905eb05f405fa050a06130617061f0621061d062106;
    inBuf[2671] = 256'h21061d061d0613060306fc05ee05da05cb05b7059b058105630542052005f904;
    inBuf[2672] = 256'hd204aa04780448041d04e703b00380034a030f03d8029b025f022502e401a401;
    inBuf[2673] = 256'h67012201df009c0053000e00cdff84ff3ffffdfeb7fe76fe36fef2fdb8fd80fd;
    inBuf[2674] = 256'h42fd0efddefca8fc78fc4efc22fcfcfbdafbb6fb9afb80fb64fb51fb44fb33fb;
    inBuf[2675] = 256'h26fb20fb1cfb1cfb20fb27fb31fb3ffb51fb64fb79fb93fbaffbcefbedfb0ffc;
    inBuf[2676] = 256'h38fc62fc88fcb6fceafc19fd4dfd89fdbefdf6fd39fe76feb1fef2fe2dff6aff;
    inBuf[2677] = 256'hadffe8ff240064009d00d700150146017801b501ec011c0251028202b302e602;
    inBuf[2678] = 256'h12033f036f039703bd03eb0310043104560473048b04aa04c704dd04f1040505;
    inBuf[2679] = 256'h1b052c053805470553055e056a05730577058105860585058805880584058605;
    inBuf[2680] = 256'h85057f057d05770571056f056a056505630559054f054e0547053c0534052605;
    inBuf[2681] = 256'h19050d05f704e304d304ba04a1048b046d044f0435041204f203d403ad038903;
    inBuf[2682] = 256'h66033c031603ed02bb028c025d022702f201bb017c0140010101bc0079003200;
    inBuf[2683] = 256'he8ffa0ff50fffefeb5fe63fe0bfebcfd64fd09fdb7fc5ffc01fcaffb56fbf7fa;
    inBuf[2684] = 256'h9efa43fae9f99af943f9ebf8a0f850f8fef7b9f770f726f7e8f6a7f664f62df6;
    inBuf[2685] = 256'hf6f5c0f591f560f534f512f5edf4cef4bbf4a3f491f48cf488f489f493f49df4;
    inBuf[2686] = 256'hadf4c9f4e6f409f531f55af58ff5c6f5faf53af67df6bef60bf75af7a5f7fcf7;
    inBuf[2687] = 256'h52f8a6f809f96bf9c6f92efa95faf8fa64fbcefb36fca8fc14fd7afdeafd56fe;
    inBuf[2688] = 256'hbcfe2aff92fff5ff5f00c10020018601e20139029902ed023a038f03da031904;
    inBuf[2689] = 256'h5e049b04cf0409053d0564058b05af05cc05e805ff050f0620062c0632063706;
    inBuf[2690] = 256'h3a0636062d06240616060406f105da05bb059d057f0556052d050605d504a404;
    inBuf[2691] = 256'h750440040a04d6039c0361032703e802ad0274023202f201b60173013401f600;
    inBuf[2692] = 256'hb0006f003200edffaeff70ff2bffedfeb0fe6cfe2efef1fdadfd70fd2ffde9fc;
    inBuf[2693] = 256'habfc6cfc27fce8fba4fb60fb25fbe3fa9ffa62fa21fae1f9a8f966f926f9f1f8;
    inBuf[2694] = 256'hb2f873f83ff803f8caf796f756f71df7edf6aff675f648f610f6d9f5abf574f5;
    inBuf[2695] = 256'h42f51bf5e9f4bcf49af46ff44bf430f40ef4f0f3dbf3c2f3b0f3a4f393f38cf3;
    inBuf[2696] = 256'h8bf384f387f391f399f3a9f3baf3caf3e9f30bf426f44ff47cf4a3f4d7f410f5;
    inBuf[2697] = 256'h45f586f5c9f506f652f6a2f6ecf642f79bf7f0f753f8b5f813f97ff9e9f950fa;
    inBuf[2698] = 256'hc3fa34fba1fb17fc8cfcfcfc75fde8fd58fecffe3fffabff1f008b00f4006301;
    inBuf[2699] = 256'hc9012a029402f5024d03ab0302045104a304f00435057b05ba05f00526065a06;
    inBuf[2700] = 256'h8506ac06ce06e706fd0612071f072507290725071a070e07fa06e106c706a506;
    inBuf[2701] = 256'h7c0652062406f005bb057e053d05fd04b80470042a04dd038a033b03ea029302;
    inBuf[2702] = 256'h4002ea018f013801de0081002900ceff6eff16ffb9fe5afe04feaafd4efdfafc;
    inBuf[2703] = 256'ha3fc4afcfdfbaffb5cfb13fbc9fa81fa42fafef9baf982f945f90af9dbf8a7f8;
    inBuf[2704] = 256'h73f849f81af8eff7cff7a8f785f76df74bf72ef71ef706f7f1f6e5f6d2f6c3f6;
    inBuf[2705] = 256'hbdf6b0f6a9f6aaf6a1f6a1f6a9f6a5f6a8f6b4f6b6f6bff6d3f6dff6edf600f7;
    inBuf[2706] = 256'h0ff725f73cf74ef76af785f799f7b9f7d9f7eff711f835f851f876f89ef8bff8;
    inBuf[2707] = 256'heaf815f93cf96cf99df9caf9fff933fa63fa9dfad6fa0bfb4afb86fbc0fb02fc;
    inBuf[2708] = 256'h3efc7bfcc3fc05fd44fd8cfdccfd0dfe5bfea1fee2fe30ff78ffbdff0c005400;
    inBuf[2709] = 256'h9900e6002c016f01bb01010244028c02d002110355039403d10310044b048604;
    inBuf[2710] = 256'hc204f60429055c058a05b805e00504062b064e06670682069c06af06c106d106;
    inBuf[2711] = 256'hdc06e706eb06ec06ed06ea06e506df06d106c106b2069c0683066a064b062b06;
    inBuf[2712] = 256'h0c06e405ba059305650538050d05db04a70475043f040904d5039c0366033303;
    inBuf[2713] = 256'hf902c0028a024f021502e201ac01740141010c01d800a700750046001a00eaff;
    inBuf[2714] = 256'hbfff9cff73ff4bff2aff08ffe9fed2feb6fe9bfe89fe74fe5ffe55fe49fe3dfe;
    inBuf[2715] = 256'h3afe36fe31fe36fe39fe3afe44fe53fe5dfe6dfe7ffe90fea4febbfed3feeefe;
    inBuf[2716] = 256'h09ff23ff45ff65ff82ffa5ffcbffedff14003e0062008900b600df0007013201;
    inBuf[2717] = 256'h5c018a01b701dc010502320259028002ab02d102f7021e03410365038903a903;
    inBuf[2718] = 256'hc903e70301042204400455046e0488049a04b004c504d404e804fb0404051205;
    inBuf[2719] = 256'h1f05260532053d05410548054b054b05500552054f05530553054b054a054805;
    inBuf[2719] = 256'h1f05260532053d05410548054b054b05500552054f05530553054b054a054805;    
    inBuf[2720] = 256'h40053f053b05320530052b0520051e051a05120512050e05060507050205fa04;
    inBuf[2721] = 256'hfc04fa04f404f904f804f104f804f704f104fd040105fb0406050c0509051505;
    inBuf[2722] = 256'h1e051e052d053705380547055505590568057705810593059e05a705bc05c905;
    inBuf[2723] = 256'hd105e605f405fc0510061e062406370644064b065b0665066706760680068306;
    inBuf[2724] = 256'h900697069806a506ac06ac06b606bb06ba06c206c606c406cc06cc06c706d206;
    inBuf[2725] = 256'hd406c906cc06ce06c606c806c706bd06bf06bd06b406b506b306ab06ab06a806;
    inBuf[2726] = 256'ha006a206a0069c06a306a1069906a206a506a006a606a906a906b406b506b206;
    inBuf[2727] = 256'hbd06c206c006cb06d006ce06d806dc06d906e306e906e706ed06f006ed06f306;
    inBuf[2728] = 256'hf106ed06f306f006e906ed06e806dc06d906d306c506bf06b306a10691067f06;
    inBuf[2729] = 256'h6a0656063b0622060b06e705c205a4057c05540531050105d004a70475044204;
    inBuf[2730] = 256'h1404dd03a40372033a030103cd02930256022002e601a8016e013501fb00c200;
    inBuf[2731] = 256'h87004e001700ddffa6ff73ff3eff0cffe0feb2fe85fe5cfe33fe0efef1fdd2fd;
    inBuf[2732] = 256'hb3fd9cfd87fd72fd68fd61fd57fd54fd55fd54fd58fd61fd6dfd80fd94fda5fd;
    inBuf[2733] = 256'hbefddcfdf7fd19fe3ffe61fe8bfeb7fedefe0dff40ff6dff9fffd8ff0e004a00;
    inBuf[2734] = 256'h8600bb00f80039017101b001f3012e026b02aa02e40221035d039003ca030404;
    inBuf[2735] = 256'h330467049b04c704f504220544056d059505b005d005f3050a0623063d064f06;
    inBuf[2736] = 256'h6106730681068f0698069b06a006a406a306a2069e0695068c067f0671066406;
    inBuf[2737] = 256'h51063c0628060d06f105d905ba0598057705520530051005e804c00498046c04;
    inBuf[2738] = 256'h43041e04f203c7039c0369033c031103de02ac027c0246021302df01a6017001;
    inBuf[2739] = 256'h3601f900c100840042000900caff84ff48ff09ffbffe81fe40fef7fdb6fd74fd;
    inBuf[2740] = 256'h2afde7fca1fc5afc19fccefb80fb3ffbf8faabfa69fa1ffad1f98ff944f9f6f8;
    inBuf[2741] = 256'hb4f86af81ff8dff794f74af70df7c6f67ff648f607f6c5f592f558f51ef5f3f4;
    inBuf[2742] = 256'hc1f48ff46bf442f41ef401f4dbf3bff3aff393f37ff377f367f35ff360f356f3;
    inBuf[2743] = 256'h54f360f365f372f387f395f3adf3cbf3e3f309f436f459f488f4bef4edf426f5;
    inBuf[2744] = 256'h66f59ff5e0f527f66cf6b8f604f749f79cf7eff73bf892f8e9f838f992f9ecf9;
    inBuf[2745] = 256'h3dfa98faf2fa42fb9cfbf7fb4afca2fcf9fc49fda0fdf3fd40fe97fee9fe30ff;
    inBuf[2746] = 256'h80ffceff120059009f00dd001e015b018f01c501f80121024c0275029602b802;
    inBuf[2747] = 256'hd602ea02ff0212031b032503300330032e0330032a031e0313030003ec02dc02;
    inBuf[2748] = 256'hc002a10286025f0234021402e801b40187014f011001dc00a00059001a00d2ff;
    inBuf[2749] = 256'h85ff46fff9fea2fe5afe0afeb1fd63fd0efdb2fc64fc0dfcaefb5cfb05fba9fa;
    inBuf[2750] = 256'h58fafcf99df94df9f4f896f847f8ebf78bf73cf7e4f686f637f6e0f588f53df5;
    inBuf[2751] = 256'he9f492f44cf4fcf3aef36ff323f3d8f2a2f261f21ef2eff1b6f17df154f124f1;
    inBuf[2752] = 256'hf8f0d8f0acf088f074f052f036f02cf014f003f0feefefefeaeff1efeaefeeef;
    inBuf[2753] = 256'hffef00f010f02ef039f051f077f08ff0b4f0e4f007f137f170f19df1daf11ef2;
    inBuf[2754] = 256'h55f29af2e2f220f36ff3bff301f456f4adf4f5f44ef5a9f5f5f552f6b2f603f7;
    inBuf[2755] = 256'h64f7c5f717f87cf8e2f838f99cf901fa59fac1fa2afb83fbe7fb4efca9fc0dfd;
    inBuf[2756] = 256'h6ffdc6fd25fe82fed6fe31ff88ffd8ff2f008100c70014015f01a201e9012a02;
    inBuf[2757] = 256'h62029f02d60207033d036e039603c203e9030704280448046004750488049704;
    inBuf[2758] = 256'ha204aa04af04af04a8049f0495048604710458043f041f04fa03d503ad037f03;
    inBuf[2759] = 256'h51031e03e502af0275023402f701b80173013101ea009d0057000c00bbff70ff;
    inBuf[2760] = 256'h1fffc9fe7dfe2bfed3fd83fd2efdd3fc85fc33fcd9fb8bfb39fbe3fa96fa46fa;
    inBuf[2761] = 256'hf5f9aff965f91bf9daf895f853f81bf8def7a9f77cf748f718f7f5f6cdf6a9f6;
    inBuf[2762] = 256'h8ff670f656f64af639f62af625f61df618f61ef623f62cf63af647f65af675f6;
    inBuf[2763] = 256'h90f6b0f6d6f6fbf626f758f78af7bff7f5f72ff871f8b2f8f3f83df984f9ccf9;
    inBuf[2764] = 256'h1dfa6bfab5fa08fb5bfbacfb04fc56fca8fc04fd5afda9fd05fe5ffeb2fe0bff;
    inBuf[2765] = 256'h63ffb9ff13006600ba0016016801b90110026202b20208035503a103f0033604;
    inBuf[2766] = 256'h7f04cb040d054e059405d0050d064a067f06b906f2061c074d078107a907d207;
    inBuf[2767] = 256'hfe0723084c0872088f08b108d308ea0805091f0934094b095d0969097c098909;
    inBuf[2768] = 256'h8d099909a0099f09a309a20999099609910985097c096d095a094c0936091d09;
    inBuf[2769] = 256'h0d09f308d008b9089c0878085b0837080e08ee07c6079807750749071507ee06;
    inBuf[2770] = 256'hc006870658062706ee05ba0582054a051805db049b0468042f04f303c0038603;
    inBuf[2771] = 256'h4a031803e102a9027c0248021102e701bc018d0165013c011301f200ce00ad00;
    inBuf[2772] = 256'h940076005600460033001d0014000900fbfffafffcfff9ff01000c0013002500;
    inBuf[2773] = 256'h3800490067008600a000c700f200140142017601a301db01150247028602ca02;
    inBuf[2774] = 256'h030347038d03c90311045d049c04e80436057605c10512065606a106ef063307;
    inBuf[2775] = 256'h7f07cc070c0855089f08dc08240967099d09e009230a540a8b0ac50af20a220b;
    inBuf[2776] = 256'h4f0b710b9c0bc30bdc0bfd0b1a0c2a0c430c570c5c0c6b0c760c750c7a0c7a0c;
    inBuf[2777] = 256'h730c740c6b0c560c500c400c240c160c020ce10bc90bad0b890b6f0b490b1b0b;
    inBuf[2778] = 256'hfc0ad30aa00a7a0a4f0a1a0af209c4098d0961092f09f608c90895085f083308;
    inBuf[2779] = 256'hff07c8079d076b0737070c07da06a9067f064b061a06f605c605930570054805;
    inBuf[2780] = 256'h1905f304cb04a20480045c0436041604f103ce03b503970374035d0345032703;
    inBuf[2781] = 256'h1103fc02e502d302c002ac029f028e027d0276026c025c025802530247024402;
    inBuf[2782] = 256'h43023a023b023d0239023d02430246024d0255025d026c0277027e029002a102;
    inBuf[2783] = 256'hae02c702de02ed0205032003350352036e038503a403c303dc03000421043904;
    inBuf[2784] = 256'h5f0484049d04bf04e404010528054c0567058e05b205cc05ef0511062a064e06;
    inBuf[2785] = 256'h71068806a606c506da06f4060e07200738074a075507670775077e078c078f07;
    inBuf[2786] = 256'h8e0795079207890787077c076d07650752073c072c071107f406da06b6069106;
    inBuf[2787] = 256'h710646061906f005be058b055b052005e704af046d043004f503ab0364032003;
    inBuf[2788] = 256'hd5028e024802f601a8015d010c01c10072001c00d0ff83ff2dffe1fe94fe3ffe;
    inBuf[2789] = 256'hf3fdabfd5dfd13fdc7fc7afc37fcf3fba9fb6afb2cfbe8faadfa73fa38fa05fa;
    inBuf[2790] = 256'hd2f99cf970f945f917f9f3f8d0f8acf890f875f85cf849f834f823f81cf810f8;
    inBuf[2791] = 256'h06f808f807f808f811f818f821f831f840f854f86ef885f89ef8bcf8dbf8fff8;
    inBuf[2792] = 256'h24f947f970f999f9c0f9f0f921fa4dfa80fab4fae4fa1cfb52fb84fbbcfbf4fb;
    inBuf[2793] = 256'h27fc61fc9cfcd1fc0bfd42fd78fdb3fde8fd17fe4efe82feb2fee8fe18ff41ff;
    inBuf[2794] = 256'h72ff9fffc5fff0ff19003c00600082009e00be00dc00f3000b01230133014201;
    inBuf[2795] = 256'h51015c0166016e016f01730175016e016801650157014a013f012a0115010401;
    inBuf[2796] = 256'he700c900b2009300700051002900ffffdcffb1ff81ff58ff28fff4fec4fe8efe;
    inBuf[2797] = 256'h57fe26feecfdb0fd7dfd40fd00fdc9fc8bfc49fc11fcd0fb8bfb51fb10fbccfa;
    inBuf[2798] = 256'h92fa52fa0dfad0f990f94ff915f9d4f892f85bf81ff8e0f7aaf770f735f702f7;
    inBuf[2799] = 256'hc9f696f66af632f6fef5d8f5a8f57cf55cf531f509f5eef4c9f4a9f495f479f4;
    inBuf[2800] = 256'h5ef44ef439f42bf424f414f40cf40ff409f40af413f414f420f434f43df44ff4;
    inBuf[2801] = 256'h6df481f49af4bcf4dbf402f52ef552f57ff5b3f5def515f651f683f6bff602f7;
    inBuf[2802] = 256'h3ef781f7c9f70bf858f8a5f8e8f838f98af9d1f922fa7bfac9fa1afb6ffbbefb;
    inBuf[2803] = 256'h15fc6bfcb7fc09fd60fdaefd00fe50fe98fee9fe37ff78ffc2ff0c0049008b00;
    inBuf[2804] = 256'hcd0002013c017701a601d80109022e02540279029502b302cc02dc02ef020003;
    inBuf[2805] = 256'h030308030e030b030303f902e902da02c702ab028f0273024b022302ff01d101;
    inBuf[2806] = 256'h9e016e013601fd00c800890046000a00c6ff7fff3cfff1fea4fe60fe15fec3fd;
    inBuf[2807] = 256'h7bfd30fddffc96fc49fcfafbb2fb67fb19fbd4fa8afa40fafcf9b5f971f937f9;
    inBuf[2808] = 256'hf5f8b4f87ff846f80cf8def7adf779f750f726f7fdf6dcf6bdf69ff686f66df6;
    inBuf[2809] = 256'h5af64af638f62df627f61ff61ef622f621f62bf63cf646f654f668f67cf697f6;
    inBuf[2810] = 256'hb6f6d1f6f4f61cf740f76af798f7c5f7f7f729f85af896f8cff805f949f98cf9;
    inBuf[2811] = 256'hc7f90bfa52fa96fae1fa29fb6ffbbdfb0bfc5afcaefcfcfc4afda0fdf1fd43fe;
    inBuf[2812] = 256'h9dfeebfe3cff99ffecff3d009900eb003b019701ea013a029002e10230038503;
    inBuf[2813] = 256'hd3031f046e04b70403054f059105d7051f065c069d06de0614074e078807b707;
    inBuf[2814] = 256'hea071d0844086c089508b608d708f30806091e0931093c094a09520953095709;
    inBuf[2815] = 256'h54094909420935091f090a09f008d408b7089008680843081308de07ae077707;
    inBuf[2816] = 256'h3a07fd06ba0678063606eb05a10557050505b60467040f04b90365030903b102;
    inBuf[2817] = 256'h5d020002a4014a01eb0092003b00dcff82ff2dffd1fe7bfe2afed3fd80fd31fd;
    inBuf[2818] = 256'hdefc94fc4cfcfffbbafb7bfb36fbf8fabffa85fa51fa1efaeaf9c0f99bf974f9;
    inBuf[2819] = 256'h54f939f91df905f9f4f8e6f8daf8d2f8ccf8cbf8cdf8d4f8def8e9f8f9f80df9;
    inBuf[2820] = 256'h23f93df95bf97bf9a0f9c2f9e8f916fa44fa74faa9fadafa0ffb4efb89fbc1fb;
    inBuf[2821] = 256'h03fc42fc81fccafc0cfd4bfd94fddcfd26fe74febafefffe4eff98ffe3ff3200;
    inBuf[2822] = 256'h7a00c20012015b01a501f3013a028102ce0212035803a203e60328046e04ac04;
    inBuf[2823] = 256'heb042f056c05a805e6051b0654068f06bf06f106250752078007ae07d207fa07;
    inBuf[2824] = 256'h2208420864088808a108bd08d908ec080109150923093409400946094f095309;
    inBuf[2825] = 256'h5309590956094e094d09410931092b091b090509f908e208c508b50899087608;
    inBuf[2826] = 256'h5e083d081408f607d007a307800756072707ff06cf069e06740640060b06df05;
    inBuf[2827] = 256'ha905710544050c05d204a2046c0435040304c903950366032b03f302c5028e02;
    inBuf[2828] = 256'h58022b02f701c301980168013a011301e400b60094006a00420024000100dbff;
    inBuf[2829] = 256'hbdff9eff80ff68ff4fff34ff1eff0afff8fee7fed7fecdfec5febafeb2feadfe;
    inBuf[2830] = 256'ha8fea8fea9fea7fea9feaffeb5febbfec4fecffedafee7fef8fe0bff19ff29ff;
    inBuf[2831] = 256'h3eff53ff68ff7fff93ffaaffc4ffddfff7ff11002900440061007c009700b100;
    inBuf[2832] = 256'hce00ed00070121013f015a0173019001aa01c301dd01f601100229023d025502;
    inBuf[2833] = 256'h6e027e029102a802b802c802db02ea02f9020703110320032e0335033f034803;
    inBuf[2834] = 256'h4e0355035d03600363036403640367036603600360035d035603550351034603;
    inBuf[2835] = 256'h41033b0332032903200314030b030003f002e502d902ca02bd02af029f029402;
    inBuf[2836] = 256'h860276026b025c024c0240023202230218020a02fa01ee01e201d501cb01bd01;
    inBuf[2837] = 256'hb301aa019b018e0187017b016f016c01630156014f01470140013d0135012d01;
    inBuf[2838] = 256'h280123011e011b01170113010f01060102010201fd00f700f300f200f200f000;
    inBuf[2839] = 256'hec00e900e800e300de00db00d900d500d100ce00cb00c700c300be00b900b500;
    inBuf[2840] = 256'hb000aa00a4009f009c00990091008a00860081007a0074006b0062005f005900;
    inBuf[2841] = 256'h50004b0045003c0038003200260020001c0013000a0007000000f8fff2ffecff;
    inBuf[2842] = 256'he7ffe3ffddffd4ffcfffcbffc5ffc0ffbaffb5ffb3ffb0ffaaffa7ffa4ffa1ff;
    inBuf[2843] = 256'h9fff9cff98ff96ff93ff90ff8fff8cff88ff87ff86ff84ff83ff80ff7eff7dff;
    inBuf[2844] = 256'h7aff77ff75ff72ff71ff71ff6eff6bff6aff67ff63ff63ff5fff58ff54ff54ff;
    inBuf[2845] = 256'h4fff4aff46ff42ff3dff36ff2fff2cff26ff1eff1cff18ff10ff0bff08ff03ff;
    inBuf[2846] = 256'hfdfef4feedfeecfee5fedafed6fed2fecbfec7fec1febbfeb9feb6feaefea9fe;
    inBuf[2847] = 256'ha6fea1fe9dfe99fe96fe95fe91fe8ffe90fe8bfe85fe85fe86fe87fe86fe83fe;
    inBuf[2848] = 256'h81fe84fe84fe84fe88fe88fe87fe8bfe8dfe8dfe90fe92fe92fe96fe99fe9afe;
    inBuf[2849] = 256'h9cfe9efe9efea1fea2fea1fea4fea5fea5fea6fea8fea7fea7fea8fea7fea5fe;
    inBuf[2850] = 256'ha2fea1fea0fe9bfe96fe94fe8bfe84fe83fe7cfe73fe6efe65fe5afe54fe4afe;
    inBuf[2851] = 256'h3ffe36fe29fe1efe15fe06fef6fdecfddbfdcbfdbffdaefd9cfd8ffd7efd6dfd;
    inBuf[2852] = 256'h60fd4efd3dfd2efd1afd09fdfdfce9fcd6fccafcb8fca5fc97fc86fc72fc63fc;
    inBuf[2853] = 256'h54fc44fc37fc27fc18fc0efcfffbeffbe5fbdbfbcefbc5fbb8fbadfba9fba4fb;
    inBuf[2854] = 256'h9cfb97fb91fb8cfb88fb84fb82fb82fb80fb80fb83fb85fb87fb8bfb8ffb97fb;
    inBuf[2855] = 256'h9efba1fba9fbb4fbbbfbc2fbcdfbdafbe6fbf1fbfbfb0afc1bfc2cfc3cfc4bfc;
    inBuf[2856] = 256'h59fc6cfc80fc91fca5fcbbfccffce3fcf7fc0dfd25fd3dfd52fd69fd7efd94fd;
    inBuf[2857] = 256'hadfdc5fddbfdf1fd0bfe25fe3ffe58fe71fe8cfea6febdfed8fef4fe09ff20ff;
    inBuf[2858] = 256'h3bff54ff6dff86ff9fffb9ffd3ffeaff010019002f004800610077008c00a300;
    inBuf[2859] = 256'hb900ce00e200f6000a011c012e014401580169017b018c019b01ac01ba01c601;
    inBuf[2860] = 256'hd301e101ed01f80100020a0215021d0223022b02320237023c02400243024502;
    inBuf[2861] = 256'h4502430241023e023d023a0234022f022a0222021b0215020c020002f301e601;
    inBuf[2862] = 256'hd801c901b801a8019701840171015e014a0134011f010a01f000d700be00a400;
    inBuf[2863] = 256'h89006e00520035001a00ffffe1ffc2ffa3ff84ff66ff46ff27ff0bffecfecafe;
    inBuf[2864] = 256'haafe8dfe6ffe4ffe2ffe12fef4fdd3fdb6fd9bfd7dfd61fd49fd2dfd10fdf7fc;
    inBuf[2865] = 256'he0fccafcb5fc9efc88fc76fc63fc4ffc3ffc30fc23fc18fc0cfc02fcfbfbf1fb;
    inBuf[2866] = 256'heafbe7fbe3fbe2fbe2fbe0fbe0fbe5fbe7fbecfbf5fbfcfb05fc11fc1cfc2bfc;
    inBuf[2867] = 256'h3cfc4bfc5dfc70fc83fc99fcaefcc2fcdafcf5fc10fd2afd45fd60fd7efd9bfd;
    inBuf[2868] = 256'hbbfddbfdf7fd17fe3cfe5efe7ffea3fec3fee5fe0bff2bff4dff73ff96ffb9ff;
    inBuf[2869] = 256'hdfffffff2000470069008a00ae00d000f10011013001520175019401b301d001;
    inBuf[2870] = 256'heb01080224023e025c0279028f02a802c202d902ef02060319032d033f034e03;
    inBuf[2871] = 256'h600372037f038e039d03a903b603c303cb03d403df03e603ec03f103f503f803;
    inBuf[2872] = 256'hfa03fc03ff03ff03fd03fd03fa03f603f403ed03e303de03d603cb03c103b303;
    inBuf[2873] = 256'ha6039b038d037f036f035b034a033b03260313030403ef02d802c402ad029502;
    inBuf[2874] = 256'h7e026302490234021c020202e701cd01b4019d01820166014c0131011301f600;
    inBuf[2875] = 256'hdd00c700ae0092007900610047002d001400fdffe7ffd0ffb8ffa1ff8bff74ff;
    inBuf[2876] = 256'h5fff4bff39ff2bff1eff0fff01fff2fee3fed7fecdfec1feb7feb1fea9fea1fe;
    inBuf[2877] = 256'h9bfe97fe94fe93fe94fe94fe94fe94fe96fe97fe9bfea3feacfeb5febdfec5fe;
    inBuf[2878] = 256'hcdfed7fee1feecfefafe07ff14ff23ff34ff44ff53ff63ff75ff85ff97ffaaff;
    inBuf[2879] = 256'hbcffceffe2fff5ff07001a002c003e0052006300750088009900ab00bf00d200;
    inBuf[2880] = 256'he500f8000801170129013801460156016401730181018d019801a401b101be01;
    inBuf[2881] = 256'hca01d201d901e401ed01f301fc01030206020b02100216021a021d021e022002;
    inBuf[2882] = 256'h22022202240224022402230222021f021b02150211020f020b0207020402fd01;
    inBuf[2883] = 256'hf601f101eb01e301dc01d501cc01c301ba01b001a801a001990193018c018401;
    inBuf[2884] = 256'h7a016e0163015601490141013a01320127011c01130109010001f800f100e700;
    inBuf[2885] = 256'hdd00d500cc00c300bb00b300ad00a5009d0096008e0086007f00790075006f00;
    inBuf[2886] = 256'h680063005f0059005500540050004d004c004700430042003e003c003d003b00;
    inBuf[2887] = 256'h380038003600370038003600370039003a003c003e003e004100450046004600;
    inBuf[2888] = 256'h4a004d005000530057005d00610066006b006e007200770079007b0080008500;
    inBuf[2889] = 256'h88008c008e00900095009a009d00a300a800ad00b300b600b900c000c400c600;
    inBuf[2890] = 256'hca00cc00cd00d100d500da00e000e300e400e700ea00ed00f000f000f100f400;
    inBuf[2891] = 256'hf400f300f500f700fa00fd00fc00fb00fc00fb00fb00fd00f900f600f700f400;
    inBuf[2892] = 256'hf100f100f000ee00ec00e800e500e500e300df00dc00d900d700d300ce00cb00;
    inBuf[2893] = 256'hc900c500c100be00ba00b600b100ac00a800a3009e009a00950090008d008b00;
    inBuf[2894] = 256'h8800860083007f007c0079007500730070006e006b0068006400640064006300;
    inBuf[2895] = 256'h6100610060005e005b005a005b005a0058005800590058005a005d005c005b00;
    inBuf[2896] = 256'h5c005e0062006500660067006800670069006c006d0070007300750077007600;
    inBuf[2897] = 256'h75007700780077007800790079007b007b007a007b007c007a00790078007600;
    inBuf[2898] = 256'h7400730070006e006d006a00670062005d00580053004d004a00480043003c00;
    inBuf[2899] = 256'h35002d00270022001a0014000c000300fbfff2ffe7ffe0ffd9ffcfffc5ffbbff;
    inBuf[2900] = 256'hb0ffa5ff9bff93ff8dff83ff77ff6fff69ff60ff57ff4dff45ff3dff36ff2dff;
    inBuf[2901] = 256'h23ff1aff13ff0bff04fffdfef8fef1fee9fee4fee0fedefedbfed8fed4fed0fe;
    inBuf[2902] = 256'hcbfec7fec4fec3fec1fec2fec3fec2fec3fec4fec4fec5fec6fec7fec8fecbfe;
    inBuf[2903] = 256'hcbfecefed3fed7fedcfee2fee7feebfef0fef4fefbfe03ff09ff10ff18ff1fff;
    inBuf[2904] = 256'h27ff2eff34ff3dff46ff4eff58ff61ff66ff6dff75ff7dff85ff8cff92ff9bff;
    inBuf[2905] = 256'ha3ffaaffb4ffbdffc5ffceffd9ffe2ffedfff6fffbff020008000d0013001a00;
    inBuf[2906] = 256'h21002a00310036003c00410047004c0050005300570059005c00620067006b00;
    inBuf[2907] = 256'h6d006e006f00710072007400770077007800790077007500750072006e006d00;
    inBuf[2908] = 256'h6900660064005f005d005b0054004d004800400039003200280021001c001400;
    inBuf[2909] = 256'h0d000500f9ffefffe6ffdcffd3ffcbffbfffb4ffa9ff9bff8fff85ff77ff6bff;
    inBuf[2910] = 256'h61ff55ff4aff3eff30ff23ff15ff08fffdfef0fee1fed6fecbfebcfeb1fea7fe;
    inBuf[2911] = 256'h9cfe91fe85fe78fe6efe63fe58fe51fe48fe3dfe37fe2ffe25fe1ffe17fe0ffe;
    inBuf[2912] = 256'h0afe05fe00fefbfdf5fdeffdeefdeafde5fde3fde2fde3fde6fde8fdeafdedfd;
    inBuf[2913] = 256'hedfdecfdf0fdf3fdf7fdfefd02fe07fe10fe16fe1bfe24fe29fe2ffe3bfe44fe;
    inBuf[2914] = 256'h4bfe55fe5ffe6afe75fe7dfe85fe91fe9afea1feadfeb7fec0fecbfed8fee8fe;
    inBuf[2915] = 256'hf8fe02ff0cff18ff20ff28ff32ff3aff43ff50ff5bff66ff72ff7bff82ff89ff;
    inBuf[2916] = 256'h90ff99ffa2ffa8ffafffb8ffbdffc1ffc6ffcbffd0ffd6ffd9ffddffe3ffe7ff;
    inBuf[2917] = 256'hebffeeffeffff0fff3fff3fff3fff4fff4fff4fff5fff4fff3fff2ffefffebff;
    inBuf[2918] = 256'he8ffe5ffe1ffdfffdbffd5ffd1ffccffc4ffbeffbaffb5ffb1ffafffaaffa6ff;
    inBuf[2919] = 256'ha3ff9fff99ff93ff8dff86ff7fff78ff72ff6dff65ff5eff58ff51ff49ff40ff;
    inBuf[2920] = 256'h37ff31ff2bff24ff1eff17ff0fff09ff03fffdfef7fef0fee9fee3feddfed7fe;
    inBuf[2921] = 256'hd4fed0fecbfec8fec6fec2febffeb9feb4feb1feaefeaafea7fea3fe9ffe9efe;
    inBuf[2922] = 256'h9cfe9afe9cfe9bfe9bfe9cfe9cfe9efea0fe9ffea0fea4fea4fea5feaafeadfe;
    inBuf[2923] = 256'hb0feb5febafebffec7feccfed3fedbfee1fee7feedfef2fef9fe02ff08ff0fff;
    inBuf[2924] = 256'h18ff20ff2aff34ff3dff47ff51ff58ff60ff68ff71ff7bff85ff8fff9bffa7ff;
    inBuf[2925] = 256'hb1ffbcffc7ffd1ffddffe8fff3ffffff09000f00180023002b0034003c004400;
    inBuf[2926] = 256'h4d0056005f006900710078007f0085008b0094009a009f00a500ac00b300bc00;
    inBuf[2927] = 256'hc100c600cd00d200d600db00de00e000e500e700e900eb00eb00ec00ee00ee00;
    inBuf[2928] = 256'hef00f100f100f300f500f500f300f200ee00ed00ec00ea00ea00e900e500e400;
    inBuf[2929] = 256'he300e000df00db00d500d200d000cb00c500c100bb00b700b300ad00a800a400;
    inBuf[2930] = 256'h9e009a00960090008d00890082007c0076006e0069006600620061005e005800;
    inBuf[2931] = 256'h5600520049004400420040003e003d003a00390037003400340032002d002900;
    inBuf[2932] = 256'h260022002100220020001f00200021002400260027002c003000310035003800;
    inBuf[2933] = 256'h39003d004100430048004d0053005d0066006c0074007b007e0084008a008e00;
    inBuf[2934] = 256'h95009e00a500af00b800bd00c400cd00d600e300f000fb00070112011b012601;
    inBuf[2935] = 256'h30013801400146014d0159016601720181018e019801a301aa01af01b601bd01;
    inBuf[2936] = 256'hc101c901d501e001ee01fa01050212021c0223022c0234023b0244024c025002;
    inBuf[2937] = 256'h55025a025e0264026b027402820290029a02a602ad02ac02ad02ab02a802a802;
    inBuf[2938] = 256'hab02ab02af02b302b702be02c502c902d102d402d102d102d102ce02ce02cd02;
    inBuf[2939] = 256'hcb02cc02ca02c502c602c902c902cc02cc02c702c302bc02b002a7029e029302;
    inBuf[2940] = 256'h8b0283027c027b02770270026b0264025b0255024c02400237022c0220021702;
    inBuf[2941] = 256'h0b02fd01f101e601dc01d601cf01c601c101b701a9019c018b01750160014a01;
    inBuf[2942] = 256'h36012a011f0118011801160110010901fc00eb00dd00cc00bb00ad009f009500;
    inBuf[2943] = 256'h8f00870081007e0078007300730070006a0064005b00520049003d0032002a00;
    inBuf[2944] = 256'h21001b001b001a001d0025002a002d002e002c002a0029002600260029002900;
    inBuf[2945] = 256'h2b002f00300035003b003f0045004e0054005a005d005e00610060005b005800;
    inBuf[2946] = 256'h59005c0063006b0071007a00830089009000950095009600960096009c00a100;
    inBuf[2947] = 256'ha400ab00b100b500b900bc00c000c600c900c900c900c500be00ba00b400ad00;
    inBuf[2948] = 256'hab00ab00ac00b000b300b500b600b100aa00a700a2009c009b009a009a009e00;
    inBuf[2949] = 256'h9e009900920087007d0077006f006b006e006c00670065005f00580050004100;
    inBuf[2950] = 256'h330027001a0011000e000900070007000200fcfffafff4ffefffecffe8ffe3ff;
    inBuf[2951] = 256'hdcffcfffc1ffb5ffa8ff9fff9eff9effa1ffa6ffa5ffa2ff9dff91ff81ff72ff;
    inBuf[2952] = 256'h62ff56ff4eff45ff41ff41ff3eff3bff38ff32ff2eff2dff2aff29ff2cff2cff;
    inBuf[2953] = 256'h2aff25ff18ff0cff01fff3fee9fee7fee8feebfef2fef6fef8fefafef6feeefe;
    inBuf[2954] = 256'he4fed5fec7febcfeb1feabfeacfeaffeb4febffec7fecefed3fed5fed9fedbfe;
    inBuf[2955] = 256'hd4fecbfec0feaffea0fe99fe97fe9bfea7feb3fec1fecefed2fed2fecdfec1fe;
    inBuf[2956] = 256'hb3fea7fe98fe8cfe87fe85fe87fe90fe98fea0feabfeb2feb8febbfeb5feaefe;
    inBuf[2957] = 256'ha9fe9efe92fe89fe7cfe74fe70fe6bfe6cfe76fe7ffe88fe90fe8ffe89fe7efe;
    inBuf[2958] = 256'h68fe51fe3bfe23fe10fe06fe03fe08fe15fe1ffe29fe31fe31fe31fe2efe24fe;
    inBuf[2959] = 256'h18fe0afef2fdd8fdc2fdb1fdabfdb1fdbbfdc9fdd7fddbfddbfdd6fdc5fdb0fd;
    inBuf[2960] = 256'h99fd7efd6afd5efd57fd5afd64fd71fd82fd90fd95fd99fd9cfd96fd8ffd88fd;
    inBuf[2961] = 256'h7dfd76fd72fd70fd75fd7dfd83fd8bfd90fd92fd99fda0fda5fdadfdb6fdbbfd;
    inBuf[2962] = 256'hbffdbefdbbfdbcfdbefdc1fdccfddbfdecfd05fe1dfe34fe4bfe5ffe6cfe76fe;
    inBuf[2963] = 256'h79fe78fe77fe77fe7afe87fe99feb1fecefeebfe04ff1dff2fff3cff47ff4fff;
    inBuf[2964] = 256'h54ff57ff58ff5dff68ff76ff8affa8ffcaffecff0c00240035003f0040003e00;
    inBuf[2965] = 256'h3d0040004b005f0078009900be00da00ec00f600f700f000e400d800d400d700;
    inBuf[2966] = 256'he200f5000f0128013f0153015e016401650163015d0157015201520156015d01;
    inBuf[2967] = 256'h6b017d018d019a01a201a1019a018e017f01700161015301480141013c013d01;
    inBuf[2968] = 256'h3f013f0141014301430142013e0136012e0124011a0111010701fa00ec00dd00;
    inBuf[2969] = 256'hcf00c600c200c100c400c900cb00c700ba00a20082005b0033001200fdfff5ff;
    inBuf[2970] = 256'h0000170030004600550058004e0038001600efffc5ff9dff7fff6fff70ff86ff;
    inBuf[2971] = 256'haaffd2fff8ff13001a000c00ecffc0ff90ff60ff35ff1bff14ff1cff35ff5dff;
    inBuf[2972] = 256'h87ffafffccffd7ffd1ffbeffa1ff83ff69ff57ff53ff5bff6cff88ffa8ffc3ff;
    inBuf[2973] = 256'hdaffecfff6fffdfffffffdfffdfffdfff8ffefffe4ffd6ffd0ffd3ffdefff7ff;
    inBuf[2974] = 256'h1a0042006f009b00be00d900e600e300d600c200aa009b0096009c00b600df00;
    inBuf[2975] = 256'h0f0146017e01af01d501e601dc01c00194015f0134011b01170132016901b101;
    inBuf[2976] = 256'h050255029102b302b40297026b0236020402e701de01e7010502320265029a02;
    inBuf[2977] = 256'hc402de02e902e102c802a7027c024d0228020f0203020c0226024b0274029502;
    inBuf[2978] = 256'ha902af02a20282025c0232020b02f301e701e501ed01f601f901f501e901da01;
    inBuf[2979] = 256'hcd01c101b801b801b701ad01980172013c01ff00c3009500800083009c00c200;
    inBuf[2980] = 256'hec000c0117010101cc0083003000e4ffb2ffa1ffb0ffd6ff03002b0045004600;
    inBuf[2981] = 256'h2e000100c6ff87ff4dff1dfffcfeedfeedfef7fe06ff17ff24ff2aff28ff1dff;
    inBuf[2982] = 256'h08ffeafec3fe9bfe78fe63fe63fe7cfea4fed2fef9fe0fff0affebfeb8fe7dfe;
    inBuf[2983] = 256'h44fe15fef9fdf4fd04fe26fe54fe80fe9dfeaafea3fe8bfe68fe43fe23fe10fe;
    inBuf[2984] = 256'h0afe13fe28fe40fe55fe69fe77fe7ffe86fe8afe8afe89fe85fe82fe81fe80fe;
    inBuf[2985] = 256'h80fe83fe83fe80fe7ffe7ffe80fe87fe90fe9dfeadfebbfec4fec6fec1feb4fe;
    inBuf[2986] = 256'ha4fe91fe80fe77fe73fe79fe94fec3fe02ff4bff90ffc4ffddffcfff99ff40ff;
    inBuf[2987] = 256'hd1fe62fe0afedafde1fd23fe94fe1bff9fff02002d001300b9ff34ff9dfe13fe;
    inBuf[2988] = 256'hb3fd92fdb3fd0ffe96fe2cffb6ff1d0050004800070096ff09ff77fef5fd97fd;
    inBuf[2989] = 256'h6bfd73fdadfd11fe8bfe03ff62ff95ff91ff54ffecfe6dfef2fd93fd63fd6bfd;
    inBuf[2990] = 256'ha2fdf4fd4bfe94febefec5feadfe82fe51fe27fe0cfe02fe07fe0efe0dfef6fd;
    inBuf[2991] = 256'hc8fd8efd59fd38fd3dfd6cfdbdfd1ffe7cfebdfed4feb8fe6cfefdfd81fd10fd;
    inBuf[2992] = 256'hc2fca6fcbdfc04fd71fdeefd6cfed9fe25ff44ff30ffe6fe71fedffd47fdc8fc;
    inBuf[2993] = 256'h7efc7bfcc9fc60fd23fef1fe9fff04000900acff01ff32fe6bfdd9fca2fcd1fc;
    inBuf[2994] = 256'h58fd1afef2feb1ff35006a004b00ebff66ffd8fe63fe1afe06fe2bfe7bfee3fe;
    inBuf[2995] = 256'h51ffb4fff9ff18001200ecffb3ff77ff45ff2fff39ff60ffa1fff0ff3b007600;
    inBuf[2996] = 256'h9700960078004000fcffbfff9cffa0ffd7ff3a00b80035018d01a50172010101;
    inBuf[2997] = 256'h6c00dbff75ff56ff89ff0700b50070010d0267026a0213027801be0013009dff;
    inBuf[2998] = 256'h7affafff2d00d2007901fe0148024f021b02bf015301eb009a006e0069008a00;
    inBuf[2999] = 256'hcb001f017201b501d901d301a4015701fd00a9006d0056006d00ad0005016701;
    inBuf[3000] = 256'hc101ff011402fb01b2014901d8007c004f006000ad002901b5012d0277027d02;
    inBuf[3001] = 256'h3502ab01fb004500b3ff69ff79ffe6ff990067012302a502d202af024f02cb01;
    inBuf[3002] = 256'h4501d6008700610063008600c6001c017f01e9014c029502b802a6025402ca01;
    inBuf[3003] = 256'h1a015f00c7ff79ff8fff1200ea00e801d7027f03b5037503d002f3011f018900;
    inBuf[3004] = 256'h50007e00fc009c0131029702bb02a6026b022102e901d001d501f4011b023302;
    inBuf[3005] = 256'h31020d02cc0184014e0141016f01d4015a02e9025d03970392035303eb027a02;
    inBuf[3006] = 256'h1a02d901c001c701e401160255029c02ef0249039c03dc03f503d5037603e102;
    inBuf[3007] = 256'h2a027801f300c000f9009b018c02a203a5045c05a3057005cb04dd03dc02fd01;
    inBuf[3008] = 256'h70015201a3014d022803ff03a704ff04fb04a60418046c03c5024202f401e701;
    inBuf[3009] = 256'h1c0284020e03a10321048004b504c004ab0483044c041004ce0383033103e702;
    inBuf[3010] = 256'hb702b302e5023f03b0031704510451041c04c1035c030703cc02b102b402ce02;
    inBuf[3011] = 256'hff0244039503ed033d047204840472043904e90391033a03ec02ab0277025902;
    inBuf[3012] = 256'h59027602b402080355038803930372033603f302b6028c02790276028402a502;
    inBuf[3013] = 256'hd20208033a0354034b032103db028f0253022a0217020f020102e901c5019e01;
    inBuf[3014] = 256'h87018f01ba01020254029102a8028e024402dd0172011501da00c900dd001501;
    inBuf[3015] = 256'h6101b101fc01330245023202fa01a1013301bd004900e5ff9dff7fff9dfffeff;
    inBuf[3016] = 256'h98005301040278028a022a026401630065ffa7fe59fe87fe23ff09000101d101;
    inBuf[3017] = 256'h5002610200024401550064ffa1fe2efe1afe5dfeddfe7bff18009d00f9002901;
    inBuf[3018] = 256'h2801f6009600100076ffe0fe6cfe33fe49feaefe52ff1600d00053017f014301;
    inBuf[3019] = 256'ha700c8ffd7fe07fe87fd75fdd4fd8cfe6fff4500dd001201dd00510097ffe8fe;
    inBuf[3020] = 256'h76fe63feb6fe57ff1600b6000301e100560089ffb3fe13fed1fdf8fd72fe12ff;
    inBuf[3021] = 256'ha6ff07001f00f5ffa5ff4cff09ffeffe04ff3dff8cffdfff2300510062005500;
    inBuf[3022] = 256'h3000f8ffb8ff77ff33ffebfea0fe58fe1ffe06fe1efe6cfee3fe69ffdcff2100;
    inBuf[3023] = 256'h2400e8ff7fff00ff89fe35fe18fe3cfea4fe47ff0c00ca004e016501ef00eeff;
    inBuf[3024] = 256'h8bfe18fdeffb59fb7bfb40fc6afda5fe9fff200019009effddfe10fe6dfd16fd;
    inBuf[3025] = 256'h19fd6afde8fd71fee5fe2bff40ff29ffeefe9efe42feddfd71fd03fd95fc33fc;
    inBuf[3026] = 256'hf0fbdefb0efc7dfc11fda8fd1afe46fe27fed0fd5ffdfbfcbffcb4fcd5fc10fd;
    inBuf[3027] = 256'h4bfd78fd8afd78fd4afd0dfdc7fc8dfc6bfc65fc80fcb3fceafc13fd14fddafc;
    inBuf[3028] = 256'h6cfce2fb5afb02fbf8fa3efbcbfb81fc36fdc9fd1dfe1ffed8fd54fdacfc06fc;
    inBuf[3029] = 256'h80fb27fb0dfb32fb8afb0ffcaefc48fdc6fd08fef0fd79fdacfca7fba4fadbf9;
    inBuf[3030] = 256'h74f990f92bfa21fb44fc57fd21fe83fe6efee8fd17fd28fc4bfbb7fa8bfac7fa;
    inBuf[3031] = 256'h5ffb25fce0fc6bfdacfd9bfd4efddafc4dfcbefb38fbc1fa6efa4cfa5efaacfa;
    inBuf[3032] = 256'h28fbb6fb40fcaffceffc07fd03fdecfcd5fcc1fca8fc8afc63fc2cfcf1fbb9fb;
    inBuf[3033] = 256'h81fb51fb2afb0dfb08fb25fb62fbbcfb1dfc68fc8ffc88fc4cfcecfb77fbfdfa;
    inBuf[3034] = 256'h9bfa6bfa7efae3fa90fb61fc2cfdb7fdd3fd72fd9efc7cfb51fa60f9d9f8dbf8;
    inBuf[3035] = 256'h5af92bfa1cfbf8fb93fce2fce6fcaafc46fcc9fb3cfbb3fa3bfadff9b0f9b6f9;
    inBuf[3036] = 256'hedf950fac8fa35fb84fba0fb7efb2afbb8fa3bfad2f98ef974f98bf9cff92efa;
    inBuf[3037] = 256'h9cfa08fb5afb8bfb94fb71fb2efbd7fa71fa11fac7f999f991f9a7f9c5f9ddf9;
    inBuf[3038] = 256'he5f9d5f9c1f9bdf9d9f923fa8efafefa56fb79fb52fbeefa6dfaf6f9b9f9cdf9;
    inBuf[3039] = 256'h28faaffa31fb7cfb7bfb2ffbacfa25fac7f9aff9eff97cfa2efbdafb53fc75fc;
    inBuf[3040] = 256'h44fcd4fb45fbc6fa73fa56fa73fabefa24fb98fb07fc5bfc8bfc94fc7bfc5afc;
    inBuf[3041] = 256'h45fc45fc5ffc85fc9ffca8fc9ffc91fc97fcbefc04fd5efdb0fde1fde4fdbafd;
    inBuf[3042] = 256'h6cfd13fdc0fc7efc58fc4dfc5afc86fccffc32fdacfd30feaffe26ff8effe8ff;
    inBuf[3043] = 256'h31005a004e0001006effa8fedffd47fd0ffd4ffdf6fdd8feb6ff51007e003100;
    inBuf[3044] = 256'h7bff89fe9cfdeefcb2fc01fdd0fdf9fe430072015502d302e202920201024a01;
    inBuf[3045] = 256'h8b00e0ff59ff04ffe6fefafe38ff91ffebff3500610066004e002400f5ffd0ff;
    inBuf[3046] = 256'hbeffc0ffdaff0b004d00a10000015e01b8010402350244022b02e70189012b01;
    inBuf[3047] = 256'he900da00fb002d014a012801b500080055ffd9fed4fe5cff5c009e01c8028103;
    inBuf[3048] = 256'h9303f302cb017a0069ffeffe3eff4200b2012f035004cc049404c20392025b01;
    inBuf[3049] = 256'h6100cfffb7ff04008f003701d0013f027e028a026a023802ff01ca01a5018c01;
    inBuf[3050] = 256'h7a017d019b01dc015002e9028c0322048904a80487042b04a4030b036c02d301;
    inBuf[3051] = 256'h5e011c011e0178011c02e802b5034b047f045704e903670318031f037e032104;
    inBuf[3052] = 256'hcd04480580056b051f05cc048d0472048904bb04e9040505f204a9044704e203;
    inBuf[3053] = 256'h9c03a003ed0373041e05be053106780691068d068f069a06a906b906b1068506;
    inBuf[3054] = 256'h49060906dc05e1050c0645067f069d06940680066a06620679069c06b306be06;
    inBuf[3055] = 256'had068306650660068906f906a10761082209a909cb098309ce08ce07c606e205;
    inBuf[3056] = 256'h48051e055805e105ae0692076708190979096c0900093f0858079c063c065c06;
    inBuf[3057] = 256'h0b0715083409300ac00ac20a430a51091808e706f30571058e0534062d073d08;
    inBuf[3058] = 256'h090959093709b6080d08850732071b073f077807b207f60739088508ef086509;
    inBuf[3059] = 256'hd709390a600a300ab609f3080908330783060d06df05df05fe0541069206ec06;
    inBuf[3060] = 256'h5b07c60723087d08c108ea080509f908bc085908ca072a07b2068006b4066407;
    inBuf[3061] = 256'h600868093b0a880a2b0a3909cc0724068f04390355022102ae02ff03fb053008;
    inBuf[3062] = 256'h190a410b450b2a0a5b086006d30427045c04350552063907a807a8075107e106;
    inBuf[3063] = 256'h9c06850690069f067606f3051e050404da02f3018101b10197020404b0054e07;
    inBuf[3064] = 256'h7c080309db080e08d006710523041d038c026e02ba025c031c04cc044c057505;
    inBuf[3065] = 256'h3e05b904f30313034c02b40163016801a60108028102f6026803e3035d04d004;
    inBuf[3066] = 256'h2b0544050605730494039a02c6013f011f016101d101360267024102d0013c01;
    inBuf[3067] = 256'ha70037000600090037008800e2003e019801e1011a0248026502780284027702;
    inBuf[3068] = 256'h4a02f7017301d00027008fff25fffcfe08ff39ff75ff9affa0ff8eff6fff5aff;
    inBuf[3069] = 256'h5eff6eff7fff86ff76ff61ff61ff88ffe2ff6300e10039014701f600540079ff;
    inBuf[3070] = 256'h87feaefd13fdcffceffc67fd12fec4fe4cff84ff66fffdfe62fec1fd39fde4fc;
    inBuf[3071] = 256'hdbfc27fdbffd94fe7aff3d00b400be005c00adffd4fef7fd38fd9bfc21fcccfb;
    inBuf[3072] = 256'h93fb79fb86fbbdfb22fcbdfc7dfd49fef8fe4eff1dff5afe1cfdb3fb92fa1afa;
    inBuf[3073] = 256'h83fac8fb88fd47ff8a00f300750046ffb7fd2afcecfa16fab1f9b2f9faf977fa;
    inBuf[3074] = 256'h19fbb7fb34fc7afc6ffc25fcc4fb6bfb41fb58fb95fbe1fb21fc39fc30fc1efc;
    inBuf[3075] = 256'h0efc1cfc56fca9fc04fd49fd40fdccfce9fb9dfa2af9e7f713f7ecf680f79af8;
    inBuf[3076] = 256'hfcf959fb5afcdafcd7fc5cfca9fb09fba5faa5fafcfa61fb94fb66fbbdfad8f9;
    inBuf[3077] = 256'h16f9c2f818f911fa49fb59fcdefc8dfc76fbe3f927f8b5f6e5f5cbf577f6cff7;
    inBuf[3078] = 256'h86f95afbf9fcfcfd32fe93fd37fc87fa00f9f6f7a9f714f8e4f8cbf97ffabffa;
    inBuf[3079] = 256'h94fa1bfa66f9aef81ef8c7f7d5f757f828f922fa02fb6dfb4bfbacfab7f9d5f8;
    inBuf[3080] = 256'h63f87df82bf936fa2dfbc6fbd2fb3ffb56fa71f9c9f897f8d4f832f975f96df9;
    inBuf[3081] = 256'hf6f83ff894f729f73cf7d9f7c5f8cdf9affa1efb16fbabfaf6f93ef9bbf877f8;
    inBuf[3082] = 256'h85f8daf846f9c0f93cfa99fad7faeffabdfa48faa2f9daf82ef8d0f7cbf729f8;
    inBuf[3083] = 256'hcaf865f9cff9e3f986f9ebf853f8f6f727f8fff844fab1fbd8fc3efdcafc9efb;
    inBuf[3084] = 256'h00fa79f873f709f73bf7d4f77cf80af96df994f99ef9a3f99df9aaf9d6f90dfa;
    inBuf[3085] = 256'h59faabfad0fac0fa7bfafdf982f949f96ff918fa38fb84fcb6fd76fe6bfe87fd;
    inBuf[3086] = 256'he5fbbff993f7d2f5c3f4a4f475f5f1f6d6f8c6fa56fc55fda7fd4ffd9bfce5fb;
    inBuf[3087] = 256'h66fb62fbe0fb9efc62fde1fdd6fd44fd4bfc1efb18fa79f952f9a8f942fac3fa;
    inBuf[3088] = 256'hfbfaccfa2ffa6af9c3f85af859f8c9f88ff9b1fa2efce2fda3ff260104020502;
    inBuf[3089] = 256'h27019affd4fd46fc37fbcffaf0fa58fbdbfb52fc9cfcbcfcaefc62fce8fb4efb;
    inBuf[3090] = 256'ha9fa2ffa01fa22fa94fa41fb00fcccfcabfd9efea9ffaa005f018e010301beff;
    inBuf[3091] = 256'h1cfe8bfc76fb3bfbdbfbf8fc27fef7fe12ff7ffe7efd6bfcacfb7ffbeafbd4fc;
    inBuf[3092] = 256'hf8fd03ffc8ff2c002b00f2ffb1ff85ff83ffa4ffc8ffd1ffa6ff3fffb1fe0ffe;
    inBuf[3093] = 256'h71fdf6fcacfc9bfccdfc31fda7fd13fe4efe48fe14feccfd96fd94fdbbfdf7fd;
    inBuf[3094] = 256'h45fe99fefcfe93ff6a0060014802e202f20263024501ceff41fecdfca1fbe3fa;
    inBuf[3095] = 256'h9efaddfaaffbfffc96fe340085013f024402a00191006eff84fe0efe23fea9fe;
    inBuf[3096] = 256'h6eff3500c200f000bb0039009eff21ffe0fedcfef3feeffeaafe16fe4bfd95fc;
    inBuf[3097] = 256'h37fc5efc26fd72fef1ff5b01730201030503a602100284012e010e011e014501;
    inBuf[3098] = 256'h50012e01e90081000700a3ff6dff6dffa9ff2400ca007001f10137022702b801;
    inBuf[3099] = 256'h0f015100a4ff46ff5affe5ffd700f401e80274036c03d102e501f80048000b00;
    inBuf[3100] = 256'h3a00a3001901690171014101f100a2009600f600cf011c03a4040906ff063e07;
    inBuf[3101] = 256'hb20699053e04f2021102b901d0014602f502b10373042805ab05e905bf050e05;
    inBuf[3102] = 256'hee038c0226011a009aff9eff1100bf006c010d02b6028703a104f20549076308;
    inBuf[3103] = 256'hef08cf081a08e8067c0537043e03ad02b2022b03da03a8046205db052b065706;
    inBuf[3104] = 256'h5c064a0609068105dc044004d003cf033f04e30494053106ac062707ba075e08;
    inBuf[3105] = 256'hf2082109b508c70786063f055904df039b036003fc026502e201b8011202f902;
    inBuf[3106] = 256'h23043205f10536061b06fd05110672062d07ff079308ca088808e5074e071007;
    inBuf[3107] = 256'h51071b081e09ed09390abc097e08d206fb04560354020c026f027503c504f905;
    inBuf[3108] = 256'he9066b078307740755072e07240722070a07f906ea06ba066406d20500052604;
    inBuf[3109] = 256'h87036603f20300053e065c07fb070408af072c07c106ba061f07e8070609330a;
    inBuf[3110] = 256'h340bea0b160cac0bde0ac30991089c07ee06820659063506e2056305a404c503;
    inBuf[3111] = 256'h280307039003e804c006a008340a210b480bf10a5e0ac90966092309da088408;
    inBuf[3112] = 256'h0b086d07c4060a065005c50477047b04ef04b405a406a6077f080f0955093709;
    inBuf[3113] = 256'hc7084b08f007f8079c08b409f40a140cbe0cdd0ca70c430cd10b5c0bac0a9709;
    inBuf[3114] = 256'h200853067c04fc02f3017801920100029e026d03520446055b06620723088508;
    inBuf[3115] = 256'h6708e7076707310787078508d109fa0ab30bb20bf50ad509aa08c50760076707;
    inBuf[3116] = 256'h9507a007370749060b05dd0337036d0375041206c507f608660921094e085607;
    inBuf[3117] = 256'h99062506000614061c06fd05b3052105530474039a02fa01d6012702d102a803;
    inBuf[3118] = 256'h4d047e043c04a7030a03c4020103c803f6043a064f07100863085b082708eb07;
    inBuf[3119] = 256'hca07d007dc07cd076f078e062f056803590156ffc1fde5fc13fd70febf008c03;
    inBuf[3120] = 256'h350601087f08a707cc05890384013700d2ff1b00a800190116018100aeff11ff;
    inBuf[3121] = 256'h11ff0600d001d2035505b3059004350258ffc1fc18fb9dfa30fb99fca3fe1801;
    inBuf[3122] = 256'hd3038a06b608d809a5092e08ea0584038e015100b6ff7fff6eff5aff46ff4bff;
    inBuf[3123] = 256'h6cffabff020049006f006b0014005fff75fe74fd9afc27fc0dfc19fc2dfc27fc;
    inBuf[3124] = 256'h0bfc26fcabfc92fdaffea1ff0200a6ff9dfe3afdf8fb3bfb49fb29fc91fd17ff;
    inBuf[3125] = 256'h4b00d300b0002f00afff8effebff7d00e800dd002e0005ffc7fdb9fc03fc9afb;
    inBuf[3126] = 256'h43fbe2fa7afa12fad1f9c5f9bbf988f91af968f8bcf77ef7ecf722f9f7faf0fc;
    inBuf[3127] = 256'h99fe94ffa0ffdafe8bfdebfb59fa2cf982f87cf815f9faf9e0fa7dfb7afbd4fa;
    inBuf[3128] = 256'hc9f99ff8c6f7a0f731f859f9b8faaffbcafbecfa43f966f713f6c3f59bf658f8;
    inBuf[3129] = 256'h60fa2efc55fda3fd43fd68fc4dfb5afab9f946f9f1f885f8aff79ef6bbf557f5;
    inBuf[3130] = 256'hb1f58bf618f7bbf63af5dbf29ef07aefbaef2cf117f391f458f5caf571f6eef7;
    inBuf[3131] = 256'h79fa98fd900098020903bb01ecfe20fb3cf705f4e3f100f104f146f166f152f1;
    inBuf[3132] = 256'h31f17bf15ef297f3d6f4a1f594f5ebf405f413f34ef2a3f1b5f084ef56ee8eed;
    inBuf[3133] = 256'hcbed70ef4cf2daf527f92cfb72fbfff95df7a0f49df299f199f132f2cff264f3;
    inBuf[3134] = 256'h1bf411f57bf61ff853f9aff90cf991f7f2f5c4f410f4a6f3f3f24ef1caee04ec;
    inBuf[3135] = 256'hc1e9eae8dfe916eca9eea5f06bf127f181f03df0f2f085f245f47ef593f566f4;
    inBuf[3136] = 256'ha9f233f1b3f09af184f373f595f644f668f4e3f1b9ef97eeebee55f0cef1b0f2;
    inBuf[3137] = 256'hbff217f25ff122f16bf113f2c5f234f390f327f413f559f696f72af8d6f7a9f6;
    inBuf[3138] = 256'hf0f450f34bf20af28ff284f350f489f4def354f28ef040efe7eeb5ef0cf1c9f1;
    inBuf[3139] = 256'h3cf14defadece3ea33ebd1edfdf127f6abf8d7f806f74af4fbf1dcf0e7f0bef1;
    inBuf[3140] = 256'hc3f297f385f4e5f5d3f73afa7cfcbdfd90fde6fb30f975f679f46df333f329f3;
    inBuf[3141] = 256'h8bf256f108f04cefdfefe6f1abf441f7d0f8f0f8fbf7a8f694f528f558f5c2f5;
    inBuf[3142] = 256'h24f655f645f61ff607f607f63cf6b3f658f7fef746f8e4f7d0f618f515f36bf1;
    inBuf[3143] = 256'h78f05af02cf1b3f298f4c6f60ef91ffbd3fceffd36fec8fde0fcabfb61fa02f9;
    inBuf[3144] = 256'h5af775f597f334f2f8f145f3e4f528f91dfceffd74fe14fe7bfd4ffdbffd7bfe;
    inBuf[3145] = 256'hfefec8fea8fddafbb4f982f79af53af48cf3bcf3bbf423f65ff7d6f743f7ecf5;
    inBuf[3146] = 256'h72f48af3aaf3b6f428f68df7b3f8c6f93cfb63fd1c00e40209051b063006b205;
    inBuf[3147] = 256'h2805e004b8044a04430385014bff11fd31fbd5f902f98cf84ef854f8a3f828f9;
    inBuf[3148] = 256'he5f9d3fad8fbf8fc44fe96ffa4001e01b40041ff0efdb1facef8fef787f822fa;
    inBuf[3149] = 256'h45fc77fe65001702f0033406c1081a0b6b0c010cdd09a4064e03d20091ff2eff;
    inBuf[3150] = 256'h03ff99fef5fda3fd50fe3e001203f005eb0796081608eb0698055c042403c301;
    inBuf[3151] = 256'h470024ffdffebaff9101bf035b05e905790560043303820256028002fd02d703;
    inBuf[3152] = 256'h2305fa062109250ba50c6f0da70da50d8d0d3e0d640c970add07b30499010cff;
    inBuf[3153] = 256'h4bfd15fc37fbe2fa6efb48fdbc006805870a5b0f3313cf1562170618c317c816;
    inBuf[3154] = 256'h28150e13d910a80e510ca40980061f032e005dfe12fe38ff1e01f5023a04c704;
    inBuf[3155] = 256'h00057d0590066308f20af70d4e11c914d117e019911a8019001715148c11fa0f;
    inBuf[3156] = 256'h7f0f3d0f2f0ee50b5d0852040e0151ff2cff5200fe01990338052707d009720d;
    inBuf[3157] = 256'h97118615a7185e1a671a04196e160913910fb70c290b5c0b050d5a0f5f111112;
    inBuf[3158] = 256'h3811850fe50d630da00e0d117f13d6143114ba11c70eca0ce60c6c0f4913e616;
    inBuf[3159] = 256'h15194a191f18cd16e6153415e613c310820b5805070059fd37feb8010b069409;
    inBuf[3160] = 256'h550bcc0b8b0c9b0e2e12aa16801a7c1c9a1c651be0192d1982196a1a5e1ba21b;
    inBuf[3161] = 256'hc51adb18f01546127a0e050b7c0884072a082c0a360da210f413f4163a197c1a;
    inBuf[3162] = 256'ha81a9f19d61739165f15af152817eb181e1a631a8d1900186616d0142f137711;
    inBuf[3163] = 256'h3f0f9e0c400a8108e7071409b80b150f71128c1467140f12320e310ac307c107;
    inBuf[3164] = 256'hf4094f0df10f6410940e5d0b4008b20600076a08be09ee094e099509ad0c1e14;
    inBuf[3165] = 256'h18208e2e5b3c9046f54aea4879412636a628ad1a6c0d1e0229fa70f650f758fc;
    inBuf[3166] = 256'hcc037d0b451128136f10e7092a0197f8adf2a4f081f283f743fea205360d9314;
    inBuf[3167] = 256'h2f1b0c20a7214b1fa4193212450bf5068905fd051607af079807c3070309990b;
    inBuf[3168] = 256'h370fea12ea152d18d319071b001c8e1c751cec1b581bf91a981a7b19ed16a712;
    inBuf[3169] = 256'h3b0d6208f405b406420ae40ee0115d11440de806f10015fe38ff53032108f30a;
    inBuf[3170] = 256'h520acb062b02b1fee5fd7ffffa01a7034a03f500f7fdacfbddfa82fb9dfcfefc;
    inBuf[3171] = 256'h16fc38faa6f8f7f82ffc7002d20a8513c61a8a1f7c2113212a1f611c1c198e15;
    inBuf[3172] = 256'hbc11d60d470a6707730585046e04d3043505fd04d703e001a4ff12fefdfd81ff;
    inBuf[3173] = 256'heb011b042505d604b303950208029f01760041fe72fb19f9b9f80ffb2bff3503;
    inBuf[3174] = 256'h7505d604660134fc60f6abf0a1ebdee72de64de74ceb3af19df727fd4e018b04;
    inBuf[3175] = 256'hb407b60a2c0c560a5b0462fbf2f267ef80f3e2fe160efc1b77242a2672222d1c;
    inBuf[3176] = 256'hcb15df0f8709c401c5f87df0bceb68ec59f214fbb002e3056b032ffc95f23fe9;
    inBuf[3177] = 256'hd6e1ccdcd4d9a1d876d9badc6ce2eee9b4f197f71cfa0af935f564f0a4ec54eb;
    inBuf[3178] = 256'hc2ec26f010f40ef703f8b7f62cf4f1f18bf12cf4d5f93c01a2083d0ece106210;
    inBuf[3179] = 256'hb80da50905052000b8fa01f597ef5febc2e9aaeba6f069f7ecfdee013602d8fe;
    inBuf[3180] = 256'hd3f8eff1b4ebcce679e37ce15be02ce020e1dae2e2e48fe609e727e691e445e3;
    inBuf[3181] = 256'h50e311e508e846eb71ed85edb9ebefe865e6ece5c0e8bfeee4f620ffd0042b06;
    inBuf[3182] = 256'h9302b0fa7ef017e6eadc20d64cd2b3d108d598dc9be792f40401500a4e0f0810;
    inBuf[3183] = 256'h410d5f08e5012df910ee57e1e9d43acc5fca19d0e0db02eaccf516fc2dfc70f7;
    inBuf[3184] = 256'hd2f021ebcde725e75fe84aea51ecf5eda2ee30ee3dec59e802e3f5dcbcd633d1;
    inBuf[3185] = 256'hdaccb0c919c879c8e7ca76cf7ad5b5db89e1afe630ebccefa7f4cef846fb30fb;
    inBuf[3186] = 256'h86f80df5f6f293f330f735fcd7ff52002efd28f749f034ea37e545e109de4fdb;
    inBuf[3187] = 256'he1d98cda50ddd1e1f1e659ebc3ee54f112f346f498f41cf3b2efd0ea21e5dcdf;
    inBuf[3188] = 256'hb7db5dd876d5bdd22fd097cea8ce4cd00ad3e7d522d830da02dd74e1ece730ef;
    inBuf[3189] = 256'h06f512f80ff81df6c4f4b4f58bf8bdfbe9fc58faeef421ef44ebbbeaa5ec60ee;
    inBuf[3190] = 256'he8edccea55e625e3f3e246e563e820ea5ce956e754e6fae7a6ec94f2d5f6bdf7;
    inBuf[3191] = 256'h53f503f12ded36eb8aeaaae905e716e255dcffd7c3d62ed9e7dd7ce255e515e6;
    inBuf[3192] = 256'h95e5bae5c0e76febd1ef7ff385f53cf65bf62bf69ef5edf34cf046eb6ae6b2e3;
    inBuf[3193] = 256'hece435ead2f168f987feb9ff79fd38f983f4dcf0b6ee75ed85ec52eb9ce939e8;
    inBuf[3194] = 256'h3ae823eaf2ed84f2d8f573f6e8f31fef52ea9ee7ede7f5ea34efd2f2eaf484f5;
    inBuf[3195] = 256'h2df5bbf46ff4ebf3edf26af1a0ef1aeef6eccdeb27ea8de72ae433e10be0a2e1;
    inBuf[3196] = 256'h57e647edaaf4effa04ff98004b00fafe54fdf2fb0afb99fab1fa2ffbb8fb01fc;
    inBuf[3197] = 256'hb8fbeefa64fad6fa9afc84ff7102d103e002bcff38fba1f6c9f295ef8fec50e9;
    inBuf[3198] = 256'hf0e545e340e22fe3bce52ae9e5ece8f08af50cfb2801d106df0af40c9e0d0d0e;
    inBuf[3199] = 256'h5d0f9a118a135113670fb207cefd4af493edf3ea06ec36ef9df2c8f451f5ccf4;
    inBuf[3200] = 256'h36f4b0f419f79dfbce01b808dc0eb2124e139f109a0b0e06d401e9ff19004c01;
    inBuf[3201] = 256'h2a02c4011a00ecfdf3fb65fa08f969f756f563f3a1f2faf3adf725fd61038809;
    inBuf[3202] = 256'h360f66140e19841c891dd51add13920951fefaf4e4efdcefaff30bf9cdfdc700;
    inBuf[3203] = 256'h4202860385054e081d0bb30c770c150bc7098e09a70a1c0c830c490bf408ce06;
    inBuf[3204] = 256'h0806a7067b07f806220476ffb2fa7df797f6b2f7acf9a7fbacfd3900c7033208;
    inBuf[3205] = 256'h7f0cd40f23120814a316cb1a112046253429bc2a6f298225111f5f16330ca001;
    inBuf[3206] = 256'h5df840f2f2efe3f0b7f38cf642f844f9c8fa2efe4204750c66158d1d8023b926;
    inBuf[3207] = 256'h94277526e4238320a51cc7188a15021303112e0fba0c9009b1065305bd069f0b;
    inBuf[3208] = 256'hc912e619b51e8d1f6d1c0c175c11d10c190ad708a2089609d80b710fd8139e17;
    inBuf[3209] = 256'h9919a1194318c71635160b1607152b12540d4308eb052e08220fd0187221fa25;
    inBuf[3210] = 256'hd7257f22e41ef31d52208e244f282e294f26e620c71a97152212d40fd40ddc0b;
    inBuf[3211] = 256'hfd09dc081b09150a8e0aae092d073a045a0394067b0eb419e224762c572e562a;
    inBuf[3212] = 256'ha422b11af5148f122713c1149b153a15b313e7114311531202151f19dc1d4522;
    inBuf[3213] = 256'had253b278926ef23e41f461b151779135210b10d950b7f0a2f0b840df510ab14;
    inBuf[3214] = 256'h4e17921899197e1b4a1f8225da2c27339d36ae35ea2f6326931a6a0e4004d2fd;
    inBuf[3215] = 256'h41fcd2ff1d07e80feb17011d7a1e3c1d6b1a55171e15d9138513a7147c17331c;
    inBuf[3216] = 256'hb622a829152f5931562f72297b216b194c1373105f10d0117913af13af111f0e;
    inBuf[3217] = 256'hfc099d066d05cc06870a201088161a1dd4235e2a6c30d035b539393bbb398034;
    inBuf[3218] = 256'h7e2b9c1f2a1269051cfce6f72ff90bffef062d0e281321159514ac12de0f660c;
    inBuf[3219] = 256'he60826069b05fe08a510361bf3254b2ddc2e902a2522b2183611da0c6e0b120c;
    inBuf[3220] = 256'h540d5f0e440fea0f271005108b0f500f6a106a133d18d71d0222012388206c1b;
    inBuf[3221] = 256'hbe15fe1143110a13b715091791157111cf0bbb062b049f047507540b3a0ec50e;
    inBuf[3222] = 256'hd20cda080604c1ff9afc9bfacef91dfafefb9200810895137420662c7d34d236;
    inBuf[3223] = 256'hd932d229521ec812df083c0179fb1af71ef4dcf22ff4c7f85100da090114ed1c;
    inBuf[3224] = 256'h66234127c128b9284328c72705276625f0210f1c1c14170ba50275fc26f960f8;
    inBuf[3225] = 256'h20f9d1f92ef9e9f65ef377ef5becefeaf0ebd5ef70f631ff2609b712611a481f;
    inBuf[3226] = 256'h1b214520c41d711adb165a13f60fdd0c8a0a6209a409390b390d360ecb0cfc07;
    inBuf[3227] = 256'h0400abf682ee09eadaeaaff06bf949022209280dd10e290fce0e2f0dfd089901;
    inBuf[3228] = 256'hedf756ee18e8c7e7a8ed9cf715026b097e0b79083f0282fbbdf636f502f77dfb;
    inBuf[3229] = 256'h5a010007210bc10c1c0b2b06eefef3f6f6ef95ebb4ea1aedaef104f7c9fb05ff;
    inBuf[3230] = 256'h390079ff38fd1dfa0af70cf5edf4eaf6a3fa15ff1203d0050407e206f6057d04;
    inBuf[3231] = 256'h2f02a1fe8cf919f317ecc6e58de194e02de3cae83df0a1f708fd6dffd6fe2bfc;
    inBuf[3232] = 256'h0df9e3f62ff6b9f6d7f7edf8faf936fb98fcbafddafd72fcfef9b2f7dbf62ff8;
    inBuf[3233] = 256'hfbfa7cfd11fe00fc06f8f8f329f198ef5aee00ece9e766e3b9e08fe137e6f6ec;
    inBuf[3234] = 256'heef237f6adf6daf517f67ff8f8fb37fe01fda9f709f02ae97ae5cfe5cbe8eeeb;
    inBuf[3235] = 256'hafed08ee1eee8cefabf209f6a8f714f67cf122eca6e877e84debd0eef6ef4eed;
    inBuf[3236] = 256'h60e73ce0bbda93d88ad96cdcbfdfc8e253e668eb24f280f922ffa9008ffd14f7;
    inBuf[3237] = 256'hb3ef55ea4be805e956ebd9edb3ef41f19bf2e7f24df10bed50e653dfe2dab1da;
    inBuf[3238] = 256'he7de76e50eeb8aed92ec88e922e74de733ea05ef47f4b8f86dfca9ff13020503;
    inBuf[3239] = 256'h2b0165fb64f21ee8e0debbd8d6d53fd4c3d1e8cc1cc65ac026bf9ac4ddd04ae1;
    inBuf[3240] = 256'ha8f1dbfe7f07e10bcd0d970e350e380c09088f011bfa31f392ed88e986e6aae3;
    inBuf[3241] = 256'h03e10edf2bdeb3de2de085e14ae255e2bde133e1dee03fe05edf6cdebfdd77de;
    inBuf[3242] = 256'h34e147e5b5e933ed8eeef2ed60ecbaeacae976e9c3e834e706e521e344e3a5e6;
    inBuf[3243] = 256'heeecacf475fbf1fe67fe88fadcf46aef27ebb2e78ce420e12fddb7d9bbd763d7;
    inBuf[3244] = 256'h91d894da6cdcfbdd72dfd6e07de23ee491e5cee695e830eb04ef82f305f773f8;
    inBuf[3245] = 256'h70f76df40bf19fee18edadeb00e910e4d8dd88d835d630d89cddc7e340e89fe9;
    inBuf[3246] = 256'h34e85ae643e67be84decbfefc3f043ef94ec6cea89ea26edc7f002f4e0f509f6;
    inBuf[3247] = 256'h48f555f40bf327f16aee13eb8fe85fe81feb67f03ff60ffa73fa52f7e6f1a7ec;
    inBuf[3248] = 256'h85e9f6e88aeae2ec5aee4beebbec1bea70e780e599e416e5bee6c0e886ea72eb;
    inBuf[3249] = 256'h18eb17ea7be9f9e9e9ebaeeebbf0def0d6ee61eb37e800e74fe88feb47ef04f2;
    inBuf[3250] = 256'h54f3b2f322f4a9f572f8cafbd0fea700c30024ffd5fbe3f6d2f06deab7e4fde0;
    inBuf[3251] = 256'hebdf17e192e338e623e87ee913eb7eedf6f011f5e1f8d1fbcdfdecfe3fff49fe;
    inBuf[3252] = 256'h21fb86f552ee76e7a4e3cde4b0ea23f3f5fa48ff24ffa2fbe6f6f8f283f0e3ee;
    inBuf[3253] = 256'h49ed49eb36e93ce801e9d8eaa5ec54ed76ec32eb78eb6bee02f4d9faa400c303;
    inBuf[3254] = 256'hfe033a021600defeeafe0900cc01c103df050a08a909f5092a08020421fe89f7;
    inBuf[3255] = 256'h23f1aeeb35e779e3d8e010e0d3e1a0e6ecede3f584fc65005601b1007500fa01;
    inBuf[3256] = 256'h4c05ff08010b200ac406cb02a100b20161056e094c0b9f091405fcffd5fc82fc;
    inBuf[3257] = 256'hc1fd35fe00fc19f7cef167effcf141f98a022e0ab20dfa0cec0927074c060007;
    inBuf[3258] = 256'h8a071c060d0249fcc2f65af3f9f236f5f6f80afd6f00aa029e031103f700e1fd;
    inBuf[3259] = 256'ha6fa59f823f870fabefe0a041409d60cf00e7d0fd90e5a0dfb0a8d071a0307fe;
    inBuf[3260] = 256'h2df99ff52df40ef5b4f70ffb43fe0501a703fb069a0b2c119616651a5a1b3619;
    inBuf[3261] = 256'hc6144d0f070a9f0518025bff8cfd08fd4efe7201a2059809320cd10cbc0bed09;
    inBuf[3262] = 256'h420811074d06e7052a06be073c0b7510e41527192f184712b1087ffe21f7aef4;
    inBuf[3263] = 256'h55f776fd490484095e0c3d0d430db60d380fc9112715cb182e1cdf1e1420271f;
    inBuf[3264] = 256'h2d1cb017aa124c0e0e0b8c082a067703d60093ffdb002505ef0b61137219361d;
    inBuf[3265] = 256'h8e1e0c1e9e1c6d1a11178112240d3d08a6054806c109b70ef6120a154415c314;
    inBuf[3266] = 256'h0b154d17d31ab11d611e101c7417df124e1060104712ba13a612d70eb609eb05;
    inBuf[3267] = 256'h04065a0a39111018321cac1cb81a0618ed15da14be137e11250e6f0ac4076b07;
    inBuf[3268] = 256'h2409e20bc10e0711f21272159b18b91bc31d8d1d231bed176d15c9140a167117;
    inBuf[3269] = 256'hff16c313ed0d5607bd02d90103052f0bfb1147171c1a821acd19cd19621ba11e;
    inBuf[3270] = 256'hc022f125e0264f259221f81c3319fb165816e6169517c0178517e81623168115;
    inBuf[3271] = 256'h8f14e4129b10b80d9e0a2308c20602079109810ea8157c1e6327ac2e44335b34;
    inBuf[3272] = 256'h4d328c2e162a8d255721f71c25188f13ee0f220eef0ec4117215f2180e1b651b;
    inBuf[3273] = 256'ha11a0c19e1169014e111e80ea30cb80b940c7d0f8913a317621b4b1e66203922;
    inBuf[3274] = 256'h4b23dd22ca20041d6918c714061323137614661521157914b2145317371ddf24;
    inBuf[3275] = 256'hcc2bf62ff22f5b2cac27e123052202221d22b6206c1d9b18ae134910b50ea70e;
    inBuf[3276] = 256'h7e0ff10f870fab0e690d310cb50beb0b070d690f8812b8155118351937183e16;
    inBuf[3277] = 256'h2b142913ef13b015701784185e1895174e17cc17f318481acd1a871a7b1a741b;
    inBuf[3278] = 256'h2d1e7722722628286926dd20f8184611b80b9109ef0a700ea912a51696199c1b;
    inBuf[3279] = 256'h491da91ecd1fa72094205a1f461d831aa5175e1598130a1265102c0e940b8109;
    inBuf[3280] = 256'ha7089d09510c7f0fda119d126811010fe00cd00b1c0cb60ddc0f1f12cf143718;
    inBuf[3281] = 256'ha51c3c223228522d8e30d430c22dd927d21fb516a70d3905d4fd12f87df4def3;
    inBuf[3282] = 256'hf8f67cfd2306f40e8a157b180718721582129110820f720e950c860901067303;
    inBuf[3283] = 256'hb102cf0346060809800bcc0df50fe2112213d512b1107a0d610aa808d908110a;
    inBuf[3284] = 256'hc90ad7090207830330013301b0038007ac0a000c6e0baa09fd074e0761078207;
    inBuf[3285] = 256'hf3062305500240ff9dfc0dfbf9fa4ffcdffe3c0298053b08b209f50997094609;
    inBuf[3286] = 256'h5709c409060a910988086e07ce06fb0675071f072c057501b4fc73f811f621f6;
    inBuf[3287] = 256'h68f8d7fb27ff7701440274015aff5efc08f907f6e2f3eaf238f399f4e9f628fa;
    inBuf[3288] = 256'h4bfe340359088c0c8a0e540d8708e300e2f710eff3e769e36be1bde1e1e309e7;
    inBuf[3289] = 256'hb6ea8aee1ff292f533f918fd510179059f080e0a820939074e04df015b00bcff;
    inBuf[3290] = 256'h48fffefdb6fbe1f82bf6a1f4aef4aef5c1f6c1f678f4c1ef3ce9e8e185db85d7;
    inBuf[3291] = 256'h39d64fd7a5d9a8dbd9dcbedd3cdf7ce29be721ed5af106f3ecf1a9ef5cee19ef;
    inBuf[3292] = 256'hd3f104f56af614f597f181ed12eb9aebb3ee3ff395f71efa9dfa6df9e6f6e9f3;
    inBuf[3293] = 256'h07f120ee6deb02e983e646e4d6e28ce247e473e841ee85f48ff96dfb9bf9cff4;
    inBuf[3294] = 256'h5aee52e82fe4f5e133e1eee0fedf61de9cdcffda20daffd9ead9bfd982d936d9;
    inBuf[3295] = 256'hb4d98cdb8adebce2b7e76dec79f06cf384f4e7f3e9f1b2ee4beba1e8d7e640e6;
    inBuf[3296] = 256'ha0e608e752e7a6e709e83be98deb32ee60f006f125ef41eb80e6e5e1b5de04dd;
    inBuf[3297] = 256'h92dba1d9bed6dfd280cf1cce0dcf6bd243d7b2dbd1de2be05fdf36dd90dab4d7;
    inBuf[3298] = 256'h76d55cd42ad412d500d749d90ddc6cdf09e32ae7d7eb5ef083f4f1f7f1f993fa;
    inBuf[3299] = 256'hf2f9e1f7d3f4e2f09eeb58e56ede30d707d13acd22cc12ce61d258d7eddb45df;
    inBuf[3300] = 256'h84e006e04bde71db60d8dfd5f9d31fd367d33bd4abd5f0d7f3daefde7fe355e7;
    inBuf[3301] = 256'h94e9aae997e7e7e440e35ee38fe5d1e844eb09ecf1ea45e86be55be300e266e1;
    inBuf[3302] = 256'h48e13ce1e8e1e7e311e72ceb2aef65f14af1f7eee8ea79e69ee24cdf88dc22da;
    inBuf[3303] = 256'he0d757d6dcd518d6d2d685d7dbd7d2d899dbbbe03ce89df060f7f6facafa66f7;
    inBuf[3304] = 256'hc9f291ee30ebc1e8a1e6fae31ee1a1decadc2cdcdddc78de35e145e56aea6cf0;
    inBuf[3305] = 256'h67f6fbfa7efdc4fd1bfc95f9cdf698f3c6effaea44e5dfdf0bdc73da39db34dd;
    inBuf[3306] = 256'hb1de05df4fde78dd28de17e1aee5f1ea78ef41f2adf37df431f526f6e9f695f6;
    inBuf[3307] = 256'he0f4dcf116eeb4ea85e8e3e718e9b8ebf5ee35f2aef4def51af6e2f5ddf5bef6;
    inBuf[3308] = 256'h53f8d4f997fad5f964f725f407f1cdee19ee9eee7fef0ff09befd7ed41eb82e8;
    inBuf[3309] = 256'h64e6c9e502e7e6e913eeadf2ebf67efa47fd78ff70010f03f203ba03fd01f1fe;
    inBuf[3310] = 256'h8efbc6f850f757f7f9f7f9f786f660f34cefddeb5cea6eebeeeeadf328f852fb;
    inBuf[3311] = 256'hc3fc02fd4efdcafeff018106d60a460dc30c5109340457ff20fce2facefa6efa;
    inBuf[3312] = 256'hbaf8a5f5ecf1bdeef6ec99ec3ced8cee6af02ef355f7ccfcf9020c091f0ea811;
    inBuf[3313] = 256'ha2131614fc1256102d0cec067401c4fcadf98cf82ff932fb44fe18026f06cb0a;
    inBuf[3314] = 256'h270e7d0f3f0e7e0a3705e0ff6dfb24f8a7f542f3def049ef83ef3df23df7f6fc;
    inBuf[3315] = 256'h8401b8037403ce014e00c0ff07006d0028003eff76fe8efed9ffea01c103ca04;
    inBuf[3316] = 256'h3505aa05f6064609d30bb90d6e0e070e680d4f0d960d970d610c54091205ec00;
    inBuf[3317] = 256'h04fe10fdd5fd6fff6801d5032407ea0bea110b181d1d2420e7203020b31ea71c;
    inBuf[3318] = 256'hf6190516a810e50a17067703a903a70596072b08dd068d045e03c404f308050f;
    inBuf[3319] = 256'hc6143d180419b517d815371541164418241a5c1a3a186214b40f5c0b82083107;
    inBuf[3320] = 256'h24073b08c7096a0b330d9f0e6f0ff80f33107d108e113a1328153d17e918301a;
    inBuf[3321] = 256'he81b4f1e5d21c0240527e92634241b1fd6182913d10edd0bf209f1075a05c602;
    inBuf[3322] = 256'hf4001b0157045d0a29125c1ae2206724d3246b226b1e9d1add17a31616174c18;
    inBuf[3323] = 256'h79195e1a721aa9198318ea16e214ae12f80fb90ca00937078306c808230eeb15;
    inBuf[3324] = 256'hd91eaf26c92be62d662db02b832a432aa82a2e2ba62aa628d5258322451fec1c;
    inBuf[3325] = 256'h521b801a091bb61c5a1ffb2292263b29c82a9c2aad28db258922801f111e6d1e;
    inBuf[3326] = 256'h59207423292659273927252657256e2654293e2d58310634b3342e34bc32e130;
    inBuf[3327] = 256'h6a2fe72d4e2c7d2b722b442c452e6730f3315d33ad3465366639d93c8c3fed40;
    inBuf[3328] = 256'h1540383dc839523619335d30382d6529e8255b239d227a24f627d12b612fa331;
    inBuf[3329] = 256'had32b7331a3538377a3af33dd640fd4288433d42bf3f103ca73779337d2fb92b;
    inBuf[3330] = 256'h9c28d32576232b22c62129226d23ff24da26bc29d52d5a33203a91402f453147;
    inBuf[3331] = 256'h2d462c431140c53d973c173ca43a6137c132872d3c293a2723270a2812295229;
    inBuf[3332] = 256'h3a29372af82c8831ed36cd3a4b3be137f43050282c209c1915157312cc10cd0f;
    inBuf[3333] = 256'ha20f23107a11b8133616b218271b281dbc1ef71f4c208b1fbc1d801a14161011;
    inBuf[3334] = 256'hbc0bdd066803a001b00161038e0526076c07ce05b2022eff2dfc92faaafaccfb;
    inBuf[3335] = 256'h34fd3dfe7efe65fea9fe9eff600180032205e505c705e804bf037d02f3002dff;
    inBuf[3336] = 256'h5afdb5fb94fad5f9c7f8d0f6c7f367f04aeef5ee13f3fdf9a501b207820a7d09;
    inBuf[3337] = 256'h6a05c5ffabf9eff3fceeb8ea5de762e5d6e4c6e507e8ccea88edf8efaaf1a2f2;
    inBuf[3338] = 256'h17f3f0f284f26cf2edf275f424f734facbfc0afe0efd04fae4f5c1f125ef1eef;
    inBuf[3339] = 256'h75f172f5bef95cfc28fcd5f889f29aeab2e2b6db6bd610d30ad139d0e0d0fad2;
    inBuf[3340] = 256'hd2d66cdcd3e22fe9e3ee49f38af602f964fa60fa8ef86ef491ee48e8cde256df;
    inBuf[3341] = 256'h36de6dded9de82ded0dc7ddad0d89dd885da43de79e20fe63ee878e82ae7f9e4;
    inBuf[3342] = 256'h02e28ddeb6da54d6f7d163cee9cbe6ca24cbcacb8ccc75cd9bce90d050d3dbd5;
    inBuf[3343] = 256'h55d7fdd695d463d1f4ce16ce2ecf59d1e9d25ed314d3ded256d4e6d71adc4edf;
    inBuf[3344] = 256'hd8dfc8dc8ad742d247ce7dcc3dccd4cbffca7dca70cba1cf54d79de05de961ef;
    inBuf[3345] = 256'h22f152ef23eb42e5aade99d7f5cff0c899c326c0bebe42befcbce5bac5b8c3b7;
    inBuf[3346] = 256'ha5b98fbebcc471ca00ceb2ce0ecedfcd27cf79d2edd6f8da2dde82e033e2f1e3;
    inBuf[3347] = 256'h6fe5bae561e414e149dc76d7a7d38ad198d150d315d67bd977dc32de5fdec4dc;
    inBuf[3348] = 256'h41da8cd8c6d88adb5de04ce5b5e8e8e90be9a7e73ee7fae77de9beeaa3eab5e9;
    inBuf[3349] = 256'h33e914ea51ed69f275f744fbf2fc2afc5cfae0f85ff8fff915fe2d048b0c9e16;
    inBuf[3350] = 256'he7208e2a4432bb365738b93792357c333832c13189322e34033631385b3a323c;
    inBuf[3351] = 256'h6e3e4041bd4462497c4ef7526e5628583058db57d7577e580e5a745ba25b8c5a;
    inBuf[3352] = 256'h2958215597529650d74e114d8c4a69478c4498428242d144db48eb4df0525356;
    inBuf[3353] = 256'h8a5790568d53e94fe14cb34aa949084931478e43d53de435012d4424361c0116;
    inBuf[3354] = 256'h14120e10f30ff610c3110d1288113310280fa50e180e200d890a7e05d0fe47f7;
    inBuf[3355] = 256'hddefebe904e517e040db9dd6ded299d1f0d2c3d5c4d8dbd9c8d759d3d6cdbcc8;
    inBuf[3356] = 256'h54c537c34fc1fbbed2bb7db838b656b589b5efb531b50fb354b0f9ad48adb5ae;
    inBuf[3357] = 256'h54b13bb492b6d1b7bcb822ba00bc35bed7bfa0bf87bd19ba3fb6a8b330b3a0b4;
    inBuf[3358] = 256'hb6b76fbbb3be8cc1f5c305c68fc887cb63ce35d165d387d477d59ad632d820db;
    inBuf[3359] = 256'h08dff8e2ede64feaa0ecabee7ff0a7f19bf22df321f394f312f580f741fbb1ff;
    inBuf[3360] = 256'ha5031b07cc092d0b910bbd0a48083705ba02bf016b0347075a0b180e3a0e820b;
    inBuf[3361] = 256'hbb07ad040203dc02f1025f01d6fde4f869f31eefe0ec23ec73ec16ed09ed52ec;
    inBuf[3362] = 256'h1feb1ae993e6f8e34de14bdfa5de3bdf0de1bbe325e6b9e71ce8b7e6d1e3fbdf;
    inBuf[3363] = 256'h5adba9d69ed244cf02cdf8cb72cb15cb73cac1c833c66bc3cac04cbf7abfc1c0;
    inBuf[3364] = 256'hc9c2fcc465c62bc7bfc713c898c841c903c95cc7f5c37cbefbb7dfb117adc8aa;
    inBuf[3365] = 256'h08ababacf5ae36b1ffb268b561b9f0be23c6d6cd0bd427d8e4d911d9bad645d3;
    inBuf[3366] = 256'h2dce07c880c14abb82b763b74eba68bfbac410c88bc934ca16cbe9cdb1d2b2d7;
    inBuf[3367] = 256'h01dcd7dee5dfaee0f7e104e354e3aae1efdc70d6e9cf8ccacec77fc712c80ac9;
    inBuf[3368] = 256'h0dcaefcae3cc7ed052d55adbeae1c9e78fec9cef1cf031ee0cea03e418dde1d5;
    inBuf[3369] = 256'haece1dc85fc2a6bd4cbacbb74cb534b2d2ad83a8b1a37ca0d09fdea156a5e9a8;
    inBuf[3370] = 256'hf1ab40ae0fb11bb638bed9c97ad869e86cf865071814491ea6258529572a9828;
    inBuf[3371] = 256'haa243c20871cfa19b519d61b761f85240b2a652e8e316c33ce331e34cb34ed34;
    inBuf[3372] = 256'h63344c32f32d38291e260226652a4132c83a5542bf47564b8e4f5855285c5a63;
    inBuf[3373] = 256'hab686a6a9b695a67ff6466642565166641673b685869196c55702175f979617d;
    inBuf[3374] = 256'hb47ecf7ee67d587cba7a72788e75157378719771f57332771d7af37bd17ba47a;
    inBuf[3375] = 256'hf979017a077b857c857c8b7a0377fa71ce6c78681364445f9c59125276490a41;
    inBuf[3376] = 256'h2b390733fe2ec22be228d4257021671c9217c012a60e550bb7074904d3016a00;
    inBuf[3377] = 256'h2f01570423086c0b090dac0b08085003b9fde0f7c4f175ea4be23adabfd2e1cc;
    inBuf[3378] = 256'h2ec9e7c6abc56bc5bfc5ecc663c9a9cc5ed06ed45bd81ddc2de037e4ade753ea;
    inBuf[3379] = 256'h66eb8aeaace8a0e63be5d3e57ce846ecc6f0eef4a9f785f9e5faa8fb92fc93fd;
    inBuf[3380] = 256'hf2fd5efe4effc900f30307090b0fe215f01c39234029302fa0343d3a1940c345;
    inBuf[3381] = 256'he64b8352f358685f6265086abe6d7c70f171b772c472e77103717e708570ae71;
    inBuf[3382] = 256'h59736f74a2748c737d71c96ffa6e1b6fe16f0a700c6f886d196cf96be86da270;
    inBuf[3383] = 256'hbb72f9720c70b76aee64be5f6b5c645b355b1e5bea5adc596c581b570e552252;
    inBuf[3384] = 256'h4f4ef048e942533d2638dd333330b42b2d26c51fa0187812710e4d0c110c8a0c;
    inBuf[3385] = 256'hb80b4909280578fff0f96ef5c8f163ef8bed13eb2de8bfe4a0e0c4dc62d93cd6;
    inBuf[3386] = 256'hccd3c6d19acf6ccdd9ca7ec7adc36ebf23bbc0b7afb542b58fb6a2b89bbafdbb;
    inBuf[3387] = 256'h55bc17bc1fbcb6bc01bea2bfacc0cbc009c0a0be52bd7bbcf8bbf2bb32bc7dbc;
    inBuf[3388] = 256'h50bdbabe94c04ec3c6c6a2ca1ccfa0d335d7b7d9abdae5d9afd8e4d7bed7e8d8;
    inBuf[3389] = 256'he2da77dcb4dd93def0deeedf20e22de55ee944eeaff266f6ecf886f9f0f8e2f7;
    inBuf[3390] = 256'haff696f60ef86cfa9dfd01014c035e040f04d4016efea9fac2f6c2f32df250f1;
    inBuf[3391] = 256'hd0f01cf04aeea6ebe4e84ee69de4f3e356e35be2e4e0b3dea1dcb3dbeadb45dd;
    inBuf[3392] = 256'h4bdf9de0b2e093dff8dc68d988d50ad14fcc07c818c41dc1c4bf6fbfe0bffac0;
    inBuf[3393] = 256'hd4c17dc25fc3edc34ac497c4e9c36ac2a6c04fbe07bc52ba7bb8b1b628b541b3;
    inBuf[3394] = 256'h94b1a2b0e1afc3af62b0f5b0eeb175b3ceb465b61cb8fbb862b952b9f7b7cab5;
    inBuf[3395] = 256'hf6b20daf1fab1da84ca693a6c9a898ab31ae8caffcae52ad4fab89a9c8a88aa8;
    inBuf[3396] = 256'hf8a7f5a61ba59fa270a0689e2e9cc7997d968d92768ff68dda8ed292c498819f;
    inBuf[3397] = 256'h9ba635ad6db360ba47c288cba7d6f3e2daefcdfc36082b115d175d1a551b051c;
    inBuf[3398] = 256'h261dbf1f0e249d28b12cd12fe8304230542ea02ac1257f20ee1a37164d13f411;
    inBuf[3399] = 256'h8312e1144718fb1cf922a4291831de384c40d747654faf56045e58647a68836a;
    inBuf[3400] = 256'h316afe67b965e6639e627362b3620d637e64fa66586adb6e68730877e679bf7b;
    inBuf[3401] = 256'hbe7c737d5a7dfd7b57794175a870e46ca26ab26a026d4470c073a276cf77a977;
    inBuf[3402] = 256'hb876d474b37286706e6d726986642b5e27571350bb48b2411c3b7334442ee728;
    inBuf[3403] = 256'h0524ea1f261c99173412dd0b7a0434fd9df682f051ebb1e6f9e1ddddbcda71d8;
    inBuf[3404] = 256'haad741d84ad9c3da60dc8eddb7ded2df1ce06ddf7fddeed932d5dfcf49caf0c4;
    inBuf[3405] = 256'h01c06ebb4db7b3b3b9b078aed5accfab70abd4ab56adfeaf71b330b781ba04bd;
    inBuf[3406] = 256'h07bf03c1a5c357c7b4cb35d05cd48cd7f4d904dcb3dd50dffce051e2b4e394e5;
    inBuf[3407] = 256'ha3e725ea21edd1ef64f245f530f891fbb2ffef034408c30cf2101b158119a51d;
    inBuf[3408] = 256'h6e21a824bf26e7278828f7281e2a872c24301935f23ace407046934be14f9b53;
    inBuf[3409] = 256'hc356fc58345a445a1c5938571c553c53fd514251bc501950fa4e6f4dbd4b094a;
    inBuf[3410] = 256'hd548704898485949784a2d4b5b4b074be849774822478b45bd439641673e7f3a;
    inBuf[3411] = 256'h83368d32312f8f2cb12919269f21371c9d164311340c1a08e304da0138ff04fd;
    inBuf[3412] = 256'h03fbe1f9abf9c7f951faddfaa0fad5f963f8f9f542f390f0d6ed92eb93e940e7;
    inBuf[3413] = 256'h9fe475e19dddb7d927d637d365d182d036d051d04bd0fccfb5cf86cfc9cfd9d0;
    inBuf[3414] = 256'h57d2eed33dd593d5ebd4acd3fad14cd0facec2cd9ccc7ccb28caf1c828c8dec7;
    inBuf[3415] = 256'h78c810ca70cca5cf40d380d63ed92adb21dcf8dc13de4edfdfe031e237e203e1;
    inBuf[3416] = 256'hbbde80db7ad849d6bcd432d478d4d4d4a1d506d788d88eda19dd5fdf88e1a1e3;
    inBuf[3417] = 256'h27e58ee61fe868e9bbea32ec25edb5edebed53ed5dec54ebece98ae83ae75de5;
    inBuf[3418] = 256'h36e301e182de57dccfda69d946d856d714d6f2d459d406d437d4d4d439d599d5;
    inBuf[3419] = 256'h1bd678d610d7ccd7dcd73bd7d7d566d3add02ace99cb66c9c8c774c61ac633c7;
    inBuf[3420] = 256'h41c90dccdece6dd09bd0c1cf46ce78cd07cea1cf32d20ad51bd781d84cd941d9;
    inBuf[3421] = 256'h05d9a8d8a9d76dd6f8d4dbd2a3d08dce6dccfeca92caeaca5dcc9acec5d001d3;
    inBuf[3422] = 256'h40d538d78ed944dc93de45e0cee09cdf84dd64dbbed98bd9b0dafddbb5dcfadb;
    inBuf[3423] = 256'h50d9cdd597d278d073d054d213d572d8f8db35dfc4e284e687e99beb4dec3deb;
    inBuf[3424] = 256'h7fe909e820e743e7f5e705e823e726e514e2f8de8bdceeda80dafddaa8db2fdc;
    inBuf[3425] = 256'h1cdc14db6ed97dd7afd591d414d4ffd31ad4d7d317d302d279d0c3ce2dcd94cb;
    inBuf[3426] = 256'h49ca7cc9b6c8f4c710c780c5a1c30bc22dc150c24ec6fecc50d65ae176ecf8f6;
    inBuf[3427] = 256'h4900e507980ea7149719c01dfa20f522d4244127362a642e37334237683a213c;
    inBuf[3428] = 256'hd73bbb3a583994379a36733641367e36d3366d3655361837c2389a3c4d42f947;
    inBuf[3429] = 256'h114d2351cc53fd5510580a5a9f5c4d5f7161bc6320668968b36b026fc5716c74;
    inBuf[3430] = 256'h937633783d7a477cb87daa7e477e597cc5798e76fa72c96f9b6c876938677065;
    inBuf[3431] = 256'h616456646b644664ed63c4622b61b15f065e905c865b375ae058885753557452;
    inBuf[3432] = 256'hff4e664a6f45c4403e3c9e381236b933a831b22f082dfd29ab269e22661e201a;
    inBuf[3433] = 256'h48154110f40ac50434fe8af7cdf0f9ea77e60be302e1f1dfeedeeadd8fdc67da;
    inBuf[3434] = 256'hf9d78bd514d327d1e9cf04cf8ece51cecfcd18cd2bccd8ca67c926c81ec776c6;
    inBuf[3435] = 256'h4dc675c6b5c6f7c609c7bbc63bc6ccc593c504c664c767c9e3cb87ce9bd00fd2;
    inBuf[3436] = 256'h29d3f4d30ed502d796d9e8dceae0e9e4cfe884ec5def85f16ff32af594f767fb;
    inBuf[3437] = 256'h4b001c066c0c35125717f51bca1f312342268728522ae12b142d7f2e51300e32;
    inBuf[3438] = 256'hdb33c2358937b939a33c0040cc439847b94a384d1f4f6e509751a0523f537553;
    inBuf[3439] = 256'h1a532d5229515150d14fc84fda4fc94f7e4fbe4ecd4d174d7f4c154cc64be54a;
    inBuf[3440] = 256'h2c498e46d442863e503a6a365b333c31692fb32dd72b39292326e4225f1f121c;
    inBuf[3441] = 256'h2f19471694131e117f0e170c160a3308e40661064d06e006d20727089107c405;
    inBuf[3442] = 256'h5f0217feb0f974f5f1f12cef9cec3eea12e809e685e490e3b4e2b8e15fe08fde;
    inBuf[3443] = 256'hc9dc85dbfada3adbeddba4dc2edd64dd54dd36dd04ddaadc41dcecdbe4db6bdc;
    inBuf[3444] = 256'ha5dd74df77e14fe3d1e4d6e56ee6d8e61fe765e7efe7d0e825ea17ec63eeb1f0;
    inBuf[3445] = 256'hbcf212f48cf486f44ef44af404f599f6faf805fc27ffd401d603ed0428051905;
    inBuf[3446] = 256'h2c0597058e06d5070e09280a190bf80b140d4e0e390fb20f9f0f060f650e070e;
    inBuf[3447] = 256'hc90d930d2f0d5a0c750b070b3f0b3c0c9a0d580edb0d1b0c54094706c4030702;
    inBuf[3448] = 256'h1801c50088003700d9ff2cff37fe28fdf4fbfdfac8fa29fbccfb3cfc9bfb9df9;
    inBuf[3449] = 256'h9df6f7f25def66ecdfe9afe7e6e54be41be3bde2d5e201e3ece202e259e07dde;
    inBuf[3450] = 256'ha9dc37db37da08d97dd7bdd5d4d376d23dd2dbd20cd478d56ed6ecd648d793d7;
    inBuf[3451] = 256'h12d8bfd821d937d9fcd83dd86ed7d1d641d621d68dd622d7ffd7fad872d971d9;
    inBuf[3452] = 256'hf5d8b8d74ed634d565d45bd420d51ad64cd789d84fd9fcd9c9da71db50dc53dd;
    inBuf[3453] = 256'hd3ddf2dda6dd9bdc87dbd4da59dab5da06dca1dd99df95e1b0e22ae320e34ee2;
    inBuf[3454] = 256'h8fe15ee14ce194e110e2f2e170e1c2e0acdfbcde3eded3dda7dd93ddfcdceedb;
    inBuf[3455] = 256'h6dda47d8f5d5e2d32cd222d196d018d08ecfb5ce69cdfacb69cac3c84bc7e6c5;
    inBuf[3456] = 256'hadc4fcc3c3c316c40bc534c674c706c9dfca45cd95d0a6d474d905dffce443eb;
    inBuf[3457] = 256'hbcf1d3f745fdc701e80400078508a009fa0ade0cf70e6a1107142416df171e19;
    inBuf[3458] = 256'h45199b184c172015da120e11ac0f3c0fde0f0311ca121e158f17751ad31d4621;
    inBuf[3459] = 256'h18250f299f2c0a302c33be355238093bd63d3a410345cc48d94ce650bb54c058;
    inBuf[3460] = 256'hab5c166011631365c865876546643562e35f4b5d8a5a0758ad558853a651a44f;
    inBuf[3461] = 256'h624dd04ad94706459e428040e43e753daa3bd63902380a365a3494321130252d;
    inBuf[3462] = 256'hc229e3258b22f31fc31d491c0d1b531945177d147610890b920589fe5ff76cf0;
    inBuf[3463] = 256'hd4e942e484df3edbcbd7e7d44bd238d025ce9bcbeec806c605c395c096bed0bc;
    inBuf[3464] = 256'h68bbedb939b8b7b657b523b43cb326b2b6b029af7ead25acb3ab33aca3adc6af;
    inBuf[3465] = 256'h01b2feb375b52cb652b6fbb563b522b541b5b2b5a0b697b75fb865b99fba3dbc;
    inBuf[3466] = 256'ha5be36c16ec34dc575c646c7bbc8f1ca14ce48d2acd6e6da27df19e319e7beeb;
    inBuf[3467] = 256'h93f072f552fa7ffe2302de05ba09640e4d14bb1a42216a27322cab2f60325834;
    inBuf[3468] = 256'h2c363a38f8393c3b003c0b3cee3b483c223d963e4c408c412e423a42ca417f41;
    inBuf[3469] = 256'hbe4195420b44c8456e47f148324a514b8f4cb14d884ede4e284e784c3b4a9c47;
    inBuf[3470] = 256'h31456c43f041af40a83f623e0f3de53b613a6638d3351e32972db82889239c1e;
    inBuf[3471] = 256'h3f1a22169712b90f1e0d040b50096107700593038301cfff9cfe68fd57fc46fb;
    inBuf[3472] = 256'hbff92ef8caf65bf528f40cf383f1bfefcfed90eb6de986e7b2e52ae4e5e2b5e1;
    inBuf[3473] = 256'hbae0dbdfe8dee8ddb1dc3adbbad94ad827d792d683d6f4d6c7d798d837d988d9;
    inBuf[3474] = 256'h70d923d9c7d85cd808d8bdd75dd71fd722d787d7a3d859da59dc7bde57e0c0e1;
    inBuf[3475] = 256'h0ce366e4f1e5ece7f3e982eb82eccfeca0ecb0ec57edb3eeddf04ff37cf555f7;
    inBuf[3476] = 256'h9ff850f9dff96ffa0cfb18fc92fd51ff68017d0320056e0666070e08d108a109;
    inBuf[3477] = 256'h050ae1091509a0073d069c05f0054b072c09a00a290ba30a1109fc06eb04f102;
    inBuf[3478] = 256'h210169ff84fd82fb99f9dff7a0f623f63ff6b4f625f7f8f6e7f515f4caf199ef;
    inBuf[3479] = 256'hffed00ed8fec82ec86eca6ec0aed8aed19ee8bee6ceea9ed6decd0ea47e92de8;
    inBuf[3480] = 256'h5fe7f0e6dae6b1e658e6c7e5aae429e3b4e17fe0f3df42e008e1ffe1dde23ce3;
    inBuf[3481] = 256'h4ce351e33ce33de337e3a0e28ae133e0b2de90ddfedc81dcebdbf0da29d91cd7;
    inBuf[3482] = 256'h62d53dd44bd494d560d77ad99ddb4ddddede81e0c4e1ace21fe3cae23be2fee1;
    inBuf[3483] = 256'h21e21be3d2e484e601e8ffe811e9afe81fe845e7a1e649e6d0e57de55de51de5;
    inBuf[3484] = 256'h16e557e570e579e559e5b1e4c5e3cde2d4e145e134e14ae15fe128e172e073df;
    inBuf[3485] = 256'h59de6dddf0dca5dc4cdca8db5bdaa1d8e7d630d5c1d3d2d219d2b7d1dfd15bd2;
    inBuf[3486] = 256'h6fd368d525d8e1dbb2e034e661ecfbf26bf9c2ffe405550b2a102d14df16b318;
    inBuf[3487] = 256'h0d1a291b091df21f56230e27402ad52b152c2f2b352940279b25dc238922a321;
    inBuf[3488] = 256'hd920fb2035220924a3266f299f2b992d662f0531633384360f3a613eef422a47;
    inBuf[3489] = 256'h7b4b8b4f2353f656d25a9e5e00639067ee6b58700d74a37687785379f378e077;
    inBuf[3490] = 256'ha07523720a6e6769df646a61fe5ea65d395dbf5ce05b885a6058ef5576538c50;
    inBuf[3491] = 256'hb24d1b4b5248e245f243e141fe3f183e603b52383035a7318c2e3b2c282aa628;
    inBuf[3492] = 256'h8c27f225f5238021101e201ace15ae10320b6b0503ffb3f8edf2aeed90e98de6;
    inBuf[3493] = 256'hf0e399e125df11dccfd8a3d598d249d0d1ced0cd46cde8cc47cc80cb92ca69c9;
    inBuf[3494] = 256'h71c8d1c761c74dc7adc761c897c97ecbdbcd5bd0c2d29ad491d5edd5f9d5dbd5;
    inBuf[3495] = 256'h08d6a2d64bd70fd8ded85fd9e1d99cda49db46dcc5dd5adf46e1a2e3d9e539e8;
    inBuf[3496] = 256'h08ebeaed4bf14df532f9fffcb000e5036f07fd0b73112d18c31ffe26b22dab33;
    inBuf[3497] = 256'h7638b83c98409a4323464348be496c4b9e4df74fa05211556856d5566a564755;
    inBuf[3498] = 256'h5854f3530c54ec542f566757b858cf597d5a0b5b1e5b8d5aab595558cc56ab55;
    inBuf[3499] = 256'hd2546254a75415557955d95592559e5453537a517e4fd94d2f4ca14a48497b47;
    inBuf[3500] = 256'h64455f432b41363fae3dd43b9139cc36fe32ba2e882a32263122a01ee01a4d17;
    inBuf[3501] = 256'h2e142d119d0e410c2209330563009dfa06f57ff030ed86eb06eb91eae2e9a2e8;
    inBuf[3502] = 256'hafe6dce487e3a7e295e2f5e22fe34ce305e315e2dee074dfe7dda6dcb9db12db;
    inBuf[3503] = 256'hc0da6fda03da8fd9e6d82ad881d79dd671d5fad3f9d1bacfafcdf7cbf4cabfca;
    inBuf[3504] = 256'h06cbc3cbe3cc2bcedbcf07d269d4f5d65ad933dbbcdc1cde4ddfa4e003e2f4e2;
    inBuf[3505] = 256'h78e374e3cbe20ae294e187e14ae2cce3ade5ffe77beab0eccbee9ff0cdf198f2;
    inBuf[3506] = 256'hedf28af2fcf182f1e5f092f097f082f08ef0d9f026f1d7f104f344f4acf518f7;
    inBuf[3507] = 256'h12f8e9f8caf976fa34fbf2fb1bfcbefbd8fa1df9eff696f4eaf152ef16ed13eb;
    inBuf[3508] = 256'ha0e9d6e848e8fae7d2e767e7f3e696e6f6e528e51fe469e24ee034de23dca7da;
    inBuf[3509] = 256'h0edae9d928dab1daf6da03dbf8da84daded957d9dcd8d9d893d9aeda1bdc80dd;
    inBuf[3510] = 256'h15dee3dd0fdd76dbafd928d8afd694d5e1d41fd493d354d3f1d2afd28fd209d2;
    inBuf[3511] = 256'h66d1bfd0aacf93ceb0cdb2cc19cc14cc34ccd5ccf3cde1cebfcf7dd09ad095d0;
    inBuf[3512] = 256'hc8d006d1c5d1f6d2ddd383d4bed43dd4c1d3b9d3f0d3b4d4a4d5e5d5a3d5ead4;
    inBuf[3513] = 256'ha2d3b1d272d280d20bd3c2d3f5d3fed30ed401d46ed470d596d603d878d96fda;
    inBuf[3514] = 256'h1fdb71db17db6eda9ad9a7d820d824d88dd868d93dda90da53da46d98ed7c4d5;
    inBuf[3515] = 256'h1bd4e9d28dd2b4d240d34fd489d5fed6f4d818db5cddd9df45e2e3e429e815ec;
    inBuf[3516] = 256'he9f092f650fcd401be066f0a290d360f9010e4119d13b115a118651c59207c24;
    inBuf[3517] = 256'h62283e2b402d672e692ed32dc22cf32afc280627f2246d239122112256222a23;
    inBuf[3518] = 256'h2024a7259f27ca29b22c2b30d9330d385e3c4c40134445478949494b5b4cda4c;
    inBuf[3519] = 256'ha14dda4ec450e653b657bc5beb5f7563f4659967fc672c67aa655c63a060fe5d;
    inBuf[3520] = 256'h3b5b6f58b6559a52534f374c16494e46f9438d41323ff43c803a463863364834;
    inBuf[3521] = 256'h0832672fef2b37289024de20ab1dd61acd17f0143d126f0f190d270bf308a106;
    inBuf[3522] = 256'hee037f00fcfcacf973f6c6f371f1eeee7eec0eea6de70ee5d4e258e0b2dd9dda;
    inBuf[3523] = 256'he0d6edd2e5ced5ca30c702c430c1f1be34bddfbb10bba6ba85bacbba77bb8ebc;
    inBuf[3524] = 256'h1ebe0cc020c20cc493c5a5c63cc782c7b8c7dbc704c85bc8d5c8b1c93bcb51cd;
    inBuf[3525] = 256'hfccf1cd317d6d2d84fdb32ddcfde7de0ffe1b1e3e9e53be8cfeabaed57f0bdf2;
    inBuf[3526] = 256'h1bf5fbf6a8f87efa2efc1dfeb900ca03b0079e0cec117017f01cc8212c26712a;
    inBuf[3527] = 256'h7a2ead322437693b7a3f3443484604498b4bb54da54f17517f51c850d24eb84b;
    inBuf[3528] = 256'h454814458042d1409e3f533eba3ca53a54385836e1340f34df33df33ff335834;
    inBuf[3529] = 256'hb1341e359735ae35713500352734323346321231c92f852e022d7d2be729bf27;
    inBuf[3530] = 256'h1925fc215f1e061b55180f1644147812f90f080dd8098c06bd03460196feabfb;
    inBuf[3531] = 256'h3bf83bf45ff0b6ec13e993e5aee119dd70d8f3d304d054cda6cba1ca5dca73ca;
    inBuf[3532] = 256'hc1ca8ecb82cc69cd56cef2ce49cfa8cfe1cffbcf0dd0c8cf46cfb7cef1cd21cd;
    inBuf[3533] = 256'h5ecc70cb97caf0c948c9b8c813c806c7e4c5d9c407c4f6c37dc40bc59fc5edc5;
    inBuf[3534] = 256'hb9c5a3c5e4c558c63fc761c871c9dbcab0ccc4ce4fd1fed35dd6add8ecda1add;
    inBuf[3535] = 256'hb4df99e26fe568e851ebf6edb0f03ff32ef58af612f7adf601f658f5dbf404f5;
    inBuf[3536] = 256'h95f529f6f6f6d9f7b9f80bfaadfb40fde5fe50002b01c9012a0221020702dd01;
    inBuf[3537] = 256'h70010501a4000f0064ffa8fed0fd3bfd39fdddfd44ff36013403f3043306c106;
    inBuf[3538] = 256'hbc0649065e0516048a02af00a3fe8efc74fa77f8a8f6e5f429f36cf18defaced;
    inBuf[3539] = 256'h01ec94ea8fe906e9bde890e862e8f7e76fe702e7b5e6cae672e784e805eaeeeb;
    inBuf[3540] = 256'hecede1efbaf127f32ff4dff407f5bef40ff4c3f216f15eefc9edccec9eecf8ec;
    inBuf[3541] = 256'hb0ed6bee9bee3eee67ed10ecaaea71e936e813e7efe581e404e39fe13be023df;
    inBuf[3542] = 256'h5fde9cddfddc87dc08dcd0db0edca0dcbedd5edf22e10ee3f4e475e6bee7e5e8;
    inBuf[3543] = 256'he6e91aeb88eceaed3fef46f0c1f0f5f0fcf0d1f0b0f069f0beefe2eee6edeeec;
    inBuf[3544] = 256'h4eecd6eb33eb3eeabde8efe670e580e459e4e2e474e5c5e5d0e587e56fe5dce5;
    inBuf[3545] = 256'h6fe606e751e7c2e6ade58de49ee3b3e336e5ebe712ec78f164f7e3fdb704460b;
    inBuf[3546] = 256'hd8115218121e41239f27a92af22ccd2e54306d321e35c537893ade3c073e783e;
    inBuf[3547] = 256'h223ec93c433ba039ad374436583586347534df3446354736a237f338d33ae23c;
    inBuf[3548] = 256'hb33ee6401f430d456f47f1494e4c364f23529b54175709594d5aec5bfa5dc460;
    inBuf[3549] = 256'h2d657b6ae56f5175aa79747c367ea17edd7d8c7c377af3766e73796f7f6b3168;
    inBuf[3550] = 256'h27656d623560d45d595bfa581156b352f84e4e4a28450e40df3a42367532be2e;
    inBuf[3551] = 256'h492b1b28c22406225920411f031f461ff61e351e0d1d111bdd189c16ba139a10;
    inBuf[3552] = 256'h560d9009f105b50259ff1efcecf846f5a5f150ee10eb39e8a9e5c7e29fdf25dc;
    inBuf[3553] = 256'h3ad867d4fed007ced0cb44ca04c900c8fbc6b5c556c4ebc276c135c04dbfc9be;
    inBuf[3554] = 256'hd2be6bbf77c0e0c195c399c50dc82fcb03cf3ed38ad762db48de60e0e7e1e6e2;
    inBuf[3555] = 256'hc0e389e4e5e410e550e599e57fe641e857eab4ec2def2ef10ff326f523f752f9;
    inBuf[3556] = 256'hcafb06fe5b0024033c061c0ae50ef21331196d1e182372279d2b512fd1321936;
    inBuf[3557] = 256'hcf384d3bbd3d07409e427a453a48ff4a8b4d8d4f5651d452de53b55427550b55;
    inBuf[3558] = 256'hc254385467539c528451e84fff4d984bd24821466943c9409b3ea83c153b233a;
    inBuf[3559] = 256'h75390739e838a1385a3854383c38433879384438c6372f3735365635de346334;
    inBuf[3560] = 256'h1e34fb33563360321c31122fa92c072ac62645238c1f2f1b9416e611090da808;
    inBuf[3561] = 256'heb04770170fe70fbddf707f405f0e5eb4ce830e53de2a0df0edd5dda15d845d6;
    inBuf[3562] = 256'he2d442d41bd41ed475d4ead45dd504d6a5d611d76ed796d796d7b3d7e3d72dd8;
    inBuf[3563] = 256'h92d8c7d8b0d836d823d7a4d5e8d3ffd148d0e9cec6cd0acda5cc5bcc65ccb5cc;
    inBuf[3564] = 256'h04cd83cd12ce62cebbce29cf82cf21d003d1e4d115d397d43cd668d80ddbcfdd;
    inBuf[3565] = 256'hd3e0dfe38fe629e9a4ebceed06f03ff23af44af656f813fac8fb48fd39feedfe;
    inBuf[3566] = 256'h61ff7dffcaff60000301e201a102a302fd01990060fef5fbbbf9b9f752f677f5;
    inBuf[3567] = 256'hb5f413f476f395f2b3f1f3f025f079ef01ef7cee18eefdedf6ed22ee89eecbee;
    inBuf[3568] = 256'heeee12ef08ef06ef41ef73efa0efdfefe9efe5ef0ef020f01ff004f05bef31ee;
    inBuf[3569] = 256'hbfecdfeae4e818e73ce579e3fbe16fe003dfcddd60dcdbda65d9b7d72fd613d5;
    inBuf[3570] = 256'h04d432d3b0d212d2add1cfd11dd2c9d2ccd374d4dcd437d539d556d5e7d570d6;
    inBuf[3571] = 256'h07d7add7ced79cd74dd77ed672d55bd4ded26ad167d0a2cf81cf13d0b4d071d1;
    inBuf[3572] = 256'h2fd268d281d2a5d260d209d29bd189d040cfe7cd18cc63cafac878c774c61fc6;
    inBuf[3573] = 256'hfdc57bc683c75bc854c986ca8ccbfdcc02cf13d15dd39fd525d739d8fad83ad9;
    inBuf[3574] = 256'h8cd910da60da9dda7cda88d90ed825d6dbd3cfd11fd0b6cedccd56cde5ccbecc;
    inBuf[3575] = 256'h9fcc63cc49cc21cceccb0ccc60cce8cce3cd02cf37d0d7d1e2d396d655dad5de;
    inBuf[3576] = 256'hdee33de947eecdf2eef688fae8fd6901e60492088a0c77106f146e18071c541f;
    inBuf[3577] = 256'h4d228b2441267827e527e927ba273227c5267e26f5255f259a2454230c22f320;
    inBuf[3578] = 256'hf21f801f901fcf1f9320c22124230f2542275529742b642d162f1d3184335436;
    inBuf[3579] = 256'he639e03dfb415c46964a764e1a5206550e576558d858a4584c58c6574657f456;
    inBuf[3580] = 256'h5b565755d3536851364e794a2646a741393db53865344b301b2c0d280524aa1f;
    inBuf[3581] = 256'h3e1bb616ec11780d89090c068403d5019200f3ffa9ff28ffacfefbfdb4fc49fb;
    inBuf[3582] = 256'hc7f9fef766f6f2f441f39ff1fbef1bee6cecfdea91e95ce829e79de5d2e39fe1;
    inBuf[3583] = 256'hd4dea4db0cd810d407d00acc37c8c1c48ec193bef0bba1b9dbb7ddb698b604b7;
    inBuf[3584] = 256'hedb7feb824ba5fbbb7bc5cbe4bc068c2a8c4d3c6edc82ccb94cd5fd0b3d34fd7;
    inBuf[3585] = 256'h3edb84dfb7e3dee7edeb55ef2cf294f443f6bdf76af9fbfac2fccefe6f00c701;
    inBuf[3586] = 256'he90255038503f1036a049205bc07610a9e0d5811e7149418931c8820b9241329;
    inBuf[3587] = 256'hee2c693092333f360039133c353fa24234468549d44c0450c1522d550457fc57;
    inBuf[3588] = 256'h6e586658f8579f574a57cf566456bb55ac547753e9510b50444e754cb44a3749;
    inBuf[3589] = 256'h8947854543438240a33d373b2939b137cd36c23584342a336c31d02fb12ea82d;
    inBuf[3590] = 256'he82c5f2c6f2b662a6d291d28e026c7254224a6220021db1ea81c811af6177415;
    inBuf[3591] = 256'h03133310600d850a3a07e8039f0018fdb8f968f6c1f200ef12ebd0e6b8e2e5de;
    inBuf[3592] = 256'h38dbeed7d7d4b0d1c3ce23ccecc986c8ebc7edc78dc88ac9bfca4ccc29ce46d0;
    inBuf[3593] = 256'ha3d200d521d7e5d826daecda54db75db83db9fdbd9db5ddc26dd26de72dfe2e0;
    inBuf[3594] = 256'h51e2d0e330e54ae634e7b9e7b4e752e77de639e5eae3a6e28be10be12de1e9e1;
    inBuf[3595] = 256'h74e385e5c7e73eeaa8ece6ee56f105f4f9f672fa28fec20148057a08430bf40d;
    inBuf[3596] = 256'h8510dd12211513178418a319621ab91ae51ad51a7f1a1a1aab193019c9185218;
    inBuf[3597] = 256'h951790163e15ae131912a110370fcb0d410c720a6408420622041b025400c3fe;
    inBuf[3598] = 256'h6cfd7cfcedfbbbfbf8fb5efcaefcebfcf4fcd8fcf1fc47fdd2fd95fe24ff21ff;
    inBuf[3599] = 256'h8dfe55fdb3fb3afa1ef97af863f870f856f810f873f796f6a8f57cf400f337f1;
    inBuf[3600] = 256'hf3ee67ecf0e99ee7a6e520e4b8e264e127e0cdde88dd8cdcaadbf6da80da00da;
    inBuf[3601] = 256'h8dd954d927d92dd983d9d6d918da4ada1bdab5d961d921d951d92ada6edb16dd;
    inBuf[3602] = 256'hfcdeb1e041e2aee3c1e4b3e583e6dce6ebe6b0e6f5e521e54fe449e369e2b2e1;
    inBuf[3603] = 256'he2e06ce06fe09fe035e1efe131e227e2e2e15de144e1d4e1bfe202e43de5f1e5;
    inBuf[3604] = 256'h57e6a4e6f9e6b9e7d6e8ffe91cebf5eb87ec1aedb3ed63ee2fefc5ef16f02cf0;
    inBuf[3605] = 256'hdcef59efc5eee7ede6ecdeeba0ea76e998e8e0e79ce7f7e7bde842eaa8eca6ef;
    inBuf[3606] = 256'h6ef3ecf79efc86016906b70a8f0ee4117714c7160f19381bc61dbb20b623fc26;
    inBuf[3607] = 256'h5d2a532d1b307832ea33d0342135b634553434342d34c534b3355736e236f636;
    inBuf[3608] = 256'h33363535fb3372325831a8304430c930f93178338d35a13735399c3a893b043c;
    inBuf[3609] = 256'hda3c0e3eca3f9542f8458b49484d6b50ac5265546b551a560b57f857e358df59;
    inBuf[3610] = 256'h525a425ae759f0589557fc55b353ee50e34d5d4ad0467143da3f2f3c5938ea33;
    inBuf[3611] = 256'h452fa22ad4254a21fe1c7b180a14ae0f3a0b4e071c04600162ffd5fd1efc75fa;
    inBuf[3612] = 256'hcbf800f7c4f53cf51cf593f52cf62ff6aff582f47cf234f0d5ed48ebece8abe6;
    inBuf[3613] = 256'h41e4f8e1cddfa4ddc4db12da4fd882d67bd418d290cfeecc4acad3c774c52dc3;
    inBuf[3614] = 256'h17c13cbfd3bdffbca9bcbfbcf7bc10bd20bd4abdd5bd1fbf13c187c34bc6edc8;
    inBuf[3615] = 256'h6dcb18cef9d069d49bd81addcbe192e6f2ea1fef51f325f7cafa40fedf00cc02;
    inBuf[3616] = 256'h3004b704f7046c05da05b2063308e209010cb50e79117914ba17a01a491dd41f;
    inBuf[3617] = 256'h02224d240a27052a672d05314d344137da39f63bf93d094006421a442646f947;
    inBuf[3618] = 256'hc549824b1a4db94e30504b51175266522c5297519550384fa94db84b6f49ec46;
    inBuf[3619] = 256'h0544f140ed3ddf3a00386335bd324330152e052c6c2a5229362811279b255323;
    inBuf[3620] = 256'h8f20891d3b1a36179314fa11b10fa00d6f0b7b09ab079f059b037d0114ffecfc;
    inBuf[3621] = 256'h0efb51f901f8bef616f54cf341f1f9ee09ed55eba4e915e82ee6b6e304e104de;
    inBuf[3622] = 256'hdadaefd711d52cd269cf8bcca6c9f7c653c4d4c1a0bf7cbd9fbb44ba53b90fb9;
    inBuf[3623] = 256'h86b962baafbb46bdc9be5bc0edc134c360c463c507c6a8c66bc74ec8bcc9b3cb;
    inBuf[3624] = 256'hebcd7cd015d352d55cd719d968dab0dbefdc09de49df76e048e1fbe15be246e2;
    inBuf[3625] = 256'h3fe24ce25ee2e7e2b6e37ae47ee58be668e785e8c0e9d3ea13ec51ed4dee7bef;
    inBuf[3626] = 256'hdaf044f217f42ff631f852fa76fc6efe9700ea02200555074709940a630bc50b;
    inBuf[3627] = 256'hb50b940b730b200baa0aec09a808160765059803fe01b60086ff76fe79fd44fc;
    inBuf[3628] = 256'heefa95f913f895f646f5f0f3a9f28df15ef034ef4fee8eed1ded3fedb8ed84ee;
    inBuf[3629] = 256'ha4efa3f061f1e9f1f1f19df13bf1b3f035f0f0ef9aef33efbdeed9ed9cec34eb;
    inBuf[3630] = 256'h78e9bce749e6f7e4e7e319e31ae2ece0a0df04de6bdc12dbc1d99bd89ed76ed6;
    inBuf[3631] = 256'h31d518d4fbd221d2a9d14ad126d141d153d19ad135d2ddd2c1d3e3d4e3d5e8d6;
    inBuf[3632] = 256'hf0d7aad855d9fed955daa2daf2daf3daf8da1adb12db3fdbbbdb36dc03dd25de;
    inBuf[3633] = 256'h33df6de0bee1b4e294e35be4abe4dde4fbe4b7e464e406e454e39de2dbe1cae0;
    inBuf[3634] = 256'hc1dfd1dee0dd56dd46dd87dd42de44df44e053e14ae20ce3c2e352e4ade4efe4;
    inBuf[3635] = 256'hede4a7e446e4b7e336e30ee331e3cce3e3e406e61fe725e8dbe898e9bbea32ec;
    inBuf[3636] = 256'h44eef8f0d3f3e9f646fa97fd1601c80423081c0b990d410f8c10ed116e139715;
    inBuf[3637] = 256'h7d189e1b041f782279254828dc2ad92c8e2eec2fa7304731e6315f3241336f34;
    inBuf[3638] = 256'h77359b368637c337bc3757377536c6354835d534eb34383557359e35c735b635;
    inBuf[3639] = 256'h06369e3677370b390e3b5a3d5340a0431547e34a754e81512c540f563d571d58;
    inBuf[3640] = 256'h6d584d580b585b577356b055d054f1532053d4511150ee4d2b4b30484d454942;
    inBuf[3641] = 256'h693fab3c99395a36e432e32eba2a8c262722041e351a6916fa12df0fba0ce409;
    inBuf[3642] = 256'h4a077d04cb0123ff3cfca6f987f7a7f56bf4a0f3b6f2d7f1dff085ef33eee3ec;
    inBuf[3643] = 256'h43eb92e9a7e744e5d8e285e040de65dcd8da46d9bcd700d6e2d39bd130cfaacc;
    inBuf[3644] = 256'h51ca2ec844c6b8c482c399c200c2a5c17bc170c17ec1b1c101c280c248c337c4;
    inBuf[3645] = 256'h5bc5c2c63ac8e7c9f4cb2acea7d07cd344d614d90edcf3de13e2b0e571e97ded;
    inBuf[3646] = 256'hd3f1e1f5c4f997fdef00090408077b099c0b980d220fa8107b125b14a3167419;
    inBuf[3647] = 256'h5c1c7c1fc922c02582281d2b482d5e2f88318a33a335d037be399e3b6d3deb3e;
    inBuf[3648] = 256'h4c40864175426f438a44c2455a471949a64afa4bca4cfe4ceb4c8b4cf74b6d4b;
    inBuf[3649] = 256'haa4aa0497c48f9462e455e434e41233f1a3de73ab138a7366f3441325930672e;
    inBuf[3650] = 256'hab2c4b2bcf29622818278225e92360226d204f1e121c5b19a8163914c911b50f;
    inBuf[3651] = 256'he70dd60bc009a507490535038501e3ff8efe53fdbcfb0efa46f837f648f474f2;
    inBuf[3652] = 256'h77f089ee8aec3feaf4e7b2e568e362e19fdfffdda4dc76db4eda42d937d817d7;
    inBuf[3653] = 256'hf6d5cfd4a9d3b0d2ffd1b5d1e8d187d277d37fd461d50cd683d6ebd696d7b2d8;
    inBuf[3654] = 256'h56da96dc3fdf1fe22de52fe800eba3edd6ef75f1a0f24df3a5f30ff493f43ef5;
    inBuf[3655] = 256'h3ef651f758f882f9a0faadfbeffc3cfe87ff09018a02ec0359058e0672074a08;
    inBuf[3656] = 256'hfe088f09450af50a7d0b070c780cda0c7e0d610e720fba10fb110a130314ea14;
    inBuf[3657] = 256'hca15c016b2177318ef181f19171905191219411972197e1925194118ea163615;
    inBuf[3658] = 256'h4c137611c70f380edf0c990b470a0a09ce0790067f057c046b0369024a01fcff;
    inBuf[3659] = 256'hb3fe4efdc4fb41fa99f8c9f618f56df3dff1aef0a7efc3ee2deeb1ed51ed35ed;
    inBuf[3660] = 256'h12edd3ec8cecf6eb29eb70eaace9fbe880e8e7e724e74be618e5a8e32ee277e0;
    inBuf[3661] = 256'haede10dd7cdb2eda62d9e0d8b4d8dbd8ead8dbd8b2d827d866d798d68fd58bd4;
    inBuf[3662] = 256'hb4d3dcd247d216d20dd260d207d39cd345d4f6d465d5e9d596d626d7e0d7b4d8;
    inBuf[3663] = 256'h48d9f7d9cdda91db9fdce3dde9deeadfd2e05ae1f6e1b3e24ae301e4b1e4fde4;
    inBuf[3664] = 256'h2ae531e5e7e4ace48ae461e486e4efe46be51ae6cde64de7c1e712e839e860e8;
    inBuf[3665] = 256'h6ae84de82de8fbe7d6e7e5e7fee71ee83de81be8d9e79de751e730e756e78ce7;
    inBuf[3666] = 256'h05e8dce8dbe934ebe8ec9aee71f07cf289f4f5f6f1f941fd12014e0575098a0d;
    inBuf[3667] = 256'h6811a7148917371a991c231ff421b9249527582a982c972e48306b315232df32;
    inBuf[3668] = 256'hdb32c132a5327632a532f032e532be32393239315c308e2fa72e092e622d902c;
    inBuf[3669] = 256'h2a2c202c682c632d942e9a2fb33089311b32f432e733f53488365d386d3afe3c;
    inBuf[3670] = 256'h9c3f09425d442f469a470b49684ad74b704db04e774fc04f3c4f294ebe4ccd4a;
    inBuf[3671] = 256'h9948384667436a40513dd8394c36a932a42e852a3b267821a01cc317be121c0e;
    inBuf[3672] = 256'hec09e805650241ff1ffc61f9f4f67df447f21df09ded30ebece8bee631e540e4;
    inBuf[3673] = 256'h8ee33fe308e37fe2e0e119e10ae010df2fde48dd97dcf7db35db71da8fd97ed8;
    inBuf[3674] = 256'h62d716d67ad499d268d01fce1bcc88ca8bc9fec883c8e8c70cc700c623c594c4;
    inBuf[3675] = 256'h54c46ac48ac4a3c4fbc495c59bc63cc818ca06cc20ce2ed06bd232d541d89ddb;
    inBuf[3676] = 256'h54dff0e27de62deaa1edfef078f4b9f705fba7fe4102f105bf09250d48106213;
    inBuf[3677] = 256'h2716d718941beb1d0a2029220d24fc250a28b229e52aa52bc02ba52bba2be62b;
    inBuf[3678] = 256'h452cc42c032d262d5b2da82d462e382f3b30453145322133f233ad343b35a435;
    inBuf[3679] = 256'he53516365d36a436db36e5368c36f4355535c634883497349e3496346134ca33;
    inBuf[3680] = 256'h11332c32c530fa2eb52cd029b82691233d20081dd91968160713b00f2e0cc708;
    inBuf[3681] = 256'h50057f01aefdeef93af617f37cf02cee61ece0ea61e922e8e8e66be5e2e327e2;
    inBuf[3682] = 256'h2be05fdec1dc43db18daf8d8b7d785d64bd51fd448d3a6d236d20ad2e6d1c7d1;
    inBuf[3683] = 256'hbcd197d16bd14cd119d1f4d0e3d0b5d085d050d0f2cfa7cf72cf2fcf10cf04cf;
    inBuf[3684] = 256'he9ce0dcf74cffdcfe0d0ebd1d9d2e4d303d523d69dd748d9d1da52dc99dd88de;
    inBuf[3685] = 256'h99dfece077e284e4d9e617e96aebb1edc3eff9f13cf44bf65cf849fadafb61fd;
    inBuf[3686] = 256'hd5fe090049017c026503450405056505aa05c00573051605af041a04b5038803;
    inBuf[3687] = 256'h62038303d50303042e043c04e2035a03b102bd01c700ebfffbfe36feb2fd2ffd;
    inBuf[3688] = 256'hcdfc8efc22fca5fb34fb9bfa01fa82f9cef8ecf7f7f6b2f550f414f3cdf18df0;
    inBuf[3689] = 256'h69efffed5becb2ead7e801e771e5e5e376e252e135e04fdfd0de61de10dee1dd;
    inBuf[3690] = 256'h6dddd4dc42dc71db94dac5d9a1d858d70fd689d41dd3f3d1bdd0b3cfe0cef8cd;
    inBuf[3691] = 256'h49cdf8ccbdccd8cc49cdaecd44ce11cfc5cf9dd091d13fd2dcd26dd3b7d313d4;
    inBuf[3692] = 256'h99d407d5a3d56ad614d7e7d7e4d8bfd9aeda9ddb35dcb9dc29dd4edd80ddc8dd;
    inBuf[3693] = 256'hf1dd4fdee2de63df0de0c1e023e181e1ebe14ee229e38ce425e60be8ede951eb;
    inBuf[3694] = 256'h6eec4fede8edb6eed2ef0bf198f24cf4d5f54ef78ef85bf9e9f931fa32fa38fa;
    inBuf[3695] = 256'h46fa54fa7ffaa2faabfab0fa98fa6efa41fae8f967f9c1f8d0f7c7f6c4f5c0f4;
    inBuf[3696] = 256'h05f4a8f37bf3a6f30bf456f4b5f425f57ff525f623f73ef8b2f965fb0ffd06ff;
    inBuf[3697] = 256'h5c01db03cd06080a130d0c10d61230158417ea19301caf1e5921e723a9268c29;
    inBuf[3698] = 256'h3a2ce72e54311b337f346a35b535de35e1359d35813568351535d53452343933;
    inBuf[3699] = 256'hec314530552eda2cd02b272b3f2b982bd92b5a2cc62c142dcb2d992e5b2f7530;
    inBuf[3700] = 256'h8e31a1322e34e135a237b5399f3b513d303ffe40e24237459247e449464c3a4e;
    inBuf[3701] = 256'hc94f1e51dc512b522d5283515850c54e764cb649af4622436c3fa23b6b371533;
    inBuf[3702] = 256'hb12efd2970253221f71c0c195f157811a80d060a4f06ee02f2ffedfc1bfa82f7;
    inBuf[3703] = 256'hcff468f27af0baee70eda6ecfcebaaebc2ebe7eb36eca8ecd6ece2ecf2ece1ec;
    inBuf[3704] = 256'hf9ec6aedfbedb3ee81ef06f02ff0f6ef2defe4ed46ec51ea26e800e6f4e31de2;
    inBuf[3705] = 256'hb3e0badf12dfb7de73defbdd5ddda1dcbfdb09dba5da6bda91da1ddbd8db0fdd;
    inBuf[3706] = 256'hdfdefde09ee3a9e6a0e9c0ec13f04ef3e6f6f1fafffe5903e407160c4e109714;
    inBuf[3707] = 256'h8e18ac1cf020d724bb28892cd02f1033603662397d3c893ff34100449b457e46;
    inBuf[3708] = 256'h3947df4732488248a2484548cf4747479d463846ea457545114595440944d943;
    inBuf[3709] = 256'hec433444cf445445a545f2450246f6451446104603461f461046fb450f46e245;
    inBuf[3710] = 256'h8f453d458644a643d642b1417040373f973dd13b193a0338d735b5332331652e;
    inBuf[3711] = 256'h9a2b4e28ca242721f91c99183214700fb80a2a066d01e5fcb6f8a0f40cf103ee;
    inBuf[3712] = 256'h24ebaae883e662e49ce231e1dcdfcbded7ddb7dcaadbb4dac7d926d9b6d849d8;
    inBuf[3713] = 256'hf7d7a8d75ed755d78dd706d8c3d88ed94cdaedda4bdb75db70db2cdbceda59da;
    inBuf[3714] = 256'hc3d93ad9b6d828d8b7d751d7e6d6abd691d691d6e1d65dd7e6d79bd849d9dfd9;
    inBuf[3715] = 256'ha3da90dbb8dc63de69e09ee20ee569e78be9a7eba8ed95efbbf1fcf34af6daf8;
    inBuf[3716] = 256'h7dfb19fedf009f033706d808500b7a0d880f4d11a712d013aa141c156b158515;
    inBuf[3717] = 256'h54152515f0149e1470144f140c14d21393132e13da12931221128f11ca10990f;
    inBuf[3718] = 256'h290eab0c140b8e093508cc0658050404b7028c01b600f1ff1dff50fe55fd35fc;
    inBuf[3719] = 256'h42fb57fa5df975f852f7e5f586f421f3c2f1a6f081ef2deee0ec69ebdbe989e8;
    inBuf[3720] = 256'h3ae7e2e5ace44be3c0e13ce076de73dc69da28d8efd519d476d222d128d01bcf;
    inBuf[3721] = 256'h12ce39cd58cca8cb44cbc9ca57ca0fcabbc9b3c91eca96ca2bcbc9cb0dcc46cc;
    inBuf[3722] = 256'habcc07cda0cd76ce1acfc3cf83d00bd19ed132d24dd229d2ddd13ad1cfd0d2d0;
    inBuf[3723] = 256'hf9d08ed17dd252d363d4b8d5f0d65dd8ecd91fdb48dc67dd13deb4de46df5adf;
    inBuf[3724] = 256'h5bdf5edf15df05df43df6cdfdfdf90e00fe1b4e174e2e8e26be3fce355e4dde4;
    inBuf[3725] = 256'h96e534e6f8e6c6e75ae8fae89fe91aea9eea05eb1eeb1eebf9eab3ea84ea4bea;
    inBuf[3726] = 256'hf3e99fe930e9cbe8b6e8d6e833e9cae93eea90eae1ea0feb5bebfaebb1eca3ed;
    inBuf[3727] = 256'hebee49f0f7f125f48ef654f976fc7dff6d024105a207cc09fb0b090e4c10ec12;
    inBuf[3728] = 256'h9b157c18881b591e10219c23982533276d281a29ae29512ad42a7e2b162c332c;
    inBuf[3729] = 256'h132ca62bce2a0f2a60298728de2733275326b4253c25c524bf24f0242525b625;
    inBuf[3730] = 256'h5c26e326a62775284929972a362c022e253037320834d8357d370a39ba3a453c;
    inBuf[3731] = 256'h9a3dd53ec53f97407c413842c9421243ba42ed41c6402f3f703d813b14395c36;
    inBuf[3732] = 256'h4b33b72f012c2528eb23a01f331b7616d511520dc10884048b009bfc0af9c2f5;
    inBuf[3733] = 256'h79f27defb6ece9e96fe734e5ece2d5e0cedeaddcdeda79d965d8e3d7b9d793d7;
    inBuf[3734] = 256'h98d7b6d7dfd75cd808d99ed922da5dda3fda0fdac6d95ed9e5d827d81ed7f7d5;
    inBuf[3735] = 256'hbcd491d382d265d12dd0d4ce5dcd00cccfcac8c9fcc847c8aac753c730c751c7;
    inBuf[3736] = 256'hd2c769c823c934ca70cb11cd47cfb3d166d47ad78bdacfdd79e118e5d7e8d5ec;
    inBuf[3737] = 256'ha1f079f492f874fc4e004404e307740b3e0fde128816611af61d7e212f25a528;
    inBuf[3738] = 256'hf42b1b2f99318f3343359f36f1375c397c3a3b3b993b783b223bd93a8b3a393a;
    inBuf[3739] = 256'hcc3923396238af371937a9362f368635b734ca33fa3278321e32db3195310f31;
    inBuf[3740] = 256'h6e30dc2f352f912ee72de82cc02b912a3229d7278026d6240d2346215b1fa01d;
    inBuf[3741] = 256'h201c751acb181c172715471382117a0f5f0d130b4d087805a902b0ffe1fc23fa;
    inBuf[3742] = 256'h2cf75bf4abf1f0ee81ec3aeadee7bee5cce3ede16ee01edfc5dd92dc60db23da;
    inBuf[3743] = 256'h17d90fd8ebd6c7d588d44fd369d2ced180d173d161d14dd150d16bd1cbd164d2;
    inBuf[3744] = 256'h04d3aed348d4d3d493d583d67ed78ad86ed917dacdda92db67dc70dd69de2fdf;
    inBuf[3745] = 256'hfedfcde0b3e1efe23fe46de596e690e771e89be9f8ea73ec34eefbefb6f1b3f3;
    inBuf[3746] = 256'hd0f5eff73efa78fc7cfea000cc02ed043a076409260bb80cfc0de90eda0fb410;
    inBuf[3747] = 256'h4711d2113a126512a212de12e812f112ed12c012b212c912cf12d812d5129712;
    inBuf[3748] = 256'h50122412f011b3116111aa108c0f390eae0c0f0b9a092808a8064a05e8037902;
    inBuf[3749] = 256'h3601eaff72fefffc6bfbb1f923f8a4f621f5caf366f2ddf06eeff5ed70ec21eb;
    inBuf[3750] = 256'hd9e98fe877e75ae633e531e41ce3fde109e10fe028df7eded7dd48ddf7dcaddc;
    inBuf[3751] = 256'h8bdcaedcd0dcfddc3add39dd1addf7dca0dc40dce9db5ddbc3da2eda77d9d5d8;
    inBuf[3752] = 256'h62d8f1d7aed7a9d7b4d701d896d834d9ecd9a9da20db7adbbfdbc5dbc9dbcfdb;
    inBuf[3753] = 256'ha9db98dbafdbccdb3bdcfddccbdddade1ee055e1c9e26ee4f0e581e705e92dea;
    inBuf[3754] = 256'h49eb5dec27edf2edb1ee16ef73efd2effdef49f0b1f0f6f05ef1edf177f239f3;
    inBuf[3755] = 256'h20f4dcf481f5f1f502f6eaf5b5f560f51df5f0f4daf4f5f429f55af56ff532f5;
    inBuf[3756] = 256'ha1f4d7f3e1f202f25bf1cff072f033f0e6efb9efbaefc8ef1df0c2f094f1e2f2;
    inBuf[3757] = 256'hc3f402f7c2f9dafcdaffd702c9057208120bad0df00f12122214fd1510187e1a;
    inBuf[3758] = 256'h001db81f6d22aa24a1264f288629b12ad22bb02cb02dc82ec02f01315d327733;
    inBuf[3759] = 256'h953466358e357535e534b8339232663129307a2f0f2f972e752e432ed42dc12d;
    inBuf[3760] = 256'hd62df72daa2e9d2fb2307d32bb344f37863ace3dce40c7435e469b48ee4a074d;
    inBuf[3761] = 256'hd94ea1500f5241538d54a4557d561c57fa562656e054ff52e050ca4e714c0f4a;
    inBuf[3762] = 256'hbe4715454242413f923b783726336e2ede29b7259421a91dea19da15cf11f00d;
    inBuf[3763] = 256'hda09d805f601cbfdd0f957f631f3cbf02defcaedc9ec30ecafeb9deb03ec68ec;
    inBuf[3764] = 256'hd5ec2eed1dedfdec01ed08ed49edacedd5edd3ed9ced06ed3fec50eb25eaebe8;
    inBuf[3765] = 256'hbbe790e683e590e49be3a0e2a8e1afe0aedfa2de70ddf2db49da9fd806d7c9d5;
    inBuf[3766] = 256'hfdd462d40fd406d420d4b1d4dcd553d73ad982dbd6dd98e001e4cfe73fec2df1;
    inBuf[3767] = 256'hf4f5b1fa61ffaa03ed07460c4f1055147118531c562085246528142c822f5432;
    inBuf[3768] = 256'he8346937a139d23bf33db03f364188426643fc433a44f5437843e4424342dc41;
    inBuf[3769] = 256'h91412541a440e43fe13eea3df43c023c3c3b6a3a8e39e2383e38ae375e37ff36;
    inBuf[3770] = 256'h9b3669362a36fa35fb35c2355835e53423345733c43210325731a6308b2f402e;
    inBuf[3771] = 256'hf82c622bc6293e285f266d2481224020f81daf1bfa1821162e13d20f710c1609;
    inBuf[3772] = 256'h6c05c5011ffe3bfa86f614f3bbefd6ec59ea03e810e667e4cce279e15ae04cdf;
    inBuf[3773] = 256'h8ade0adeb1dda7ddd3dd19de97de3adff1dfc4e091e143e2e0e269e3f4e393e4;
    inBuf[3774] = 256'h36e5cde52ee635e6f3e579e5eae480e43ce415e418e435e46ae4e1e488e53ee6;
    inBuf[3775] = 256'h00e797e7e7e720e84ce875e8cee839e98ee9f1e955eab8ea63eb4fec56ed9bee;
    inBuf[3776] = 256'hf8ef40f1b3f24cf4ecf5d6f7f1f901fc37fe6e00660256042806a7071809720a;
    inBuf[3777] = 256'h830b8c0c8a0d470e050fba0f1b1042100f10330fe10d420c480a490875069704;
    inBuf[3778] = 256'hc8021c0153ff89fdecfb3bfa81f8e2f61af53df395f1f5ef6fee3eed0aecbaea;
    inBuf[3779] = 256'h78e9eee723e671e4ade2fee0cedfdbde2fde08defcdd08de64deacdee4de3bdf;
    inBuf[3780] = 256'h3edff4de9bdee1dd0bdd70dcbbdb0cdb79da7cd934d8d7d619d555d3cdd126d0;
    inBuf[3781] = 256'h99ce45cdcacb74ca6cc952c862c7a8c6c1c5fec48ac41ec408c44dc476c4b6c4;
    inBuf[3782] = 256'h12c53bc58cc51ec695c62dc7d9c736c89bc824c995c95dca89cbb7cc28cebbcf;
    inBuf[3783] = 256'hefd00ed216d3bad381d485d56ed6a7d71cd956dac5db5eddaede11e056e1ece1;
    inBuf[3784] = 256'h42e263e214e202e237e23de26be292e249e218e214e2f8e130e295e2b9e2fae2;
    inBuf[3785] = 256'h53e396e330e40fe5dfe5d4e6c6e781e853e931eaf7ead0eb96ec23eda2ed02ee;
    inBuf[3786] = 256'h3eee80eea8eeadeea5ee72ee1ceec5ed5bedf4ecafec6bec33ec06eca5eb16eb;
    inBuf[3787] = 256'h6dea9de9f8e8cce81be919eac6ebceed2cf0d0f26ff528f8f5fa84fdf2ff4302;
    inBuf[3788] = 256'h510484061509e60b360fe1126416cb19e21c501f6c213c239124e9254c278f28;
    inBuf[3789] = 256'h302a142ce32de82fc93112331634963461340f349133d232603200326b31ff30;
    inBuf[3790] = 256'h5e30492f352ef02c762b622a9e293629a829b42a392c702ee830683313368038;
    inBuf[3791] = 256'h9c3aa63c6b3e0e40e341b5438e45844733499a4acb4b804cdc4cf84c8f4ccb4b;
    inBuf[3792] = 256'hcb4a5b49c44722462744f6417e3f5f3cd538f7348b30ec2b352727221f1d3e18;
    inBuf[3793] = 256'h47139d0e480ae905c101bffd85f96ef593f1c3ed77eac3e75ae57ce304e288e0;
    inBuf[3794] = 256'h45df30de10dd3ddcaedb29dbf4da02db29dba8db5ddc02dda6dd11de1ede04de;
    inBuf[3795] = 256'hc9dd74dd2dddd9dc66dce1db3edb93daf3d95ad9cad82ad865d784d670d53bd4;
    inBuf[3796] = 256'h14d3ead1e8d041d0cbcfa5cfeccf55d002d110d236d3a5d480d670d8abda50dd;
    inBuf[3797] = 256'hfedff1e23fe67de9dfec7ef0f3f389f769fb35ff35038207a80be00f37144518;
    inBuf[3798] = 256'h4c1c692042241028de2b3c2f4a3208352337da38593a763b763c6c3d163e973e;
    inBuf[3799] = 256'hf73e0e3f1c3f393f463f663f843f7a3f6c3f513f1a3fe33e7a3ec13dd73caf3b;
    inBuf[3800] = 256'h783a8939c7383538d4373c377336ad35c234f1336a33c832143259313130db2e;
    inBuf[3801] = 256'h8c2df42b5a2ae02820275e25b523c021ca1fed1dc81bab199e173315b2122410;
    inBuf[3802] = 256'h420d7f0afa0767050d03d10056fef8fbccf9adf7ecf560f49ef2c1f0b2ee61ec;
    inBuf[3803] = 256'h3fea65e8b8e656e506e493e225e1bedf6bde61dd96dcfadb9bdb64db4edb5fdb;
    inBuf[3804] = 256'h80dba7dbccdbe6db00dc1edc40dc74dcb1dcf0dc44dda2dd00de70dedade3bdf;
    inBuf[3805] = 256'hb5df41e0dee0abe182e249e317e4d4e47ce543e611e7d0e79fe863e918ea0eeb;
    inBuf[3806] = 256'h4aecc8edb4efd7f1f3f323f646f846fa65fc89fe830077023e04b10516076208;
    inBuf[3807] = 256'h78098d0a820b2b0cc10c430d980d000e740ec30e110f490f360ff70e8d0ed70d;
    inBuf[3808] = 256'h040d320c430b580a800987087e0786067b0572048e03960289018f0081ff6dfe;
    inBuf[3809] = 256'h8cfd9ffc91fb82fa30f9a1f724f699f40df3bef16cf013eff1edd3ecc7eb0deb;
    inBuf[3810] = 256'h64eacce971e909e995e83ee8b7e70ae763e685e592e4b9e3bae2ade1aee079df;
    inBuf[3811] = 256'h33de05ddb7db7bda77d978d8b7d75ad727d73dd791d7bdd7c9d7b8d75cd7fcd6;
    inBuf[3812] = 256'hc5d68ad671d674d64ad61dd606d6d9d5c6d5cbd59fd567d533d5e4d4c6d4edd4;
    inBuf[3813] = 256'h1ed57cd5fad55dd6e7d6a6d766d85fd97fda82dbabdcfcdd3cdfa7e01ee246e3;
    inBuf[3814] = 256'h58e449e5ece5a7e681e744e843e96cea7cebb4ecf0edd9eea7ef48f09af006f1;
    inBuf[3815] = 256'ha0f14bf241f35bf44ef53af6fbf66cf7b4f7bff77af715f794f60af6a9f563f5;
    inBuf[3816] = 256'h32f515f5d8f479f4fef349f382f2bcf1e2f028f09aef12efc0eea3ee86eea5ee;
    inBuf[3817] = 256'h01ef63ef09f0f2f0e7f13cf314f549f730fabbfd700154052a09800c9e0f9d12;
    inBuf[3818] = 256'h50151718f81aa11d65204b23192628295a2c2f2fc531dc3326352636fb369937;
    inBuf[3819] = 256'h82388b39593a3b3be93b1b3c3c3c003c1b3bfb396838583692341133db317d31;
    inBuf[3820] = 256'h88319831f2311a32df31d831d531e03190329733dc34c536e838223bbb3d3d40;
    inBuf[3821] = 256'h7d42b7448b460b489e49154b974c604e005064518c520353e35257522051884f;
    inBuf[3822] = 256'hc04d814b1b49ad46eb432441643e3c3be6374f3405305e2b76261621cc1bc716;
    inBuf[3823] = 256'hc411260de908a104a300edfc28f9aef578f228ef12ec3be96ae610e43fe2b6e0;
    inBuf[3824] = 256'hb8df24dfa9de84dea5ded9de61df18e0bce078e12ae2b0e246e3cde322e460e4;
    inBuf[3825] = 256'h53e4e2e334e339e2fee0b5df53dee4dc80db15daa2d82cd7a4d51cd49ad227d1;
    inBuf[3826] = 256'hdacf9fce74cd68cc64cb8dca17cae8c91fcacbcaa3cbc1cc4fce21d077d27ad5;
    inBuf[3827] = 256'hced883dc9de0aae4d0e832ed72f1c1f542fa93feec027e07f10b78103215b519;
    inBuf[3828] = 256'h241e9822b4269d2a652ead318b340c37e8384c3a5b3bf03b413c693c3f3cea3b;
    inBuf[3829] = 256'h6d3ba53abc39bd38a1379c36ab35be34f9333e338432f5317231f7309e303430;
    inBuf[3830] = 256'hbd2f672f152fed2e1e2f6c2fde2f803002317d310d326e32c03211331233ef32;
    inBuf[3831] = 256'hc2324832c031363157305a2f442ec12c122b3629dd265524a8219a1e851b6218;
    inBuf[3832] = 256'hda142b113f0dd8085f04e7ff4efbf5f6d0f2a4eec0ea14e77be341e054dd8dda;
    inBuf[3833] = 256'h2ed822d650d4f8d2fdd148d100d1fbd026d19dd130d2d8d2b4d3a2d4b3d500d7;
    inBuf[3834] = 256'h53d8aed90edb3ddc5cdd89dea0dfbbe0c8e179e2dce2f6e2ade24ce2eae15ee1;
    inBuf[3835] = 256'hcde02ce04ddf6cde92dd99dcb2dbc2da92d95fd82dd7f6d518d596d457d49ad4;
    inBuf[3836] = 256'h43d528d683d72cd9efdafedc22df24e14ae370e57ae7c6e942eccbeeadf1b0f4;
    inBuf[3837] = 256'h8df77afa47fdc5ff5602ec045807df09510c5a0e3110bb11b7126513ac133d13;
    inBuf[3838] = 256'h5212fb101a0f180d260b1d09330774059d03da014800adfe1cfd9ffbe7f90bf8;
    inBuf[3839] = 256'h38f651f484f200f18bef2aeef5ecb6eb81ea83e98ce8b5e728e7bce699e6ede6;
    inBuf[3840] = 256'h7ce744e83fe90ceaabea32eb65eb72eb7deb47ebfceac2ea5beafce9bfe94be9;
    inBuf[3841] = 256'hbae817e80ce7d4e5a2e439e3dde1b5e06bdf2dde1adddcdba7da9cd965d833d7;
    inBuf[3842] = 256'h28d6f5d4d9d3fcd210d24dd1cdd03dd0cecf9ccf5bcf43cf6dcf8ccfe0cf7ed0;
    inBuf[3843] = 256'h18d1eed106d306d425d55cd655d755d85cd91fdaf6daeadbb4dca7ddbcde8bdf;
    inBuf[3844] = 256'h55e005e141e16ce194e178e17ce19ce184e184e19be17fe187e1b4e1bce1ebe1;
    inBuf[3845] = 256'h3ee279e2e1e273e3f2e395e450e5ece599e643e7bce725e867e871e872e861e8;
    inBuf[3846] = 256'h42e83fe83ce83ee85ee870e87fe89ce895e88ae8a2e8b6e8fbe889e915eab7ea;
    inBuf[3847] = 256'h78eb0decb3ec98ed85eec0ef6cf13ff37df541f830fb74fefc0148057308830b;
    inBuf[3848] = 256'h290ec0107113fb15ad18901b4c1e28211b24c1264829882b1e2d612e572fe52f;
    inBuf[3849] = 256'h9330623116320433f73399344135ac358e354435983468334c3239312230872f;
    inBuf[3850] = 256'h1f2fa42e6f2e2f2ebe2d902d6d2d3f2d7f2dfc2dae2e0630b2318033a335af37;
    inBuf[3851] = 256'h8439723b3d3dec3ec4407342f3437c45c846ee471e49014a9c4afd4acb4a2d4a;
    inBuf[3852] = 256'h4849d74715461d44a341f13e203cea3897352a32452e302af5254f21ac1c2618;
    inBuf[3853] = 256'h7b130f0feb0ab806cd0221ff53fbb3f73af49cf044ed45ea64e7ffe416e35fe1;
    inBuf[3854] = 256'h24e062dfd2deabdecaded5deebdefbdedadecedee7de07df54dfbcdf17e079e0;
    inBuf[3855] = 256'hd8e019e141e142e106e19ae00de06ddfc6de25de83ddcbdc05dc38db56da77d9;
    inBuf[3856] = 256'hadd8ded72bd7b0d64fd637d680d6f1d6add7c8d8ffd983db6bdd6ddfbae166e4;
    inBuf[3857] = 256'h1ce713ea63edaaf01df4ccf754fbf3fec5026706170ae80d7411fd14a518121c;
    inBuf[3858] = 256'h901f3723a626172a962dc030c433a236f638eb3a8b3c983d663e153f793fd23f;
    inBuf[3859] = 256'h19401640fc3fc43f5a3ffa3e963e103e973d0c3d673ce73b6c3bf73aaa3a423a;
    inBuf[3860] = 256'hb93933396e3881379e3685355c345e334e326031c1301630812f192f7c2edd2d;
    inBuf[3861] = 256'h5b2d9a2cd32b232b2f2a3d296f2865275c265725e8235222a420881e531c141a;
    inBuf[3862] = 256'h7217c1140f12190f3e0c82099406b703dc00b8fda2faa6f793f4c3f133efa5ec;
    inBuf[3863] = 256'h60ea53e843e66ce4b7e2efe04edfd0dd5adc36db65daccd995d9a3d9c4d905da;
    inBuf[3864] = 256'h3bda43da30daf9d9a1d957d926d91cd94dd9abd930dad6da80db31dce2dc7fdd;
    inBuf[3865] = 256'h1ddebfde63df2be00fe1f8e1f7e2e6e3a4e451e5d7e52ce686e6dae624e7a7e7;
    inBuf[3866] = 256'h56e824e942ea83ebb9ec0fee5bef81f0c2f103f323f466f5b4f6f7f778f91efb;
    inBuf[3867] = 256'hb5fc6bfe10006d01c5020e042205400656072b08fd08c909630a030b9d0be00b;
    inBuf[3868] = 256'hed0bc30b2d0b670a92098108620753062205f9030003f901f6000700e1fe94fd;
    inBuf[3869] = 256'h4afcd9fa64f924f8e8f6baf5bff4b8f3a8f2b2f19cf072ef64ee45ed2eec59eb;
    inBuf[3870] = 256'h9dea0fead4e9afe9a6e9cae9d0e9bce9a7e94fe9d5e868e8dae756e700e791e6;
    inBuf[3871] = 256'h20e6c4e52de582e4e4e308e31ce240e12ee020df41de4add6adcbadbe0da0ada;
    inBuf[3872] = 256'h5bd985d8bdd722d75fd6afd538d5b6d471d483d49bd4e9d467d5b5d503d653d6;
    inBuf[3873] = 256'h55d64ed64dd618d607d62cd64bd6b4d65fd7fcd7d1d8c7d988da5edb31dcb5dc;
    inBuf[3874] = 256'h47dddedd43dedcdea3df59e053e173e267e373e477e52ee6f2e6bfe76ae84be9;
    inBuf[3875] = 256'h4dea34eb39ec34ede7ed88eef3ee01efeaeea5ee31eed6ed8aed52ed54ed5ded;
    inBuf[3876] = 256'h5eed69ed49ed0eeddaec87ec43ec37ec33ec72ec13edcfedd3ee20f04ff18ff2;
    inBuf[3877] = 256'hedf31cf580f646f82bfa8dfc77ff7d02e1059809220dbb10511470176a1a531d;
    inBuf[3878] = 256'he81fa32299257328822b9f2e4c31c633e035443760382f398c39013a7c3ac33a;
    inBuf[3879] = 256'h443bc43bfa3b493c673c133cc13b343b523ab2392339893860384538ff37f537;
    inBuf[3880] = 256'hca3757371637bb3639361f3637368f36a9372d39f43a393d733f71416f430f45;
    inBuf[3881] = 256'h5e46ba47e8480e4a724bb74cde4df64e884fa44f684f844e414dcd4be349db47;
    inBuf[3882] = 256'hd1456e430141823e803b4038b93484300f2c682741221c1d0d18c712ca0d2009;
    inBuf[3883] = 256'h69040e0006fce4f709f474f0cdec80e999e6c9e373e194dfd5dd7bdc79db80da;
    inBuf[3884] = 256'hd1d96dd91ed923d971d9ccd955daf4da74dbf7db74dcd0dc27dd6cdd8add96dd;
    inBuf[3885] = 256'h8cdd6cdd4fdd31dd14ddfbdcdddcc0dc9fdc77dc4adcffdb91db0edb65dab1d9;
    inBuf[3886] = 256'h16d985d81dd8fdd7ffd747d8f3d8c9d9e9da6fdc18de0de073e2fde4d2e706eb;
    inBuf[3887] = 256'h34ee80f102f555f8a5fb14ff44027205d008110c720f1a13a216311ae01d5421;
    inBuf[3888] = 256'hbb243328602b5e2e39319f33b835a2372a39803ab93ba53c6a3d0f3e693e993e;
    inBuf[3889] = 256'h963e443ec33d0d3d203c243b053ac2387a370d368d342433b3315a30372f0e2e;
    inBuf[3890] = 256'hf42cfa2bd92ab229a428762760268525a224e22350239422d9212a213f20561f;
    inBuf[3891] = 256'h851e841d961cc31bbf1ac219c618761713169214b512d010e00ea50c6e0a2a08;
    inBuf[3892] = 256'h990511038500bcfd0bfb52f859f579f2a7efc2ec2beac8e763e536e311e1c6de;
    inBuf[3893] = 256'h9edc80da57d86bd69fd4e9d28cd16fd090cf1dcfe0cec8cee5cefcce0dcf2dcf;
    inBuf[3894] = 256'h27cf15cf18cf0acf21cf78cfe0cf81d056d11cd201d3ffd3d8d4c2d5b9d687d7;
    inBuf[3895] = 256'h7ad893d99ddad5db11ddfbddc9de65dfa9df00e066e0aee020e196e1d4e12fe2;
    inBuf[3896] = 256'h99e2eae27be32fe4cce4a1e591e669e779e8a0e9a0eabfebdfeccbedd1eed7ef;
    inBuf[3897] = 256'ha9f098f199f284f3b4f41ef686f721f9c8fa2dfc81fdb0fe7eff2c00bc00fe00;
    inBuf[3898] = 256'h3c0183019501a2019b0132019600dbffd4fec8fdd2fcb3fb8ffa73f916f89bf6;
    inBuf[3899] = 256'h1cf55bf383f1c5effaed5bec18ebf6e903e94de883e7b8e60de649e589e4f6e3;
    inBuf[3900] = 256'h5ce3e3e2bae2abe2d2e241e3a0e300e47ce4cfe41ee586e5b5e5c8e5dfe5b7e5;
    inBuf[3901] = 256'h8ce58fe56be540e51be597e4e2e32de330e22be147e02cdf12de25dd19dc32db;
    inBuf[3902] = 256'h91dad0d91dd985d8a6d7c4d6fdd503d524d474d3a0d2fdd199d125d1f7d011d1;
    inBuf[3903] = 256'h1cd166d1ead14ad2d7d283d3f9d39ad46cd52ed644d7a5d8f5d973dbf9dc30de;
    inBuf[3904] = 256'h68df9ce09be1c8e21ee46be5f3e68fe8f6e94beb5aece9ec30ed1fedb7ec4cec;
    inBuf[3905] = 256'hd6eb59eb0aebb9ea58eaffe974e9b8e8f0e7eee6dbe5eee404e45ae328e338e3;
    inBuf[3906] = 256'hbee3c6e4f0e54fe7dee83feab8eb7aed55efb7f1c9f432f827fc9200e3043f09;
    inBuf[3907] = 256'h930d72113515fa187c1c27200b24c527a02b7d2fe032fe35ac38813ad73baf3c;
    inBuf[3908] = 256'he53c0b3d2b3d173d363d4e3d053db13c083ccc3a7539d537de353834ca328b31;
    inBuf[3909] = 256'h0c31f230f7307531f5313932bb322c337a333d343935603632384e3a803c143f;
    inBuf[3910] = 256'h9141c7430346e7476c49f24a3d4c6c4ddf4e4b50b15128532b54aa54b954fd53;
    inBuf[3911] = 256'hb7522b511f4fe94cbc4a3e48ad450f43eb3f743cb4384d34ab2ffe2a01262021;
    inBuf[3912] = 256'h791caa171013be0e520a290652026cfed4fa9ff776f4b2f15def1aed31ebb4e9;
    inBuf[3913] = 256'h59e86ee700e7b8e6bde602e735e78ae70be87ee80ee9b3e930eaaaea29eb8aeb;
    inBuf[3914] = 256'hf0eb4aec66ec4aeceeeb42eb6aea71e949e801e797e50fe489e21be1cfdfa4de;
    inBuf[3915] = 256'h8cdd75dc53db34da2bd940d894d73cd72ed78bd75dd873d9d3da68dcefdd8edf;
    inBuf[3916] = 256'h68e162e3c7e5b6e8e0eb65ef45f319f7fffafffead023406b609e90c1b108313;
    inBuf[3917] = 256'hc916161a771d80205623152668287a2a5b2cbf2dd72ec92f6f300c31b6313e32;
    inBuf[3918] = 256'hcf326233cc333334803488346c3415347933dc3230327231d33020304e2f8e2e;
    inBuf[3919] = 256'hb92dd92c252c692bab2a1a2a8229f728a92858280d28e727a52767275b274a27;
    inBuf[3920] = 256'h4f277a27752750271f27a7261e26ad252025a3244324ab23f4221722c520301f;
    inBuf[3921] = 256'h761d6d1b681980177a1584138d11490fe40c5e0a820792049d0178fe70fb95f8;
    inBuf[3922] = 256'hbbf522f3c2f063ee35ec36ea3be87de6ffe49de38ae2c7e13fe11ce153e1c0e1;
    inBuf[3923] = 256'h66e222e3d1e37fe421e5bbe567e61be7e8e7dbe8dde9fcea2bec37ed24eee1ee;
    inBuf[3924] = 256'h45ef7def97ef7def67ef58ef2aef0eeffdeec7ee96ee5ceee6ed69edf0ec69ec;
    inBuf[3925] = 256'h1eec18ec2fec83ecf2ec39ed78eda0ed94ed94eda6edb1edebed46ee9bee14ef;
    inBuf[3926] = 256'ha4ef24f0c6f080f126f2e7f2b5f35cf40cf5c0f54ff6f3f6b5f76bf844f93dfa;
    inBuf[3927] = 256'h13fbe2fbaafc2bfd91fdf5fd26fe51fe8dfe9bfe92fe7dfe14fe6ffda4fc7cfb;
    inBuf[3928] = 256'h24fac3f82bf784f5ebf328f261f0bcee0ded89eb51ea2ae92be85de774e68be5;
    inBuf[3929] = 256'hbae4cde3f3e256e2c3e168e161e168e194e1ece11ee24be28ce2b7e20be3b3e3;
    inBuf[3930] = 256'h7ce48ce5dee614e834e930eab5eaefeaf9eaa8ea44eaece962e9d3e845e86ae7;
    inBuf[3931] = 256'h7ae692e57be47ae3a4e2aae1bee0e7dfdcdee3dd17dd39dc8ddb21dba6da5dda;
    inBuf[3932] = 256'h50da35da51daa9daedda61db04dc86dc27dddedd53decade46df84dfe4df74e0;
    inBuf[3933] = 256'hf0e0a6e188e23de303e4cee44ee5cee553e6a0e604e783e7d7e72fe873e85ce8;
    inBuf[3934] = 256'h19e8b1e713e78ee63ce613e640e6a4e60ee770e786e72be772e654e509e4e9e2;
    inBuf[3935] = 256'hfde173e162e17de1bce119e24be27ce2dde24de319e47de54be7b6e9d4ec43f0;
    inBuf[3936] = 256'h05f408f8dcfb86ff0203ff05bc08740b100ef8105b14f717e51bfc1fb9232427;
    inBuf[3937] = 256'h1f2a622c392ebd2fcf30d631df32b6339b345b3593356d35bf346433e6316830;
    inBuf[3938] = 256'hfb2e262ec92da02ddd2d212e1b2e132ecc2d2a2dac2c3e2cf42b5a2c4a2da52e;
    inBuf[3939] = 256'ha430cb32c934cd368138e339663be13c693e554057425c4488466548d749ec4a;
    inBuf[3940] = 256'h404be54a164aa348db460745f642ec40063fe43cb03a62388b356332f92e0c2b;
    inBuf[3941] = 256'h0f273723511fc31b8b183415ea118e0eb20aae06a3026bfe8afa32f72ff4d1f1;
    inBuf[3942] = 256'h0bf06fee17ede0eb76ea1ae9e4e7bee6fee5b2e5a5e5f3e576e6e3e64fe7aae7;
    inBuf[3943] = 256'hd5e702e83ae86ae8bae81be969e9b2e9dde9c8e97be9e9e800e8d4e675e5f6e3;
    inBuf[3944] = 256'h74e208e1b4df68de20ddd6db7bda2bd903d8f5d619d682d511d5e7d430d5ced5;
    inBuf[3945] = 256'hd7d65bd808dad8dbe0ddecdf25e2cee4bae700ebc2eea0f290f6a2fa78fe2002;
    inBuf[3946] = 256'hd3055f09f20ccd10a6147918471c981f542290240a26ee268727be27c227c127;
    inBuf[3947] = 256'h83270d276c2671253524df226221e61f841e2e1dfd1bfb1a1a1a6719cc182e18;
    inBuf[3948] = 256'h9517f2165216e01591156d157f159a15c9152a16ab166c177c18a219d71a0e1c;
    inBuf[3949] = 256'h121df91dc71e4d1f9c1faa1f4d1fb61ef81d001d021cf81aba197c184217f215;
    inBuf[3950] = 256'hbd148213f3112310f40d4f0b9908f4055d031301f5feb8fc76fa14f86ff5cdf2;
    inBuf[3951] = 256'h3af0b0ed75eb98e905e8e5e61ee67ce506e59ee42fe4e2e3c0e3d1e33ce4efe4;
    inBuf[3952] = 256'he1e513e74ee877e990ea76eb32ece5ec7eed14eebfee5ceff9efa3f032f1aff1;
    inBuf[3953] = 256'h17f232f20af2a5f1e4f0f3efedeeb6ed79ec43ebf5e9c2e8b6e7aee6cfe513e5;
    inBuf[3954] = 256'h49e4a3e32ee3cde2bbe2f1e232e39ee324e496e433e509e6f8e636e8bbe94deb;
    inBuf[3955] = 256'h0eede7ee9ff057f2fff369f5c9f624f861f9b9fa2afc80fdccfee9ff9000d300;
    inBuf[3956] = 256'ha900f4ffedfeb1fd35fcb8fa52f9e7f79bf66cf527f4dff29bf13ff0f9eeefed;
    inBuf[3957] = 256'h09ed61ecfbeb9feb53eb1eebdaea9fea7fea54ea2eea1dea05ea09ea48eaaaea;
    inBuf[3958] = 256'h4aeb26ec07edf5ede9eeb4ef7bf04bf104f2ccf2a4f34ff4e4f45bf579f569f5;
    inBuf[3959] = 256'h3bf5c8f447f4d5f344f3c6f26ff204f2a4f152f1c4f018f063ef74ee79ed92ec;
    inBuf[3960] = 256'h86eb73ea69e928e8d1e681e50be4a9e28fe1a5e027e02fe06fe0e2e065e18ee1;
    inBuf[3961] = 256'h76e13be1c5e075e083e0c4e06de184e2abe3fae462e67be769e83ae9b6e93dea;
    inBuf[3962] = 256'h04ebd2ebe1ec28ee36ef21f0e0f015f1ecf072f062ef02ee81ecceea45e913e8;
    inBuf[3963] = 256'hfee61de64fe53ee4f9e27fe1bbdfefdd3ddcb0da89d9c8d85ad841d83ed82cd8;
    inBuf[3964] = 256'h12d8d2d794d79ad7e2d7a4d803dac7dbfedda1e050e315e6f5e8a6eb68ee6af1;
    inBuf[3965] = 256'h71f4b4f73ffba3fefa014a053508f90aba0d2a108e120b155417b219361c7f1e;
    inBuf[3966] = 256'hb520cb225b24a725ba265b27e6276a28ad28052965298129a529ae2956290729;
    inBuf[3967] = 256'hb8284c2848289428f328c529c42aa22bc02cdd2dbb2ed02fed30f2316e333e35;
    inBuf[3968] = 256'h3b37cc39903c313fed415b44464617489949d14a3b4ca14dfa4e8b50df51cd52;
    inBuf[3969] = 256'h7d538853ff523e521051b14f704efd4c744bf1490148b9452a43e93f323c3a38;
    inBuf[3970] = 256'hc5333e2fe12a6f264e229c1eff1ac217dc14d211df0e050cf7083006e003ca01;
    inBuf[3971] = 256'h45003eff32fe4efd82fc71fb6bfa7bf956f84af76ff695f509f5d3f49af46df4;
    inBuf[3972] = 256'h2cf488f3adf2b1f17bf03beffeedaaec69eb49ea32e92be81ce7d6e559e4b5e2;
    inBuf[3973] = 256'hfde060dffbddcedcdadb1bdb8bda29dafcd9f5d9f7d902da21da5bdae1dacadb;
    inBuf[3974] = 256'hf0dc47deb6dffde036e287e3dfe473e666e87beac7ec61effff1b3f48df736fa;
    inBuf[3975] = 256'hc2fc5cffcb013c04e9068509190cbc0e1a1145136d155c172c19071bb21c431e;
    inBuf[3976] = 256'he21f6121d52250249825b526a8274828b028ec28ee28e928e928e128ef28f628;
    inBuf[3977] = 256'hc7286828ad278d264d25fa23b722cd212121ab2085207420622067204020e81f;
    inBuf[3978] = 256'h881ffb1e5e1eef1d8b1d421d411d4c1d701dcb1d181e591ea61ebd1eb71ec71e;
    inBuf[3979] = 256'hba1ea01e821e0d1e451d411cd81a3c19a317e31520147412af10f60e670dcd0b;
    inBuf[3980] = 256'h490aed08830737061e050004fb0210020301f3ffecfebffd8ffc67fb21faedf8;
    inBuf[3981] = 256'hedf70ef780f64ef649f678f6ccf61ef781f7f3f754f8b3f803f933f956f961f9;
    inBuf[3982] = 256'h4cf924f9d2f855f8cbf72bf78ef616f6acf55df539f51af508f509f5e1f493f4;
    inBuf[3983] = 256'h25f46ff39cf2ddf11ef185f01ef0aaef35efcbee43eecfed8fed58ed42ed52ed;
    inBuf[3984] = 256'h47ed40ed5ded6bed8dedc9eddeede9edf9ede0edcbedd2edbeedaaeda1ed64ed;
    inBuf[3985] = 256'h15edc5ec42ecb7eb47ebc8ea6aea47ea22ea0aeaffe9b7e951e9e6e847e8a7e7;
    inBuf[3986] = 256'h20e776e6cae527e555e486e3d7e21ae287e136e1e1e0afe0a8e086e078e096e0;
    inBuf[3987] = 256'ha2e0d5e041e1a4e12ae2dae264e3f6e3a0e426e5c7e5a2e679e77be89de985ea;
    inBuf[3988] = 256'h4febfbeb54eca4ec0bed54edaced07ee10eef0eda6edf4ec1cec2bebe9e99fe8;
    inBuf[3989] = 256'h66e712e6f6e425e460e3dce29be255e243e26ce285e2bde215e33ce366e3a7e3;
    inBuf[3990] = 256'hc4e3fae357e49ae4f5e473e5cfe53de6c6e628e79ee737e8bfe873e950ea05eb;
    inBuf[3991] = 256'hbceb68ecc5ec19ed72ed99edceed09eef9edd0ed8aedefec46eca1ebd1ea1cea;
    inBuf[3992] = 256'h8fe9f9e893e85de814e8cce771e7d4e617e640e53ce42fe315e2e6e0c8dfc0de;
    inBuf[3993] = 256'he4dd5add06dde7dc04dd31dd89dd35de13df3fe0bee136e3b3e446e6bce758e9;
    inBuf[3994] = 256'h4ceb54ed90ef0df275f4fcf6c9f99efcbcff2f0392060a0a960dd9100b143217;
    inBuf[3995] = 256'hfc19aa1c431f7e21b023d62598273c29ad2a962b532ce12cff2c1a2d2b2df32c;
    inBuf[3996] = 256'he12ce32cb72cc62ce92cd22ce42cf92cd62cf32c2f2d592de52dae2e872fe530;
    inBuf[3997] = 256'h9a327734cd363c39783bc53dd13f8a4168433c450b473649614b5e4d5b4fd750;
    inBuf[3998] = 256'hb0512952f1512d514550fd4e824d1f4c784aa848e146bb445a42e73fef3caf39;
    inBuf[3999] = 256'h6a36dc32662f462c22293b26a023d7201b1e7a1b861886159112510f300c6109;
    inBuf[4000] = 256'ha60660049e02f900a2ff95fe74fd84fcd9fb30fbc9faa2fa70fa5dfa5cfa29fa;
    inBuf[4001] = 256'heef99df9fff841f855f718f6cef485f337f227f14af078efbaeee4edc6ec7feb;
    inBuf[4002] = 256'h0eea71e8d5e637e586e3d4e113e03ede76dcc0da22d9b3d77fd68ed5e7d491d4;
    inBuf[4003] = 256'h8cd4c5d438d5edd5ddd61ed8c7d9afdbbfddeddf02e2fde30de621e83bea73ec;
    inBuf[4004] = 256'h92ee90f09ef2b0f4eaf687f955fc3bff4a023505e5077c0ab80c7d0ef10fed10;
    inBuf[4005] = 256'h8811151294121413b9133f147c1484142f147f13b712e4112311ab107c109810;
    inBuf[4006] = 256'h051194111e129812e6120313fe12dc12a0124412d0114b11b11015108a0ff50e;
    inBuf[4007] = 256'h500e9f0dc70ce30b1f0b8c0a500a860a040ba60b400c8c0c7a0c030c170bec09;
    inBuf[4008] = 256'ha30846070d060b053f04ca03a903bc0303045a049904c604cf04b104a1049f04;
    inBuf[4009] = 256'ha604c704d504a60436045903fe014f004ffe1dfc07fa24f887f65cf598f42df4;
    inBuf[4010] = 256'h23f44ff497f4f2f427f51bf5d2f42ef440f335f20cf1e0efdeee08ee74ed3aed;
    inBuf[4011] = 256'h38ed58ed8aeda0eda4edb9ede9ed4eeef1eea9ef67f01df1a1f105f255f265f2;
    inBuf[4012] = 256'h47f2fdf164f1aff0f8ef3befa1ee3deef9edf9ed49eebfee5eeff8ef3bf03af0;
    inBuf[4013] = 256'h06f09bef42ef13efe2eec8eeb3ee72ee44ee41ee41ee6deebceef2ee43efc1ef;
    inBuf[4014] = 256'h49f013f113f2f6f2d0f391f4f7f434f555f51bf5b0f424f443f34cf263f166f0;
    inBuf[4015] = 256'h84efd2ee1cee87ed29edd4ecafecd4ec19ed97ed54ee11efcdef74f0c2f0c4f0;
    inBuf[4016] = 256'h85f0ebef20ef46ee52ed79ecd7eb55eb1deb25eb34eb57eb6deb3aebfceacfea;
    inBuf[4017] = 256'ha5ead2ea5debf0eba2ec5aedbdedf4ed0deec4ed56ede4ec40ecc0eb96eb8eeb;
    inBuf[4018] = 256'he8ebbeecbded02ef86f0cef1d5f28ff398f318f34cf214f1bcef80ee32edfaeb;
    inBuf[4019] = 256'hf4eaefe918e97ae8d8e767e72fe7f8e6fee64ce796e70be8a9e813e962e9c1e9;
    inBuf[4020] = 256'hb9e97de94de9c4e846e8fce79de767e76ae766e7a1e726e8b2e867e922ea86ea;
    inBuf[4021] = 256'hbfead8eab2eaafeae9ea29eb8aebefeb0aecebeb8eebe0ea0fea24e91ce81de7;
    inBuf[4022] = 256'h23e633e56ae4b4e31ee3c9e297e29fe2efe24ce3b8e337e4a0e42ce509e617e7;
    inBuf[4023] = 256'h91e884ea9becf4ee9af147f42cf758fa7cfdb800ff030007f009de0c950f5f12;
    inBuf[4024] = 256'h4515fd17b91a631da81fc321a82324259226f3271b29652ab42bce2c082e392f;
    inBuf[4025] = 256'h1c300d31d9313432823298324132f831a3311d31ef30ed30db3028318d31c131;
    inBuf[4026] = 256'h3f32d3324d33353453356c36fc37b239433b0e3dab3ece3fea40ca416c427c43;
    inBuf[4027] = 256'hca443d4645485f4a3b4c304ebf4fb9509151d05153519a50484f654d8b4b7149;
    inBuf[4028] = 256'hfd46a844fc41d13eae3b3b388c342531a22d212a242738247a21511f1e1dc41a;
    inBuf[4029] = 256'h7f18bb159312870f500c3209a40643042902a60048ff1afe4bfd69fc85fbd9fa;
    inBuf[4030] = 256'h1ffa91f970f969f98cf9ebf923fa47fa6efa49faf6f987f9c8f8f4f741f795f6;
    inBuf[4031] = 256'h28f608f6ebf5d0f59ff513f53ff42df3bff11ff066ee8cecbeea14e98ce751e6;
    inBuf[4032] = 256'h75e5e7e4a7e4a8e4bde4d2e4f8e442e5c3e59ee6dce758e9feeac6ec93ee79f0;
    inBuf[4033] = 256'h94f2cef427f795f9dbfb02fe2500220218042a062508120a140cf70dc50fa211;
    inBuf[4034] = 256'h5c13f3148116d017dd18be19471a781a651aee1926192a180617e515d814da13;
    inBuf[4035] = 256'hfe12251241117f10cc0f100f5a0e730d4e0c2f0b1f0a4209e108d708fe082209;
    inBuf[4036] = 256'h0d09a808fe072c075106b80553052f05860537064107d408c20ad40cf30ed210;
    inBuf[4037] = 256'h46125613e9130a14df136613c01222128f111911cc1081103510f10fa40f5c0f;
    inBuf[4038] = 256'h2b0ff20ea80e3e0e890d820c2a0b76098b078905770376018cffadfdfefb8dfa;
    inBuf[4039] = 256'h49f942f86cf7a5f6f3f55bf5edf4cef4fcf46af511f6b4f62cf78cf7d8f725f8;
    inBuf[4040] = 256'habf864f93cfa27fbf3fb91fc13fd6afd9cfdb8fda0fd5ffd0dfd99fc32fcfffb;
    inBuf[4041] = 256'hd8fbc2fbb3fb60fbc6fae1f974f8a6f6aaf476f263f0ccee9bede2ec91ec35ec;
    inBuf[4042] = 256'hb4eb12eb24ea32e979e8d2e75ae724e7ebe6c9e6dfe6f4e615e746e73be7f6e6;
    inBuf[4043] = 256'h8fe6efe559e504e5dfe41be5c0e579e63de7ebe733e841e83de807e8e2e7f4e7;
    inBuf[4044] = 256'h07e831e867e85ee841e82ae8dce775e703e763e6dbe589e53be51de52ce51de5;
    inBuf[4045] = 256'h0de5fce4b3e459e4e2e319e34ae293e1dfe086e08de0a7e0f0e04ee188e1e8e1;
    inBuf[4046] = 256'h7be217e3fee318e510e61ce739e821e91bea27ebf6ebbfec8eed28eed3eeaaef;
    inBuf[4047] = 256'h7af07bf1aef2c5f3dff4f0f5aaf635f79bf79ef769f700f727f60ef5bff313f2;
    inBuf[4048] = 256'h54f09deec0ecfeea6be9d8e77ce671e594e426e422e43ae489e4fae435e560e5;
    inBuf[4049] = 256'h84e56ae54de53de511e516e56de5ede5cbe607e856e9c5ea43ec8cedb6eeb1ef;
    inBuf[4050] = 256'h44f096f0b3f08af05ff045f01bf0f7efbeef3def99eee2ed12ed50ec96ebc1ea;
    inBuf[4051] = 256'he4e9fce813e858e7d6e69ae6b4e606e77de70ee897e824e9c9e96aea1eebf1eb;
    inBuf[4052] = 256'hbeeca2eda7eeaeeff8f0abf2a1f4f9f6a2f937fcb5fe10010503cd0488060b08;
    inBuf[4053] = 256'h9c095b0b120df00e08111a134a159417b219c21bac1d251f50201a215b217621;
    inBuf[4054] = 256'h9121ad212222d22277233924e0244a25d9257426ea267d27e727ec27e927cd27;
    inBuf[4055] = 256'h9d27d5274d28d428b129972a582b492c332df42dda2eac2f56302f310a32df32;
    inBuf[4056] = 256'hf83310351b36583783389c39e03af93bd53c943ddf3dbd3d623d8a3c583b0d3a;
    inBuf[4057] = 256'h67388e36bb34a8327730482ec12b042941263e234020811dbe1a2c18e815a313;
    inBuf[4058] = 256'h9311d50f150e8b0c500b0b0ae208da07990658053804f802e20116014c00aaff;
    inBuf[4059] = 256'h30ff80febdfd04fd2afc70fbf0fa6cfafcf99bf90af95ff8a6f7c6f6eaf518f5;
    inBuf[4060] = 256'h39f476f3d1f22cf29cf112f17ff0faef7fef04ef9aee24ee88edd4ec05ec38eb;
    inBuf[4061] = 256'haaea73ea99ea16ebbbeb5aecdbec30ed6ceda4ede1ed2aee6beea5eef2ee59ef;
    inBuf[4062] = 256'hf7efe7f004f22af346f421f5b6f530f68df6edf695f781f8b8f955fb21fdf0fe;
    inBuf[4063] = 256'hae000d02ee027303980375034a031803ed02f80225036903d5034b04b6041e05;
    inBuf[4064] = 256'h68058e05a805a80582054405dd045a04db035f03e902900247020f02fd010e02;
    inBuf[4065] = 256'h39028602ec025c03cb03250466049004a704ba04e1043905d905bf06d607fb08;
    inBuf[4066] = 256'hf209930adf0ad00a720aee095009a008e40710072a06500591040304b6038d03;
    inBuf[4067] = 256'h68033703e3026e02eb016401e0006500eeff78ff08ffa6fe62fe3dfe37fe5bfe;
    inBuf[4068] = 256'h9dfee7fe3cff92ffdcff1a00410055006c008c00bd0005014d0182019a017b01;
    inBuf[4069] = 256'h2801b000090045ff6dfe70fd66fc71fb92faf1f9aaf999f9b0f9d4f9c0f96bf9;
    inBuf[4070] = 256'he6f827f855f795f6cdf5faf424f427f323f250f1a4f030f00bf003f00ef035f0;
    inBuf[4071] = 256'h4bf051f056f02df0d6ef68efd3ee3deec7ed54edfdecd8ecb8ecb3ecdfec0eed;
    inBuf[4072] = 256'h4bed8eed88ed41edd6ec34ec9feb4feb21eb2eeb77ebb2ebe5eb1aec1fec18ec;
    inBuf[4073] = 256'h22ec14ec0bec1fec2cec57eca8ece5ec1ded4eed41ed12edcfec5aecddeb71eb;
    inBuf[4074] = 256'h04ebc9ead6ea10eb98eb5fec2bed0eeef1ee92ef00f035f009f0b3ef58effbee;
    inBuf[4075] = 256'hdeee0fef68ef05f0e3f0e0f11cf386f4daf510f7fff777f8a5f8a2f86af832f8;
    inBuf[4076] = 256'hf6f793f733f7def686f666f687f6c4f631f7b2f70ef855f874f83df8d6f74bf7;
    inBuf[4077] = 256'h9bf612f6d1f5d1f531f6d5f67cf72bf8dbf871f902fa7efab3faa8fa63faf6f9;
    inBuf[4078] = 256'hb0f9c1f934fa0cfb17fc0cfdc8fd25fe0bfe97fde2fc0bfc56fbe4fac0faf1fa;
    inBuf[4079] = 256'h58fbc0fb13fc3efc43fc42fc49fc49fc38fcfafb85fbe8fa40fab8f96ff96cf9;
    inBuf[4080] = 256'ha9f918fa9afa24fba6fb09fc54fc85fc92fc91fc83fc4dfc06fcb7fb5bfb2afb;
    inBuf[4081] = 256'h4dfbc7fbb8fc09fe66ffbd00ee01c1025503bd03e5030004200435047604ed04;
    inBuf[4082] = 256'h7e05560665078208da095f0bde0c6b0ede0f03110a12e9128f134c141615c915;
    inBuf[4083] = 256'h9d167a172e18e5187419ac19cb19c7199f19b419fb19501ae31a7a1bdd1b471c;
    inBuf[4084] = 256'h9e1cce1c221d781db71d281eb11e411f232034215922c8233d258926cc27b728;
    inBuf[4085] = 256'h22294e291b299328172891270f27e226de26f6265d27cc27242885289f286028;
    inBuf[4086] = 256'h012856277a26b825df2404246223bc221d22b1211b215620861f651e1a1df71b;
    inBuf[4087] = 256'hd61ae3195719e8189e18951875183b18f4173c171416a214c012b110ca0ef50c;
    inBuf[4088] = 256'h650b500a850918091c0947099009ec090c0af009a60900091508fb069a052304;
    inBuf[4089] = 256'hc30271015e00a3ff16ffc4feb5feb3fec2fee1fedafeb4fe80fe29fecefd90fd;
    inBuf[4090] = 256'h56fd28fd12fdeffcc5fc9ffc62fc10fcb2fb29fb80fad7f931f9a9f85bf83ff8;
    inBuf[4091] = 256'h56f8a9f826f9bef966fa09fb95fb0afc6dfcc6fc23fd8efd04fe83fe05ff83ff;
    inBuf[4092] = 256'hf9ff6100b200e900110134015f01a30101026b02e1025603bd031b0464047804;
    inBuf[4093] = 256'h4804c903eb02cd019d0073ff65fe7dfdadfcf7fb77fb3ffb62fbe7fbb7fcbdfd;
    inBuf[4094] = 256'hf2fe3a008201c202c7035e046f04df03b30227016dffb5fd35fcf6fa01fa6ef9;
    inBuf[4095] = 256'h31f935f972f9cef938faadfa17fb7afbe4fb33fc5ffc6dfc3afcc9fb36fb6efa;
    inBuf[4096] = 256'h85f99bf89cf7a9f6f6f57ff563f5bff567f653f76ff86bf937fad0fafbfacffa;
    inBuf[4097] = 256'h67fa9bf992f877f720f6b3f458f3eef1a8f0bcef00ef8fee7fee86eeb1ee12ef;
    inBuf[4098] = 256'h60efa8efefefd9ef6befb7ee7fedfdeb79eacfe834e7d8e57be438e33be250e1;
    inBuf[4099] = 256'h91e00fe082df09dfc8de91de91ded7de12df4edf81df61df1cdfc9de37dea1dd;
    inBuf[4100] = 256'h1edd81dc16dc03dc1edc98dc5fdd14dec8de63dfa8dfebdf40e07fe0f3e093e1;
    inBuf[4101] = 256'h1be2cee29ce33ae4d6e44fe554e51be5b2e40be494e365e355e39ae312e470e4;
    inBuf[4102] = 256'hd9e438e563e5a5e5f9e53be6a8e62ce786e7d9e703e8d2e784e72ce7c3e695e6;
    inBuf[4103] = 256'hb2e619e701e858e9f8eaf6ec18ef12f1e3f25af460f529f6aff6f4f63ff78cf7;
    inBuf[4104] = 256'hddf767f817f9cbf987fa15fb60fba1fbe3fb42fcfbfcf2fd07ff380047011002;
    inBuf[4105] = 256'ha802f102e402b602710224020502100234027002aa02d202f90220035303a303;
    inBuf[4106] = 256'h08047f0404058505f5054e067e06810660062a06f105c305ac05b005c505e805;
    inBuf[4107] = 256'h21066906bb061007430745072407ed06c106c206f1064607b5071b0860087d08;
    inBuf[4108] = 256'h5f08fc075e078f06b005ee045304e3039a034603ce024902bf0143010401fd00;
    inBuf[4109] = 256'h0e01360162018e01de015402e5029b035504f3048605fc054406790681064f06;
    inBuf[4110] = 256'h1406e405cc050b069d065f0757085c094b0a3e0b200cd00c660dc90de40dd50d;
    inBuf[4111] = 256'h920d230dcd0c970c810cbb0c2b0db20d680e180f960f03104810591072108810;
    inBuf[4112] = 256'h9210c610041130117b11c8110e12881209137913041469148514a014a0148114;
    inBuf[4113] = 256'ha81404157b1541161617cc179d185a19ec19a01a421bb71b431cb51cfa1c661d;
    inBuf[4114] = 256'hd91d481efe1ec01f66202621c7213122a522f7221a234a2358233e2341234723;
    inBuf[4115] = 256'h5823ad230c246324cb24fe24f324cf2457249923d622f4211a2193203a200d20;
    inBuf[4116] = 256'h1a20172002200220ec1fda1fe21fa01fff1e131ea91cf11a3f198517ed15a314;
    inBuf[4117] = 256'h75137712db1175114911591152112b11f3107510bf0feb0eca0d6b0cf60a6009;
    inBuf[4118] = 256'he707c506e60555050e05c9047a041404650385029d01bc001700c1ff9effabff;
    inBuf[4119] = 256'hc7ffb7ff80ff18ff72feb3fdd7fcd0fbbffab2f9bcf80ff8b6f7b2f712f8b4f8;
    inBuf[4120] = 256'h73f937fabbfad0fa6bfa74f90af883f60df5d7f306f379f212f2c3f162f1f8f0;
    inBuf[4121] = 256'ha3f05bf02ef027f023f029f049f063f07af097f09bf094f093f080f069f051f0;
    inBuf[4122] = 256'h09f0a0ef37efcfee9eeec0ee0aef74efefef43f082f0bbf0d0f0dbf0e1f0bbf0;
    inBuf[4123] = 256'h92f081f06ef080f0bdf0eef01ef14cf155f157f14ef114f1d2f094f03cf002f0;
    inBuf[4124] = 256'hecefcfefd4ef00f027f069f0b7f0cbf0b4f063f0b8ef03ef77ee0fee06ee56ee;
    inBuf[4125] = 256'hbaee45efe0ef4cf0b9f03cf1b3f14ff219f3d8f3a2f45ff5bcf5c3f577f5b7f4;
    inBuf[4126] = 256'hcbf3f1f22bf2c4f1d9f130f2caf28bf31cf47cf49cf442f492f3a1f256f101f0;
    inBuf[4127] = 256'he6ee00ee8eeda3edf2ed6feee7eefbeeb7ee1eee0dedd1eba6ea88e9cce894e8;
    inBuf[4128] = 256'hb1e838e902eaa0ea1aeb6deb6beb5deb70eb8bebdaeb52eca7ecfbec5aed9bed;
    inBuf[4129] = 256'hf7ed78eee2ee5eefeeef4cf09ef0edf001f102f1edf088f0ffef60ef83eeabed;
    inBuf[4130] = 256'h04ed70ec26ec34ec5eecb7ec27ed64ed80ed76ed12ed83ece1eb19eb74ea12ea;
    inBuf[4131] = 256'hd9e9fae970ea01ebbaeb80ec1bed9fedfced19ee36ee65ee9eee13efb3ef46f0;
    inBuf[4132] = 256'hddf05df1aff10cf27ff202f3c4f3baf4c0f5e0f6f9f7ebf8c4f972faeafa53fb;
    inBuf[4133] = 256'hadfbf5fb4bfca1fcecfc3dfd85fdc0fd01fe3efe75febbfe0bff70fffbff9a00;
    inBuf[4134] = 256'h4401ed017a02e3022603390334032a032403420394030f04ae045f05fe057906;
    inBuf[4135] = 256'hbb06c706cb06df061a07a20776088509c60a060c100dcc0d110ed90d5e0dce0c;
    inBuf[4136] = 256'h580c3d0c850c250d110e0c0fe30f8b10dd10ca106d10c40fd90ed50db70c920b;
    inBuf[4137] = 256'h9f0ae2096109390948096b099e09b909b509b409aa099f09b409cd09e109010a;
    inBuf[4138] = 256'h0c0afe09f709e509d109eb092d0a960a340bd40b5b0cda0c3a0d7e0dc70dfc0d;
    inBuf[4139] = 256'h0b0ef80d9d0dfd0c470c750ba10afc09750917091b096b09fc09df0acf0b9f0c;
    inBuf[4140] = 256'h5b0dd10df20df00db40d490df30c9e0c4e0c450c560c640c990cc40cda0c240d;
    inBuf[4141] = 256'h830dec0da50e7b0f481041112c12db128113e813f9130414f013c213d3130214;
    inBuf[4142] = 256'h4314e314b1159116c4170919331a6d1b711c191da41de31dc91dac1d751d2d1d;
    inBuf[4143] = 256'h2f1d5c1d9f1d2b1ebe1e3d1fe21f7a20fb20a0212522682297227022e6214821;
    inBuf[4144] = 256'h7f20a11f011f771efa1db71d711d261d101dfe1cfa1c3c1d811dc41d211e4c1e;
    inBuf[4145] = 256'h461e4a1e2e1e051e011ee91dc01da31d481db51c0d1c221b141a1a1915182b17;
    inBuf[4146] = 256'h7516ae15d914fe13e812bf11ad108f0f890eac0dc20cdf0b100b2d0a5c09a908;
    inBuf[4147] = 256'hf50769071607db06d106de06bc066e06e005f604e403bd02850174008dffc3fe;
    inBuf[4148] = 256'h38fedffda1fd86fd5efd04fd82fcb0fb87fa30f998f7c9f505f453f2d2f0c5ef;
    inBuf[4149] = 256'h1cefcaeedfee22ef7cef01f081f0f0f067f1b3f1c1f1a6f136f173f083ef5aee;
    inBuf[4150] = 256'h20ed19ec41ebbaeaa2eac3ea0beb72ebb7ebceebb5eb3eeb80ea95e972e85ee7;
    inBuf[4151] = 256'h8ce6eae5a1e5bae501e68be651e714e8dfe89ee906ea2bea12eaa5e931e9dde8;
    inBuf[4152] = 256'ha3e8c1e840e9eee9e1eaf5ebd6ec91ed12ee2fee2aee21eefeedf3ed02eefded;
    inBuf[4153] = 256'h09ee25ee33ee65eebeee0fef70efcdeff3ef01f0f9efc3ef96ef7eef6bef94ef;
    inBuf[4154] = 256'hfbef81f048f13ef227f312f4e4f46ef5cbf5eaf5adf543f5b8f40ff49af369f3;
    inBuf[4155] = 256'h68f3c2f356f4e5f489f52bf699f6f9f63cf737f720f7f9f6abf673f656f636f6;
    inBuf[4156] = 256'h43f679f6b9f630f7d8f782f846f90cfa99fafafa17fbc0fa15fa1ff9daf78df6;
    inBuf[4157] = 256'h63f561f4b4f35bf32bf32ef34cf35cf370f382f378f36ef35cf31ff3caf254f2;
    inBuf[4158] = 256'hadf100f163f0d9ef94ef9cefd6ef53f001f1b1f168f212f38bf3e2f315f419f4;
    inBuf[4159] = 256'h11f407f4f4f3fcf31df43cf472f4b7f4f1f42df561f574f573f54ff5f7f48af4;
    inBuf[4160] = 256'h11f48af310f39bf211f280f1e8f04bf0d8efa6efb3ef03f073f0ddf036f16df1;
    inBuf[4161] = 256'h74f168f15ef166f1a0f11bf2cbf29ff379f432f5bef522f66cf6bcf624f7a0f7;
    inBuf[4162] = 256'h29f8aff820f980f9ddf944fac3fa5dfb03fca1fc27fd81fda4fd96fd63fd17fd;
    inBuf[4163] = 256'hcdfc97fc7dfc8efcd6fc51fdfafdcbfeacff87004b01d7011102f4017701a800;
    inBuf[4164] = 256'hbaffdbfe39fe00fe2ffeadfe64ff2800d3006501d701270267029402a802b002;
    inBuf[4165] = 256'haf02a902b502df022b03a3033c04e904ab056c062607de0782080f0994090a0a;
    inBuf[4166] = 256'h780af40a6d0bd30b1e0c2f0c040cbb0b5f0b020bc30a8f0a5d0a450a3e0a480a;
    inBuf[4167] = 256'h780aad0ac40ab90a700aed096909f208900870088308b9082b09c309610a130b;
    inBuf[4168] = 256'hb60b300ca10c000d470d980dd70de40ddf0db80d7a0d720db00d350e1f0f3a10;
    inBuf[4169] = 256'h53117212671310148e14c614a7145b14d51320137c12df115511181110113511;
    inBuf[4170] = 256'hb0114d12e6128713f2130d140514bd133a13bb12221276110211bb10ab101411;
    inBuf[4171] = 256'hc711a112ae1390140f153f15ed1428145a139b121d123a12ce12ac13d314e915;
    inBuf[4172] = 256'hbb165f17a5178e175717ef1675164016451693164b172e181c19251afe1a901b;
    inBuf[4173] = 256'hea1bd41b4d1b8f1a8e1973188217a216df155015c4144114e4137d131113b212;
    inBuf[4174] = 256'h2e129211fb104a10940ff50e490e9a0df40c340c6d0bb40af0094009c5087608;
    inBuf[4175] = 256'h7308c4084009e109840ae00ae80a8c0ab3097e080c076c05da0383027b01e600;
    inBuf[4176] = 256'hbe00d900230166016d013001910088ff39feaffc03fb6ef9fff7c9f6ecf55af5;
    inBuf[4177] = 256'h11f51df55bf5baf530f67bf67bf629f663f53ef4f4f292f14df05befabee4eee;
    inBuf[4178] = 256'h4dee6cee97eec6eec4ee98ee56eee1ed53edc5ec20ec8beb2eebf1eaf9ea55eb;
    inBuf[4179] = 256'hcdeb66ec20edc1ed4ceebceedaeeb7ee66eecfed26ed92ec05eca2eb76eb62eb;
    inBuf[4180] = 256'h7bebbfebf9eb30ec58ec47ec18ecdbeb7eeb33eb12eb0beb42ebb6eb3aecd6ec;
    inBuf[4181] = 256'h74edebed54eeb2eef1ee3aef8befc8ef14f075f0d9f064f10af29ef230f3b2f3;
    inBuf[4182] = 256'hfef33df47bf4acf401f57cf502f6abf664f7fcf783f8e9f819f946f981f9bdf9;
    inBuf[4183] = 256'h27fab2fa30fbb1fb26fc70fcb5fcf3fc0ffd28fd30fd07fdcffc8ffc43fc1efc;
    inBuf[4184] = 256'h27fc4bfca3fc17fd76fdcffd0dfe10fef4fdbafd5afdfefcaafc4efc04fcc9fb;
    inBuf[4185] = 256'h90fb82fbb2fb1efcdafcc8fdb7fe9aff4d00ac00cf00be007b003100edffa4ff;
    inBuf[4186] = 256'h66ff27ffd5fe8dfe57fe37fe49fe84fecbfe17ff51ff5dff46ff07ff98fe10fe;
    inBuf[4187] = 256'h7afde4fc77fc3cfc2bfc42fc64fc78fc7efc75fc5dfc40fc1afce5fbb1fb84fb;
    inBuf[4188] = 256'h63fb5efb6efb85fba0fbb4fbc0fbcefbe2fbfdfb25fc5cfc9efcf0fc56fdcdfd;
    inBuf[4189] = 256'h4ffed5fe54ffc1ff15004a005e005c005000440043004e005b00640060004500;
    inBuf[4190] = 256'h1600daff8cff37ffedfeb8feaafecefe1cff89ff06007800d40019013b013d01;
    inBuf[4191] = 256'h2c010f01fd000c014501b20157022103fd03d6048d0519067f06bc06e2060d07;
    inBuf[4192] = 256'h47079d070d087d08d80810090c09d90896085608390855089708ef0844096909;
    inBuf[4193] = 256'h5009fb086308a007da0625069f05630562059305e8053b068106bb06d506ca06;
    inBuf[4194] = 256'ha0064806cb054c05d9048b047f04a104e10439058f05da052306550668066c06;
    inBuf[4195] = 256'h5d06460647065d068406c306020738077607b207e1070408ff07c60773070e07;
    inBuf[4196] = 256'haa066b0648062b061206db057305ea043c047703c6023302d101c101ee013c02;
    inBuf[4197] = 256'ha302f40210030103bc024e02ec01a9019e01f2019102600350042b05ca052f06;
    inBuf[4198] = 256'h4b062206de05890533050a050d053b05a3052406a0061c077907a807c207be07;
    inBuf[4199] = 256'h980770073c07f806c50699066f065b0647061c06ea059c052b05c20468042604;
    inBuf[4200] = 256'h29046704d0046c0512069806fe0624070007bb0660060a06ec0506065306e906;
    inBuf[4201] = 256'ha70772084709fe09790ac80adf0ac30aa40a8e0a920ad70a510bf30bc30c980d;
    inBuf[4202] = 256'h4d0edd0e210f0f0fc10e390e880ddc0c390cac0b510b170bf60afe0a150b340b;
    inBuf[4203] = 256'h630b800b770b3e0bb20ad309c908ac07ac060006a905ae050b0693062707b807;
    inBuf[4204] = 256'h1c0842083208e4076907e4065a06de05850544052105260542057605c1050e06;
    inBuf[4205] = 256'h5a06a106ce06dd06cc068c062806a70508055b04a303df021b0257019500e2ff;
    inBuf[4206] = 256'h3aff90fee9fd36fd74fcb6fb00fb62faf6f9baf9a6f9b7f9ccf9cbf9b0f966f9;
    inBuf[4207] = 256'hf3f86ff8e4f767f719f7f1f6ebf608f723f72af71ef7eef6a1f650f6faf5b4f5;
    inBuf[4208] = 256'h96f595f5b7f501f650f694f6c1f6b4f66df6fdf55ef5b0f417f497f351f359f3;
    inBuf[4209] = 256'h98f309f49af418f571f59cf579f51bf593f4d9f30ef352f2a9f136f110f11cf1;
    inBuf[4210] = 256'h5ff1cbf132f294f2f2f22ef35cf386f394f39bf3a4f39af398f3adf3c6f3f9f3;
    inBuf[4211] = 256'h47f48ef4d8f41ff545f562f57ef58af59ef5c3f5dff500f624f62af61ff603f6;
    inBuf[4212] = 256'hc6f586f557f52df51ff52cf533f53ff54cf542f536f52bf505f5d7f4a4f45cf4;
    inBuf[4213] = 256'h1df4f9f3e4f3f5f329f460f49ff4daf4f0f4f3f4e5f4b7f489f466f443f43bf4;
    inBuf[4214] = 256'h4ff462f47ff49bf497f486f46df443f42ef438f455f498f4f3f445f593f5ccf5;
    inBuf[4215] = 256'hd4f5bef589f52cf5cff480f43ff432f459f4a2f418f5a9f532f6b7f622f757f7;
    inBuf[4216] = 256'h62f741f7f2f69ef659f62cf637f678f6d5f654f7def759f8d1f83cf988f9c1f9;
    inBuf[4217] = 256'hdef9cff9acf97bf93df90cf9e3f8b6f891f86ef847f835f836f845f870f8acf8;
    inBuf[4218] = 256'heef845f9a6f907fa6ffaccfa11fb4dfb7afb9bfbc7fbfdfb40fca6fc2afdcdfd;
    inBuf[4219] = 256'h9dfe86ff780069013802ce022a033f031a03d80287023c020d02f201ea01fa01;
    inBuf[4220] = 256'h15023f027f02c30204033b0352034d033b0320030f03100310030703e802a002;
    inBuf[4221] = 256'h3e02db0187016a0196010602bb02a00391047f055206ec065407870788077707;
    inBuf[4222] = 256'h63074e074c0750074a0749074a0752078107d8074c08e3088209100a910af40a;
    inBuf[4223] = 256'h320b5d0b6c0b5d0b440b1a0bdd0aa50a680a260af709d309bb09c109d209df09;
    inBuf[4224] = 256'hed09e109b909940970095a09690985099d09b509b709a709a1099d09a209c109;
    inBuf[4225] = 256'he709170a670ac80a390bbf0b330c840cb20ca10c550ce80b520bac0a1b0aa409;
    inBuf[4226] = 256'h5a094e095f097809890969091709a8081c088d071507a5064006e5057905fd04;
    inBuf[4227] = 256'h7c04eb035c03de026502f40193012f01d500950064004f005d007900a500e600;
    inBuf[4228] = 256'h28016d01b501ec0113022f023a024002520269028e02c602030342038103aa03;
    inBuf[4229] = 256'hb4039e035903e9025b02b20101016100d6ff6eff2fff08fff2fee9fee3fee5fe;
    inBuf[4230] = 256'hf5fe0cff20ff2cff1efff8fecbfea5fe9cfec2fe15ff89ff1100950004015e01;
    inBuf[4231] = 256'h9e01cb01f5011f024b028002b702e702150337034d0364037f03a403df032604;
    inBuf[4232] = 256'h6d04ad04d404e004dc04d004c404c504ce04da04ef040905270552058405bb05;
    inBuf[4233] = 256'hff054a069906f0063f077a079f07a30788075a071907ca067b063006f705e605;
    inBuf[4234] = 256'hfe054006aa0622079a0704084e087108710850081d08ee07c507aa079b078907;
    inBuf[4235] = 256'h7107590744074107570778079a07a9078e074107c40618064f057c04a803e402;
    inBuf[4236] = 256'h33028f01fc0079000400abff6eff49ff3cff3bff38ff32ff1dfff5febcfe6dfe;
    inBuf[4237] = 256'h08fe99fd20fda5fc3bfce9fbbefbccfb13fc8bfc27fdc8fd55fec0fef9fefdfe;
    inBuf[4238] = 256'hd1fe6bfed0fd0dfd2bfc44fb78fad3f967f939f938f957f984f99ef995f960f9;
    inBuf[4239] = 256'hfaf878f8f6f782f734f713f713f730f765f7a2f7e9f73ff897f8f8f862f9c3f9;
    inBuf[4240] = 256'h18fa56fa6afa5bfa31faf6f9c9f9bdf9d2f907fa4afa7dfa93fa85fa4dfa03fa;
    inBuf[4241] = 256'hbbf97ff96df98ef9def95efaf9fa8bfb00fc40fc3efc0efcc5fb76fb3cfb20fb;
    inBuf[4242] = 256'h1ffb42fb8afbf1fb78fc0bfd8cfdf0fd2ffe4efe6dfe9efee7fe4dffc0ff2c00;
    inBuf[4243] = 256'h8e00dc0008011101eb0095002000a6ff3dff03fffefe27ff77ffe1ff5200bf00;
    inBuf[4244] = 256'h170143013d01010199001c00a2ff39fff3fed5fedffe0fff5bffadfff3ff1500;
    inBuf[4245] = 256'h0400bcff48ffb3fe10fe71fde4fc79fc3bfc2afc40fc73fcaffce7fc16fd37fd;
    inBuf[4246] = 256'h4dfd58fd4efd28fdebfc9ffc5cfc40fc5afcb0fc37fdd5fd6ffef3fe4eff7bff;
    inBuf[4247] = 256'h7eff58ff17ffd2fe96fe73fe70fe7cfe88fe8bfe7cfe63fe54fe54fe65fe85fe;
    inBuf[4248] = 256'ha2feb3feb8feadfe8ffe63fe1ffec6fd63fd00fdaefc83fc81fcaafc01fd76fd;
    inBuf[4249] = 256'hfdfd8cfe0dff71ffb2ffc6ffb2ff8aff5bff38ff35ff4fff7bffa7ffb5ff92ff;
    inBuf[4250] = 256'h41ffc8fe3ffec4fd63fd1ffdfbfce7fcdafcd0fcbcfc92fc51fcf1fb7bfb0afb;
    inBuf[4251] = 256'haffa84fa9afaedfa6ffb0efca9fc25fd73fd87fd6dfd40fd1afd16fd46fda2fd;
    inBuf[4252] = 256'h14fe89fee3fe16ff27ff1afffcfed9feb1fe83fe55fe28fe05fe01fe21fe68fe;
    inBuf[4253] = 256'hd0fe42ffa7fff3ff15000e00e9ffaeff6bff32ff0bff03ff25ff6bffcfff4000;
    inBuf[4254] = 256'ha300e000ea00b8005700e7ff80ff42ff3bff61ffa1ffe1ff0200faffc8ff73ff;
    inBuf[4255] = 256'h10ffb9fe7bfe66fe7efeadfedffefbfee9feaffe60fe14fef1fd09fe5dfee3fe;
    inBuf[4256] = 256'h83ff18008a00c100ad005600caff1fff77fee3fd72fd2ffd18fd25fd56fd98fd;
    inBuf[4257] = 256'hdbfd18fe3dfe42fe2efefafdaffd61fd1bfdf7fc0ffd63fde4fd7cfefbfe49ff;
    inBuf[4258] = 256'h60ff41ff04ffc7fe91fe70fe72fe8efec7fe19ff65ff9cffb3ff95ff52ff02ff;
    inBuf[4259] = 256'habfe66fe41fe31fe3dfe5ffe7bfe8cfe86fe55fe0dfec5fd88fd77fd9efde5fd;
    inBuf[4260] = 256'h46fea8fee6fe05ff06ffeafed4fedefe0bff76ff1e00e700cd01b80283033504;
    inBuf[4261] = 256'hca043b05a70515067a06e2063d077607a007c207e00721088308f9088809170a;
    inBuf[4262] = 256'h8a0aeb0a2a0b3d0b3d0b2b0b0a0bfc0a000b120b3e0b6f0b8f0ba30b9b0b6e0b;
    inBuf[4263] = 256'h360bf70ab90a9c0a980aa20ac30adf0aea0af50af70af30aff0a120b2d0b640b;
    inBuf[4264] = 256'haf0b0a0c7b0ce00c260d4c0d440d180de50ca80c620c170caf0b230b850ad509;
    inBuf[4265] = 256'h2a09a2083e080408f607f807f707e807b0074907bf0611064e058c04ca031003;
    inBuf[4266] = 256'h6402be01220197002100cdffacffbbfff5ff4e00a700ec000a01f500ae004300;
    inBuf[4267] = 256'hc1ff41ffddfea8feb0fef4fe64ffe7ff6000b600dd00d500a60061001000bfff;
    inBuf[4268] = 256'h71ff23ffd0fe71fefffd7ffdf4fc68fceafb7efb25fbddfa9afa4ffafbf99cf9;
    inBuf[4269] = 256'h38f9e5f8aef89ff8c2f806f953f991f9a0f974f918f99ff82bf8e2f7d1f7fbf7;
    inBuf[4270] = 256'h5bf8d8f85ef9e3f955faaffaf6fa29fb53fb8afbd3fb30fc9bfcf9fc39fd58fd;
    inBuf[4271] = 256'h55fd45fd45fd59fd88fdcffd22fe82fef7fe7eff1400b00033018b01b0019701;
    inBuf[4272] = 256'h4901d300370084ffd1fe34fed2fdcbfd27fedefed2ffcb009a011c023902fe01;
    inBuf[4273] = 256'h8701fb00870052006a00d4007f0146020803a6030b0439043c0425040704f103;
    inBuf[4274] = 256'he403e503ec03f603fe03ff03f603e303c5039d036c032803d0026202e3016601;
    inBuf[4275] = 256'h0101c200b900e1002f01960105026902b602db02cd0294024102f001c401cd01;
    inBuf[4276] = 256'h09026d02d7022d03640373035d0337030b03e602d802da02dc02d1029d023702;
    inBuf[4277] = 256'hb2012601bb009900c4002c01b30125025b024702e1013a017700acfff2fe67fe;
    inBuf[4278] = 256'h15fe0cfe59feecfeaaff7000000135010a018700d9ff37ffbcfe78fe6ffe90fe;
    inBuf[4279] = 256'hd2fe37ffabff18005f004f00ceffe8febcfd8efcacfb44fb6efb21fc26fd40fe;
    inBuf[4280] = 256'h2fffafff98ffe6fea8fd1efca9faa2f95bf9fbf95bfb2afdfefe650024013801;
    inBuf[4281] = 256'hc40009004fffb4fe48fe0dfee7fdc1fd8dfd34fdbbfc3ffce2fbdafb4ffc3dfd;
    inBuf[4282] = 256'h77feb3ff9100c7003f0007ff62fdb1fb4cfa82f980f93ffa8dfb1ffd90fe88ff;
    inBuf[4283] = 256'hd5ff66ff5cfefffc97fb6ffac0f999f9f3f9b3faa3fb8dfc47fda1fd7dfddafc;
    inBuf[4284] = 256'hbffb4dfac1f851f732f68df564f5a8f542f60af7dcf7a1f836f984f984f935f9;
    inBuf[4285] = 256'hadf821f8bcf7aaf704f8b7f894f966faf5fa26fb08fbbafa69fa3efa40fa65fa;
    inBuf[4286] = 256'ha2fae1fa1afb4cfb64fb4dfbf8fa5bfa87f9b0f807f8b4f7caf733f8cff885f9;
    inBuf[4287] = 256'h3ffaf6faa8fb44fcb3fce6fcd7fc99fc56fc2dfc34fc6afcbafc0ffd6bfdd8fd;
    inBuf[4288] = 256'h6ffe3dff2800fb007301560197005cffeafd92fc91fbfffae2fa35fbf6fb21fd;
    inBuf[4289] = 256'ha3fe3e009a01540227020a013aff26fd48fb0bfab3f960fa10fc9efec1010505;
    inBuf[4290] = 256'hd607a009fc09cf08630652035c0035fe56fde9fdc5ff7a026f05f80776098009;
    inBuf[4291] = 256'hfe073a05d801b2fe93fc01fc10fd5fff440202050007ef07c707b5060c052a03;
    inBuf[4292] = 256'h71014000dcff5c00a1014e03ed04130687064c069a05bb04e50332039c021302;
    inBuf[4293] = 256'h97013c01210164010402da02a3031204eb031d03c101110062fe01fd2afc00fc;
    inBuf[4294] = 256'h81fc82fdbefeddff8f00b0005500c1ff50ff3fff8dfffcff2a00c0ffabfe21fd;
    inBuf[4295] = 256'h8efb6ffa22fac4fa38fc32fe470007020c03ff02bc015fff46fc14f985f632f5;
    inBuf[4296] = 256'h74f536f7faf90afda4ff2c016301640090fe76fcaafa98f984f975fa2cfc46fe;
    inBuf[4297] = 256'h4400a9012b02bf01950015ffacfda3fc20fc1efc78fc0ffdcefd99fe60ff0500;
    inBuf[4298] = 256'h5f005800e9ff19ff12fe00fd0cfc63fb2cfb7bfb60fccefd8eff5201b9026103;
    inBuf[4299] = 256'h1e03ff014f0098fe68fd26fd02fedbff4a02d8040d0788082009cd08a207e305;
    inBuf[4300] = 256'he90321020801fa000d0210048106b4081a0a610a8b09f7072206770441038c02;
    inBuf[4301] = 256'h3602220235026b02e002aa03d004510602089d09d30a440ba70afa087906a903;
    inBuf[4302] = 256'h4001d5ffb6ffd900d402170523079e085a09560990080e07f404810219003ffe;
    inBuf[4303] = 256'h55fd89fdc2fe9f00a3025d047505c1054405150464028000c5fe96fd48fdfbfd;
    inBuf[4304] = 256'h8cff9b01a0031a05b90568054f04bd0202016dff41feb5fdebfde0fe5700d901;
    inBuf[4305] = 256'hd502d702b901c6ff9cfdf4fb54fbe2fb54fd22ffbc00b601e50155013700d0fe;
    inBuf[4306] = 256'h75fd7cfc3bfce8fc7bfea500da027f042505ba048b0326022101d0003101f501;
    inBuf[4307] = 256'ha702e6028b02a0015a00fbfeb1fda9fc0bfcf7fb89fcc4fd79ff5601ef02d103;
    inBuf[4308] = 256'haf0374023c0069fd8efa4af834f7abf7a7f9c1fc46005a035305dd0501052203;
    inBuf[4309] = 256'hd30097fee6fc12fc40fc80fdadff650216051007ac079c060b0496003afdf6fa;
    inBuf[4310] = 256'h72fadffbd7fe7f02de0514088c0831076004d4008dfd81fb5afb47fdd7000f05;
    inBuf[4311] = 256'hc808000b290b61094806c102b7ffcefd47fd1afeecff3a02810445062f072407;
    inBuf[4312] = 256'h36069c04b002c6002eff2afed7fd27feeffee0ffb4004b01b0011202a6027003;
    inBuf[4313] = 256'h4104c804b504ea0397021801d5ff18ffe8fe20ff90ff10009b003b01ee019502;
    inBuf[4314] = 256'hfb02e00230020e01caffc3fe36fe1ffe4bfe7afe8cfea0fef4feb8ffe4002402;
    inBuf[4315] = 256'hfa0209033b02d1004bff1afe79fd65fdaefd20feabfe4bff0700db00ab015902;
    inBuf[4316] = 256'hd2020b03ff02ab020002fe00c9ff9efecafd8cfde5fda4fe7eff28008b00c100;
    inBuf[4317] = 256'hec00290173019d0188013c01da009d00a200c100ae001a00e2fe45fdbffbc3fa;
    inBuf[4318] = 256'h97fa28fb22fc42fd7cfeecffbd01d003980559067d05ee024fffbafb3bf974f8;
    inBuf[4319] = 256'h5df95dfbc6fd19002402f6038d05ac06f9062c064404b80140ff82fde4fc5afd;
    inBuf[4320] = 256'h78fec5ffdf008d01d101b0011c011400a6fe0afdb4fb1ffb93fb0ffd2dff4201;
    inBuf[4321] = 256'hb602280388021c014cff7afdfffb11fbc2fa15fbe8fbeffcdefd70fe7cfe19fe;
    inBuf[4322] = 256'h7afddcfc7bfc7bfce2fcb0fdcafee9ffb700ce00edff2efe09fc2cfa44f9a8f9;
    inBuf[4323] = 256'h31fb61fd93ff44014702b402b6027202e8010701deffadfed2fdb0fd6afebeff;
    inBuf[4324] = 256'h26010602f401f90086ff37fe99fdddfdd0fe0c0031010e02b7025003de033204;
    inBuf[4325] = 256'hfb03ee021a01f5fe3afdb4fcdbfd9b0058041a08d90ae10b000b8c084a051f02;
    inBuf[4326] = 256'hc3ff9ffeb4feb5ff4001fb029a04e805ad06a1069a059b03f20038fe1dfc1ffb;
    inBuf[4327] = 256'h60fb97fc29fe7dff2e0021007fff89fe69fd3bfc14fb17fa84f99ff97bfae9fb;
    inBuf[4328] = 256'h7bfdacfe24ffe2fe29fe61fdd9fc97fc78fc57fc2afc19fc5dfc05fde6fdaffe;
    inBuf[4329] = 256'h13ff07ffd2fed2fe4dff2f0009015001b30045ff85fd21fc8ffbe5fbd7fcddfd;
    inBuf[4330] = 256'h8dfec5fea5fe73fe70feabfe11ff89fff7ff52009500ab007200d8ffddfeabfd;
    inBuf[4331] = 256'h85fca1fb1dfb05fb5efb3cfcbffdd9ff2b020c04ae049603fb00c4fd3efb7dfa;
    inBuf[4332] = 256'hc7fb6dfe2d01c502a3021a0110ff6dfda1fc74fc60fc0efc9ffba3fbb6fcf9fe;
    inBuf[4333] = 256'he5017f04c905440528032e0031fddefa80f924f9cff974fbeffdd6006a03d304;
    inBuf[4334] = 256'h88049302aefffffc8bfbcefb99fd2f00ac026404ff0479040b030101c6fee7fc;
    inBuf[4335] = 256'hf4fb5bfc30fe0401060455065307e90690050104e7029e021103e403a8040f05;
    inBuf[4336] = 256'hfd049304fe036c03ff02c502be02e7022e036f038203340366022401a5ff44fe;
    inBuf[4337] = 256'h66fd55fd1dfe8eff38018d020f037102b7004bfedefb3ffa1dfabcfbd3fe9702;
    inBuf[4338] = 256'hf005d307aa0785051f02a5fe45fcc0fb20fdb8ff660219043504ce028a0035fe;
    inBuf[4339] = 256'h5ffc29fb5dfabff964f9b3f91efbc0fd15010c048505de044d02d6feccfb3afa;
    inBuf[4340] = 256'h7efa37fc90feb7002a02c702bf026202f101a601a501f601870219035203e502;
    inBuf[4341] = 256'hbc01050033fec1fcf7fbd2fb01fc14fcbffbfbfa05fa4df938f9fcf994fbbbfd;
    inBuf[4342] = 256'h0100e701ff02f802d101d2ff81fd80fb57fa3cfa15fb8cfc33febafffc00e701;
    inBuf[4343] = 256'h7a02a80259028001220053fe41fc2afa59f831f715f738f88bfa9cfdb3001a03;
    inBuf[4344] = 256'h58044e043503640122ffb2fc5cfa88f8c0f770f89ffae0fd65014f0414069806;
    inBuf[4345] = 256'h1506e20440034b0131ff45fdf5fb97fb22fc17fdc6fdaffddafcebfbc4fbfafc;
    inBuf[4346] = 256'h6eff470249047f04b10270ffdcfb14f9c5f70ef89cf9e8fb7cfefa0006034904;
    inBuf[4347] = 256'h77047203760108ffc2fc18fb2cfacff9c4f9f0f961fa3efb8afcf8fd09ff45ff;
    inBuf[4348] = 256'h71febcfca5fab9f869f7eaf635f725f87ff9ebfa0afc8efc5dfcbdfb3cfb6afb;
    inBuf[4349] = 256'h8efc70fe5a007a014701c0ff71fd30fbb2f95df931fadefbfafd1400c101ab02;
    inBuf[4350] = 256'ha502ba014000c1feb9fd6cfdc8fd68fedefee5fe68fe8bfd76fc3ffbfcf9dff8;
    inBuf[4351] = 256'h3bf87df8e3f93dfce6fe0501ea0179013900f3fe46fe47fe74fe24fe03fd4efb;
    inBuf[4352] = 256'hcaf942f909fad2fbe1fd74ff3d0070007f00c6004101900148013d0094febafc;
    inBuf[4353] = 256'h28fb2afae4f963faa7fba8fd3a00f4023f058d0680062205dc024100edfd5efc;
    inBuf[4354] = 256'hd9fb7efc44fee500eb03b806a7084d09aa081c074a05da03250323038303cf03;
    inBuf[4355] = 256'hc0035d03eb02c9023f0343048d05bb067907b1079507730795071408c2084509;
    inBuf[4356] = 256'h40097608f206140568038502de0285042c07390ae10c740e900e2c0da60aa507;
    inBuf[4357] = 256'hd904d402e401ef0195025e03e003fe03ef03030479044c051d066d06f305bc04;
    inBuf[4358] = 256'h3a0310029f01e3017d02ed02fb02e80237035c045b0698081f0a2e0a8f08d305;
    inBuf[4359] = 256'h0b033101b8007101b002d803be049a05d40696087b0abe0ba00bc8098d06d602;
    inBuf[4360] = 256'ha1ffa4fd1ffdcffd3afff900bd026004d405fd06be070308af07a906f704bd02;
    inBuf[4361] = 256'h620093fefdfd0bffa201f504d4072c096408b5051002a9fe94fc72fc3efe7701;
    inBuf[4362] = 256'h4f05cf08130b8b0b0c0afa063403b8ff4ffd50fc74fc23fddefd70fe17ff5100;
    inBuf[4363] = 256'h6b024a055e08c30aa90bb90a17086c04af00befd37fc5bfcf9fd91007f031206;
    inBuf[4364] = 256'hbc073c088707d4059003320138ff14fe01fef4fe9a004d0263038203c202c601;
    inBuf[4365] = 256'h7301630288041507c40883081806390251fed5fb84fb2ffd0000f8028b05c907;
    inBuf[4366] = 256'h010a460c240e9d0ec10c59081f02a8fbc3f6b1f4bcf547f91dfe000308079a09;
    inBuf[4367] = 256'h630a500984068c0265fe31fbddf9c4fa73fdef00270450062307c5068005a003;
    inBuf[4368] = 256'h790176ff23fe0ffe70ffec01b704d806ab073607fa059a04760377024f01e8ff;
    inBuf[4369] = 256'h92fef1fd8ffe5c009a023e047b044c037c0124000d00450118038804e9042704;
    inBuf[4370] = 256'hbe026501a500a40042013c0253035c041b0545059704f2028a00e9fdc1fbaffa;
    inBuf[4371] = 256'h0ffbd9fcabffed02e305d7073e08db06d603ccffa3fb52f89bf6d5f6ddf835fc;
    inBuf[4372] = 256'h1f00cc038406c4074d074a05450206ff5dfcd8fa96fa49fb64fc57fdd9fdf8fd;
    inBuf[4373] = 256'hf5fd1efe95fe33ffa5ff97ffe6fec3fda7fc17fc6cfca4fd58ffee00df01ef01;
    inBuf[4374] = 256'h450149005cffb4fe4bfeeefd80fd19fdfbfc70fd96fe3900e201ff021c031602;
    inBuf[4375] = 256'h39001efe83fc08fce3fcc6fef8008f02d902ad0170ffe6fcd9fac5f9bdf98ffa;
    inBuf[4376] = 256'heefb95fd45ffa5004801e4008affcffda9fce5fca1fe260128037903be01a7fe;
    inBuf[4377] = 256'h8cfbbef9caf93dfb11fd43fe62febafdf8fcb1fc1ffd0dfe08ffb0ffceff4eff;
    inBuf[4378] = 256'h51fe1efd21fce1fbaffc58fe26000e0137009ffd36fa6bf794f61cf84bfbcafe;
    inBuf[4379] = 256'h48011a0280013b00fefe30fed4fdbffdf1fd73fe10ff60ffc6fed5fcdef9e8f6;
    inBuf[4380] = 256'h41f5f5f524f9e8fde702d806eb0803094f07fd0367ff22fa1ef5baf121f1aaf3;
    inBuf[4381] = 256'hb0f8a1fe91032206d4050903e3feb3fa95f76ef68ef77ffa3efe5c017a022601;
    inBuf[4382] = 256'h03fe79fa2df803f8a4f9fafbb6fd11fe4ffd3efc8afb7cfbbbfbb5fb55fb07fb;
    inBuf[4383] = 256'h62fbe2fc4bffa201d9023602aeff20fcbff88cf635f6a4f719faaafc69feaffe;
    inBuf[4384] = 256'h94fdb7fbe7f9f5f818f9d7f993fabbfa2bfa69f909f93af9cef92dfacdf9d8f8;
    inBuf[4385] = 256'hf2f7cdf7ddf8c6fa85fc38fd6cfc5ffafff730f65df59df59af6d8f71af91efa;
    inBuf[4386] = 256'h80fa05fa93f864f644f408f324f388f471f6cff710f830f7aef568f4edf34bf4;
    inBuf[4387] = 256'h60f5daf65bf8b3f98afa61faf9f867f639f383f02aef6fef08f122f3eff44bf6;
    inBuf[4388] = 256'h83f7e9f888fabbfb7efb4af96df519f114eea2ede5ef01f464f88cfbdcfc84fc;
    inBuf[4389] = 256'h2cfbb6f9a7f808f8b9f770f7e0f6fff5dbf4a0f3c6f2b8f29ff374f5c2f7d7f9;
    inBuf[4390] = 256'h4cfb07fc32fc36fc3efc0efc53fbcaf97bf7fbf4f8f2e2f1e4f1b2f2c6f3e3f4;
    inBuf[4391] = 256'h00f627f777f8d2f9d1fa2efbcefadbf9e1f869f8baf8e5f98efb0dfdd4fd7bfd;
    inBuf[4392] = 256'he0fb72f9e7f6fcf45bf426f5d6f699f87ff9e8f8fef68bf4acf284f291f46cf8;
    inBuf[4393] = 256'h22fd66010e04a5045703b2007dfd51fa86f77af585f4e3f4baf6a2f9a5fcbefe;
    inBuf[4394] = 256'h34ff06fe2afceefa3efb3efd0e003e02b9022b011afea0fab3f7c3f5ecf416f5;
    inBuf[4395] = 256'h3ff6a6f852fcb200b7040d07c206ef03afffa5fb4cf91ff96ffafefb97fcbdfb;
    inBuf[4396] = 256'h11fac6f8f4f811fb8ffe1e026c049e04ae0273ff10fc7bf93df832f8d1f899f9;
    inBuf[4397] = 256'h36faaafa52fb7efc38fe3400c90141023a01cffea9fbc9f800f7b9f6e6f707fa;
    inBuf[4398] = 256'h81fce2fed6001a027602b901f5ffaffdb4fbdcfa89fb57fd4cff5d00f3ff57fe;
    inBuf[4399] = 256'h7afc4efb42fb05fcc7fceafc73fc08fc89fc5efe1601b3033905420556047c03;
    inBuf[4400] = 256'h7f037904af050006bb040102befe3ffc68fb4ffc66fec0009b02c00351048304;
    inBuf[4401] = 256'h87045b04f20373031303f2020d030b0384027101200030ff51ffb300f4026d05;
    inBuf[4402] = 256'h69078208d4088e08c60776067a04fd01b6ff88fe2affc801920523093e0b280b;
    inBuf[4403] = 256'h0e09fc05230371015d019e0291049b061c08c208a708ff07260795066e069106;
    inBuf[4404] = 256'hcc06b6061806240522046f036503f903fc045106b8070d09490a1d0b330b740a;
    inBuf[4405] = 256'he208e4064505a0044a052f078d097b0b5a0ccf0b200a2708a5062506da064808;
    inBuf[4406] = 256'hb909af0ac50a0d0a0909180880077707d6078908b009380b120d2a0f0c115212;
    inBuf[4407] = 256'he712a7129911d30f1b0d5209d504540010fd72fc04ff4604ca0a6d109213ec13;
    inBuf[4408] = 256'h3c120f10ea0e280f2510d6103810380ecd0b0d0abe09e90a7d0c420da00ca00a;
    inBuf[4409] = 256'h3708cf0633076e09df0c3e108412691317134112c011c2110b1233129d112810;
    inBuf[4410] = 256'h630ee90c590c000d4c0e5b0f7f0f4e0e350c5b0abc09fc0a1b0e0f1289158b17;
    inBuf[4411] = 256'h6d175e154e121b0f970c550b380bf60b4b0db30ed70fa410e610b9108c109e10;
    inBuf[4412] = 256'h271140126113f413b413931221114d107b107e1197127c127310f00c34091c07;
    inBuf[4413] = 256'h4108c20c64131e1a911e631fbc1cb2170912760db20ab609090ac40a530bb00b;
    inBuf[4414] = 256'he30b3f0c280d800e09108c11a21238139913df132e148e148814bb131b12a80f;
    inBuf[4415] = 256'hd90c730af308c4081c0a8c0c630fcc11ae127211660e780a480773067c08bd0c;
    inBuf[4416] = 256'ha3111c15ef1547143011270e3c0c490b8c0a5d098f07e5058705e5068909420c;
    inBuf[4417] = 256'h890db80c6a0ade077f0612071a097e0b290d480dd50b58095c0682037d01cc00;
    inBuf[4418] = 256'he401d904d908990ccb0e870e130cbe08fe05dd047105b9068a073807c005dc03;
    inBuf[4419] = 256'h7502e8012e0204030d043d05a206f507c5089e0839070405eb02be01d801d202;
    inBuf[4420] = 256'ha80384033c025300dcfecdfe59000f030e0657085409e008120756044e01b1fe;
    inBuf[4421] = 256'h4cfda7fd93ff39025204a904ee02e7ff0cfdf0fb5dfdd900fe0425081c09c107;
    inBuf[4422] = 256'hdb049001eafe67fde6fc0bfd71fdd6fd3bfebbfe68ff58008401bf02bf031d04;
    inBuf[4423] = 256'h7a03c9015cffe3fc3cfbf1faf4fba8fd19ff77ff8bfebbfcd6fab0f9a8f99ffa;
    inBuf[4424] = 256'h21fca4fdd6feb6ff5d00de0035013301b700dcffd2fed9fd1dfd85fce5fb21fb;
    inBuf[4425] = 256'h43faa2f9aaf97efaf3fb89fd7cfe3afea3fcfdf9f2f64ff4aaf268f2a5f30ef6;
    inBuf[4426] = 256'h1ef91afc16fe6cfef5fc15fad5f677f4c4f3e9f44af7abf9f8faa4fac5f828f6;
    inBuf[4427] = 256'hd1f376f288f200f44cf6ccf8d5fab1fb0efb0df921f636f338f193f047f1c2f2;
    inBuf[4428] = 256'h03f46bf4ddf3a5f297f170f151f2fbf3c4f5c1f687f621f5e1f27df09aee76ed;
    inBuf[4429] = 256'h48ed18eeb3ef22f243f57af824fb7bfcbcfbecf8bdf436f0adec02eb32ebcfec;
    inBuf[4430] = 256'h06efe6f023f2c5f2cef281f2eef1e4f09bef78eeceed1fee88ef82f180f3dbf4;
    inBuf[4431] = 256'hfaf4f9f336f206f019eef6ecc7ecd7ed17f0dbf26ef5e4f65cf6dcf30bf0dceb;
    inBuf[4432] = 256'ha1e819e71ee74fe805ea9beb2cedf9eef6f016f3daf476f5aef49af287ef40ec;
    inBuf[4433] = 256'h5de913e7cee5c7e5e6e641e971ec7fefb9f193f2dcf15cf00fef97ee66ef21f1;
    inBuf[4434] = 256'hc1f289f3dbf272f0eeec23e9d3e508e44de46ee6f4e9d0ed9bf098f191f0f2ed;
    inBuf[4435] = 256'h0aebffe84ee81de9cfea63ec75edf5ed05ee45ee00ef0bf059f1a4f28df31bf4;
    inBuf[4436] = 256'h29f463f3d3f188efb9ec3eeac9e898e8d0e901ec5fee8ef059f29cf381f4d8f4;
    inBuf[4437] = 256'h2df46ff2b9ef84ec00ea22e938ea22edf5f051f460f6bcf686f5abf312f242f1;
    inBuf[4438] = 256'ha1f1f6f296f405f6b9f646f6e5f4edf2c5f034efc6ee9cefc4f1d1f4eef770fa;
    inBuf[4439] = 256'hb7fb65fbd3f988f707f501f3c0f11cf10ff171f1fef1c0f2a3f35ff4eff442f5;
    inBuf[4440] = 256'h50f56ff5daf587f671f73cf860f8bcf75af672f4b4f2bef1d4f118f335f564f7;
    inBuf[4441] = 256'hfdf86bf95cf830f67af3c4f0adee66edb6ec90eceeecd6ed99ef50f29ff508f9;
    inBuf[4442] = 256'hcbfb23fddbfc0cfb09f88df43df191ee2bed6ded50ef9ff2a2f629fa3dfc34fc;
    inBuf[4443] = 256'hf4f945f649f209ef5aed59ed73ee05f05bf1f2f1e8f199f15af19cf17df2b8f3;
    inBuf[4444] = 256'h04f5f7f533f6c1f5d3f4b4f3f3f2e7f292f3edf4a0f623f827f978f9fff802f8;
    inBuf[4445] = 256'hcaf68df592f4e8f372f33af33bf36df3f7f3d5f4d5f5dbf6acf716f82df811f8;
    inBuf[4446] = 256'hcaf765f7b6f686f5e1f3faf13ef052ef88efcaf0caf2f8f4ccf61df8f7f882f9;
    inBuf[4447] = 256'hf5f94cfa71fa6bfa42fa09fad8f97af99df817f7f0f49cf2f2f09ff0eaf18ef4;
    inBuf[4448] = 256'hb8f773fa0dfc43fc5ffb01fab9f801f825f81af9b4fab4fcb8fe68008701f001;
    inBuf[4449] = 256'hb7010601f7ffb6fe6bfd2bfc2afb8dfa49fa47fa5cfa68fa96fa3bfb9afcc9fe;
    inBuf[4450] = 256'h6a01cc035505a405cc046003e901ab00bfff08ff78fe65fe46ff770106055809;
    inBuf[4451] = 256'h630d2b10e410500ffb0bc407b603e900f9fff8009203df06d109b70b3b0ca60b;
    inBuf[4452] = 256'hc80a4c0a8b0a750b5b0c7c0c870b7c09d90682041d0303034f049d066b09520c;
    inBuf[4453] = 256'hcb0e7c1051111e11f10f300e2e0c5f0a60097209a10ad00c650fab1114131613;
    inBuf[4454] = 256'ha211430f9b0c7f0ab9095b0a040c1a0eab0f2310920f420ed70c000ce10b570c;
    inBuf[4455] = 256'h2d0df90d9f0e580f281015111812c412cd1240122011ad0f560e3c0d870c6a0c;
    inBuf[4456] = 256'hc10c700d5b0e010f0e0f870e7b0d5e0cdb0b250c280d930eaa0f0010a80fd40e;
    inBuf[4457] = 256'hff0da40dac0dd90df80dc00d5d0d530dd40de70e55106c11aa111411ea0fd40e;
    inBuf[4458] = 256'h7d0eee0eda0fc91012118f10b20fe30e880eca0e290f100f300e5e0cfc09d107;
    inBuf[4459] = 256'h5f060706fc06e5085b0b030e3e109e11fc112d11780f960d1f0c9b0b540cdc0d;
    inBuf[4460] = 256'h820fac10ce100010ed0e230e120ed90ee70f95109d10ec0fe20e1f0ec20d9f0d;
    inBuf[4461] = 256'h6c0dac0c580bff0924093a09670a1b0cae0dca0e380f330f430f7c0fb80fc80f;
    inBuf[4462] = 256'h4a0f3a0e0e0d260ce60b8d0cb50dd20e800f4c0f280e870cc50a5409ae08cd08;
    inBuf[4463] = 256'h8c09cf0a340c800dbb0eb20f42106910df0f8e0ec70cd30a37099d082409950a;
    inBuf[4464] = 256'h800c000e640e980dce0bc10975085f088209870b880dda0e6d0f5d0f190f1a0f;
    inBuf[4465] = 256'h310fe70ee20dcd0bff087106f50420050807d109650cf80dff0dad0cd50a2109;
    inBuf[4466] = 256'h1a08090899086f096d0a650b630c980dcb0eb90f3610fd0f2b0f430e940d670d;
    inBuf[4467] = 256'hea0dc70e9a0f2b101d10550ffb0d130cee0924081e074107c4082e0bc60de10f;
    inBuf[4468] = 256'hd7109210860f1e0ed10cf30b620b040bee0a1a0ba50b9a0c930d250e090e040d;
    inBuf[4469] = 256'h5c0bca09e4082a09cc0a540d11105312631308138411350fb10c8f0a08093208;
    inBuf[4470] = 256'h08084308b6084e09d909490aa80acb0a8d0ad7097e08a906db04b403f5031006;
    inBuf[4471] = 256'ha909cc0d3d11c81203127a0f450ca30952081f084508ec0791068704cc025402;
    inBuf[4472] = 256'hac039b06110ac90ccb0db30cf0098506740390013f016302a1047d07580aa80c;
    inBuf[4473] = 256'hfb0df80da90c890a4608a3061b0691067a07220802081e07f9052e052b05ee05;
    inBuf[4474] = 256'hfd06d6073d0847085808c7088509210a0c0ad8089d06f603b701a7002401fe02;
    inBuf[4475] = 256'ha60564088d0aba0bd50bf70a5f0963075005750323029d010d0272038705d807;
    inBuf[4476] = 256'hdf09250b7d0b0a0b140ae908b7077a061e05ab035d029a01b301b4024804cf05;
    inBuf[4477] = 256'h9a064706e004db02e30098ff4cfffcff5301d3020104840449047d037602a401;
    inBuf[4478] = 256'h6501d401d102180455054506b9069306b8050a0488017ffe8cfb71f9dff820fa;
    inBuf[4479] = 256'hdafc31000f0389043c0459027cff75fcf7f969f8e9f74cf82ef92dfaf3fa53fb;
    inBuf[4480] = 256'h74fbaffb50fc7dfd0fff97009e01d8013e011800b3fe36fdbbfb50fa0af937f8;
    inBuf[4481] = 256'h2cf803f98ffa50fc9ffd0efe7cfd0cfc26fa3bf8a9f6dcf52cf6b6f75cfa85fd;
    inBuf[4482] = 256'h2e007601ec00bffedafb60f919f837f845f97cfa5dfbc8fbe9fb25fca1fc1efd;
    inBuf[4483] = 256'h55fd19fd65fc85fbc2fa2bfab5f93ff9b8f85df872f8fdf8d9f98cfa87faaaf9;
    inBuf[4484] = 256'h40f8cef610f671f6d8f7eaf91ffcebfd08ff44ff72fea5fc13fa25f7a4f44cf3;
    inBuf[4485] = 256'h6af3eaf42cf737f960fa6ffa99f97ff8abf741f72ff719f798f6a9f574f427f3;
    inBuf[4486] = 256'h19f277f134f159f1e8f1c8f2f7f358f5a1f6a6f738f82cf89ff7b0f673f52df4;
    inBuf[4487] = 256'h18f354f22ef2d5f227f4eff5baf7e4f80bf910f828f602f451f287f1e4f127f3;
    inBuf[4488] = 256'h9ff4b6f5fcf530f59df3ccf143f094ef04f064f15ff361f5bef62ef7b3f67df5;
    inBuf[4489] = 256'h18f402f36af27bf229f327f451f585f683f73ef8aff8bcf87af8e0f7bdf61df5;
    inBuf[4490] = 256'h1ff3f7f04defcfeebbef06f219f5e9f7b0f908faf6f81ef72df57ff355f2a0f1;
    inBuf[4491] = 256'h16f1b1f07df075f0dbf0e1f179f3a5f527f856fa98fb68fb83f968f6f3f2fdef;
    inBuf[4492] = 256'h52ee21eedceeedefcdf014f1eff0b6f092f0b6f020f18cf1f8f15bf28af2a2f2;
    inBuf[4493] = 256'hb1f29ff292f299f27af22af294f190f064ef70eedeede2ed56eebbeed9ee96ee;
    inBuf[4494] = 256'hf6ed75ed6dedcfed98ee97ef6df022f1c7f137f26bf22bf21ef167ef58ed51eb;
    inBuf[4495] = 256'h03ead2e9a0ea54ec8ceeaaf063f269f35ef35bf2b0f0caee7eed61ed76ee79f0;
    inBuf[4496] = 256'h9bf2cff3adf340f2f1efbced6fec4fec7ceda8ef28f288f440f6cbf628f68ff4;
    inBuf[4497] = 256'h6ff2acf0e5ef21f031f168f2f7f2b4f2e8f112f1f4f0d5f15ef322f586f613f7;
    inBuf[4498] = 256'hf3f660f678f577f456f3f1f195f0a1ef61ef33f0fff136f459f6dff76ff839f8;
    inBuf[4499] = 256'h77f756f62cf514f412f387f2b8f2adf35df54af7a6f8f0f8eff7e7f5b7f326f2;
    inBuf[4500] = 256'h95f114f21af3e3f317f4abf3ddf247f247f2dff202f461f5a2f6aff767f8a7f8;
    inBuf[4501] = 256'h78f8d2f7c2f6a8f5d6f47af4c7f48ff559f6cef6abf6daf5b3f499f3e5f2e8f2;
    inBuf[4502] = 256'h94f39bf4c3f5c0f659f7aaf7cff7dcf7fbf72df850f85df833f8a5f7baf67cf5;
    inBuf[4503] = 256'h11f4ddf23bf262f272f31ff5d3f60df865f8b9f76df61ef55af48ff4b5f563f7;
    inBuf[4504] = 256'h1af95afadefaccfa68fae1f956f9a6f895f729f6a1f469f309f3bef352f552f7;
    inBuf[4505] = 256'h23f943fa96fa31fa43f912f8cdf697f5c7f4a8f457f5bef671f8cff96dfa37fa;
    inBuf[4506] = 256'h77f9c3f884f8c1f83ff98ff95bf9bef816f8c4f717f8fdf810fae2fa1efba4fa;
    inBuf[4507] = 256'ha7f976f860f7adf673f6a2f62bf7f0f7d6f8e0f908fb2dfc26fdb1fd93fdd5fc;
    inBuf[4508] = 256'hb8fbaafa25fa50fafafab8fb08fcaefbf1fa55fa61fa5cfbfcfc94fe71ff23ff;
    inBuf[4509] = 256'hccfd0afc95fafbf964fa70fb89fc37fd31fd86fc81fb6dfa98f93ef979f961fa;
    inBuf[4510] = 256'hf4fbf8fd1500e001ed021a03870278015a008fff41ff85ff52007a01c402dc03;
    inBuf[4511] = 256'h5f0423042d03b901540087ff90ff7200de014c035c04cd048c04dc0308035002;
    inBuf[4512] = 256'h05024602f702fa030905d9056a06bf06d906d706aa062e068505ef04ca048e05;
    inBuf[4513] = 256'h41076c09780ba30c7d0c5f0bec09d908bc0881099e0a920be50b830be80a7f0a;
    inBuf[4514] = 256'h900a440b4a0c1f0d800d2b0d290cf50af1096e09bd09b80a030c6d0d9f0e700f;
    inBuf[4515] = 256'hff0f2810b90fb40efd0cc80ad708c107f4079e09260cb70ec210d511fb11be11;
    inBuf[4516] = 256'h5b11e3106810a30f840e700d980c280c420c7e0c7b0c420cde0ba00b0e0c210d;
    inBuf[4517] = 256'h920e23104d11da1115121412fa11fd11d6116211db105210ff0f2d108f10ca10;
    inBuf[4518] = 256'hc11042108d0f450f910f57104d11ad110811b00f1f0e1f0d720ded0efe100f13;
    inBuf[4519] = 256'h6114cb14c714931462144f14f0131e133612801171116412e4134c1530162416;
    inBuf[4520] = 256'h5b1592142a145c142915e8151e16c815e214d11338133113b513ae1491150b16;
    inBuf[4521] = 256'h2b16d215291594140b14911349130313c712e2123f13dc13be147015a4157215;
    inBuf[4522] = 256'hd7142314e1131414a814841528165e1659161316ac15641506157614dd132413;
    inBuf[4523] = 256'h6512e81183112011f010e61031112a12a0134115bb1666170217e9156014e812;
    inBuf[4524] = 256'h1812f0115312411365149215c31685177d17a616eb14b612f5103810dd10ef12;
    inBuf[4525] = 256'h9715dd171719b218d0164b14e3115b104f10831172139615181788170d17c215;
    inBuf[4526] = 256'h0d1498129b114711da111213a3144a165d1771179f160d155a137612bd122b14;
    inBuf[4527] = 256'h7416a418f219231a211951177315d613b312421242128e123313df136014bb14;
    inBuf[4528] = 256'hab14261473139912c31146111e1158112012321350145515c41562155c14c112;
    inBuf[4529] = 256'heb10750f930e710e3a0f9d104212dd13d414d014e0131712f70f4a0e6f0d9c0d;
    inBuf[4530] = 256'hce0e6a10db11cc12dc121712dc10590fd60da50cc10b430b5e0b020c310de80e;
    inBuf[4531] = 256'ha210d1110112b810090eb00a9007ad05b7057407250acb0c510e560e320d6f0b;
    inBuf[4532] = 256'hba098b08c4072f07ba0660066c06320794083b0aaa0b490cec0bc90a25096a07;
    inBuf[4533] = 256'he70597048903e902d4027403d2049b065f08a7090f0a9b098f082c07c7059504;
    inBuf[4534] = 256'h9103c2023e0210024f02e9028a03d3036a032402460063fe1afdf8fc14fe0700;
    inBuf[4535] = 256'h2e02d1036704d6035f027700a6fe55fdc1fc09fd0ffe8fff3b01a1025b033d03;
    inBuf[4536] = 256'h4802b700f4fe58fd2cfc91fb6ffb9afbe1fbfdfbc9fb43fb73fa90f9ddf879f8;
    inBuf[4537] = 256'h71f8b7f810f94ef953f90af98bf803f88ff76bf7c3f783f891f9affa6cfb85fb;
    inBuf[4538] = 256'he6fa99f9fbf77bf668f50df57af56af694f78cf8c6f815f891f686f4a3f294f1;
    inBuf[4539] = 256'h99f1abf257f4d4f59df678f66bf5f2f389f263f1b7f08bf0a9f016f1d3f1aaf2;
    inBuf[4540] = 256'h8af34ef4a8f49df44af4bef343f3f9f2b0f25df2e7f119f12ff076ef05ef17ef;
    inBuf[4541] = 256'hafef6af012f16cf132f190f0beefd0ee20eeddede0ed37eeccee48efa3efd5ef;
    inBuf[4542] = 256'haeef5eef09ef98ee38eef9edaaed6ced47ed07edd0ecabec66ec3aec4eec7eec;
    inBuf[4543] = 256'he5ec6beda6ed7aedd4ec8eeb0ceaade894e732e7b5e7d5e87dea56ecb2ed55ee;
    inBuf[4544] = 256'h21eefaec6ceb0bea11e9e0e873e94fea46eb23ec8fecb7ecb3ec49eca6ebdcea;
    inBuf[4545] = 256'hc3e9ace8dee755e75ae7f8e7d4e8dce9c2eaf4ea65ea1ae90ee7f0e467e3bae2;
    inBuf[4546] = 256'h51e314e546e777e931ebf4ebfeeb95ebbdead3e9f8e808e86ee77fe730e8ade9;
    inBuf[4547] = 256'ha5eb35edf6edb4ed65ecccea8ee9c3e884e86ee8d6e7d6e6c2e5d7e4afe463e5;
    inBuf[4548] = 256'h58e641e7cce7b0e769e75fe788e7fce772e856e8c3e7f2e605e69ae5f4e5c4e6;
    inBuf[4549] = 256'hfee75be958ea0aeb86eba9ebc2ebe7ebcfeb96eb2deb4cea40e945e859e7eae6;
    inBuf[4550] = 256'h1ae794e74ee8ffe820e9bbe8eee7cee6f9e5d9e55fe6a0e741e986ea3feb55eb;
    inBuf[4551] = 256'hb0ead6e927e995e856e85fe866e89ee81ee9b4e97bea4eebc3ebf4ebf6ebb3eb;
    inBuf[4552] = 256'h81eb78eb4ceb16ebd8ea73ea3dea67eac3ea5bebf2eb15ecd9eb5deba8ea38ea;
    inBuf[4553] = 256'h50eac1ea90eb83ec25ed7eeda2ed8aed93eddfed2dee7eeeafee7cee1deeb5ed;
    inBuf[4554] = 256'h24ed92ecf6eb1aeb50eaf3e92aea3eeb05edd1ee2df0b5f037f037ef47eea1ed;
    inBuf[4555] = 256'h8cede8ed3cee7deeb7eeeaee60ef1df0cdf057f1a1f189f15bf148f13af148f1;
    inBuf[4556] = 256'h61f156f158f186f1bbf102f23af21ff2caf159f1c4f02bf081ef9beec1ed56ed;
    inBuf[4557] = 256'ha5ed0bef57f1bcf376f5e8f5e1f40ef361f196f028f1dcf2ebf4b5f6c3f7e7f7;
    inBuf[4558] = 256'h7ff7f9f697f6acf63df70af8e3f876f96cf9c8f8b6f783f6b2f586f5e8f5b2f6;
    inBuf[4559] = 256'h8af720f886f8def83bf9acf9fff9dbf927f9f7f7a1f6bcf5b6f5abf677f88cfa;
    inBuf[4560] = 256'h39fc0afdcefcbdfb7dfabaf9e8f922fbf8fcb7fecfff01008eff16ff1affbfff;
    inBuf[4561] = 256'hba0061012601f3ff33feb0fc2efcf6fcc5fee7008c023303d702cf01b100f8ff;
    inBuf[4562] = 256'hc4fffdff5b0090008b006800590099003201f0019902f002db0298027c02cb02;
    inBuf[4563] = 256'hae03f304310621079807af07c8072408c7088909fd09c409e3088e0730066705;
    inBuf[4564] = 256'h8905a506a8081d0b660d000f650f600e560ce109cc07ed06710701090e0bc60c;
    inBuf[4565] = 256'ha80dca0d660dd80c8b0c800c9e0cfd0c8c0d450e370f0e107a1081102c10d00f;
    inBuf[4566] = 256'hfd0fb910b1117a1272126111c90f400e6c0dd30d2f0ff110ae12e9138514dc14;
    inBuf[4567] = 256'h081519153a153215e81493142b14be138f1381138813c813061419140c14a113;
    inBuf[4568] = 256'hd712131280115e11031234139a140616fb1642170e175b164d15441439133812;
    inBuf[4569] = 256'h8e1132114011101285137815d217f719631bf51b791b281ab9188717d916e816;
    inBuf[4570] = 256'h38175017121746162415521409145c144c15371691164b164a15ee130713e212;
    inBuf[4571] = 256'h9a132a15d91604188618311849177e16fa15ce1515166c16a8160d1788171a18;
    inBuf[4572] = 256'hdd1859193f19bf18ec172a171a179c174f18e018a7187b17ef1575149213c013;
    inBuf[4573] = 256'ha414bf15d9167d1792177217061748167a15841494132f135a13031426153216;
    inBuf[4574] = 256'hcd161d171717e316e016d61693163716a3150715f4146a154c1687178518eb18;
    inBuf[4575] = 256'he1185e189117e8163d167415c714191489138313dd135814e114001596141414;
    inBuf[4576] = 256'ha31381130114c4146b15f0150f16d915bb159915541505156b1497130f13f212;
    inBuf[4577] = 256'h51133e141f157f156315b214c3135013841369140916c6171819c9196a19f517;
    inBuf[4578] = 256'hf215b913da110b114a115912ed133915bb158515971453136112e011d3114a12;
    inBuf[4579] = 256'hd1121c133c130813a3128112a2120913c1134a144114a6135a12ab10490f7e0e;
    inBuf[4580] = 256'h820e7a0feb106612c313a51409153c153215f714b91441148913d4122212a111;
    inBuf[4581] = 256'h9911d81121124612c9118310c10ec30c150b5f0aaf0ae50bbd0d880fd6109111;
    inBuf[4582] = 256'h9b111e117110980fa80ed80d1d0d990c8c0cd60c5e0d170eb40e1f0f790fac0f;
    inBuf[4583] = 256'hb60f960ffd0ed70d610cdd0ad209c609af0a3a0cda0dc10e8a0e5b0d910bda09;
    inBuf[4584] = 256'hd808a8081d09dc09560a500ae5093f09b9089d08d4082a095909ff080608aa06;
    inBuf[4585] = 256'h3f054c0442042905c6069b08f109560ab50941088a062905670449048a04a904;
    inBuf[4586] = 256'h5d04a403b90216021d02db0219045b050e06e705ed046803dc01bb0035004800;
    inBuf[4587] = 256'hb80038019701c401c901ce01e401fd01f7019501a70035ff77fdd6fbd6fac1fa;
    inBuf[4588] = 256'h99fb0bfd81fe6eff89ffd4feacfd92fce5fbd0fb4efc1bfdf2fd9bfee1feb2fe;
    inBuf[4589] = 256'h1afe28fd14fc1ffb66faf9f9d3f9cbf9daf916fa87fa3dfb1afcbffcd4fc29fc;
    inBuf[4590] = 256'hb8fae1f829f7e4f550f566f5d3f561f6e7f633f746f72af7d6f676f63ef63ff6;
    inBuf[4591] = 256'h94f623f792f7b0f770f7e0f669f668f6e4f6c0f79cf8ecf87ef865f7d7f556f4;
    inBuf[4592] = 256'h4cf3cbf2dcf250f3bdf3f1f3c9f31df323f226f14ff0ebef10f077f0f0f044f1;
    inBuf[4593] = 256'h35f1f5f0cbf0d0f031f1def177f2e5f228f331f33bf355f336f3c5f2f8f1d3f0;
    inBuf[4594] = 256'hdeef9bef1ef05bf1d3f2b5f3aef3c4f227f179ef23ee12ed41ec99ebfdead2ea;
    inBuf[4595] = 256'h76ebdcece9ee1af19af213f374f2cef0b9eebeec11eb18ea08eab9ea2eec21ee;
    inBuf[4596] = 256'hedef3bf1caf16df19bf0d3ef40ef1def44ef27efabeed9edc8ec0bec05ec99ec;
    inBuf[4597] = 256'haaedccee4bef00eff7ed47ec90ea51e9a2e8c2e8a0e9ccea2bec89ed7eee0fef;
    inBuf[4598] = 256'h32efadeeb8ed7fecfaea8fe984e8dae7e5e7bfe81beae3ebc1ed16efc2efbaef;
    inBuf[4599] = 256'hf7eefced2fed8dec34ece9eb27ebf3e984e81be780e62fe7f5e883eb0bee76ef;
    inBuf[4600] = 256'h6def06eea5eb55e9dee75ee7e3e70ae92eea45eb5bec4eed42ee05ef07ef37ee;
    inBuf[4601] = 256'hafeca3eae0e800e814e832e9fbeab1ec04eea8ee48ee2aeda9eb09ea04e90ee9;
    inBuf[4602] = 256'h11eaf1eb19ee98ef10f066efbaeddeeb88eaf6e96beaa7ebf8ec0aee94ee53ee;
    inBuf[4603] = 256'habed06ed94ecbfec88ed78ee5cefedefdeef75efedee38ee7deda4ec6aeb1fea;
    inBuf[4604] = 256'h2de9e0e8b5e9a0ebeeed0ff061f16af184f037efe6ed26ed1fed8ded69ee87ef;
    inBuf[4605] = 256'h89f067f1f2f1d2f130f144f03defa5eeb3ee24efcaef3df008f053ef6bee8fed;
    inBuf[4606] = 256'h46edb7ed95eeabef95f0d9f086f0c6efc1eefbedbfedfaedb9eec3efaff071f1;
    inBuf[4607] = 256'hf5f117f207f2d6f168f1f4f09af060f08ef039f128f247f351f4dcf4e7f475f4;
    inBuf[4608] = 256'h86f374f27ff1aff03ff034f05ef0c6f051f1c6f13af2adf205f360f3b0f3b4f3;
    inBuf[4609] = 256'h65f3b3f29af182f0d3efc7ef9df028f2e1f367f564f6a5f671f60bf690f532f5;
    inBuf[4610] = 256'hf1f4b2f4a4f4e2f45ff517f6c7f60ef7e3f65ff6aef531f505f5fcf401f5f9f4;
    inBuf[4611] = 256'he5f414f5b6f5b3f6daf7c1f800f99bf8c3f7bdf6eaf570f53bf54df59ff527f6;
    inBuf[4612] = 256'h02f724f858f97cfa59fbc2fbc1fb66fbc8fa25faaef97bf9a4f90bfa6dfaaafa;
    inBuf[4613] = 256'haffa95faa2fafdfa92fb28fc6cfc2cfc9bfb20fb21fbd9fb0dfd33fecdfe9afe;
    inBuf[4614] = 256'hc5fddffc76fcd0fcd4fd02ffc2ffbdffeffeb2fd97fc13fc57fc4efda0feefff;
    inBuf[4615] = 256'h0501d201700202038303d003b5030b03e3018c006affdbfe06ffcaffdf00fb01;
    inBuf[4616] = 256'hea02ae035a04f7047d05c2059905fe041504240383026502c9028e0374044105;
    inBuf[4617] = 256'he6056006b406f1060607df06880610069c0565057805c7053a06a206e4061807;
    inBuf[4618] = 256'h5107a5072b08c4084409950997094609c7082d088d071a07ea061b07da071609;
    inBuf[4619] = 256'h990a1d0c250d540da90c560bd209c0086508b80876091c0a580a4d0a3f0a8d0a;
    inBuf[4620] = 256'h760bb00cb00d0e0e870d5c0c410bb50af00ad30bc60c3e0d200d810cc00b5b0b;
    inBuf[4621] = 256'h6a0bd90b980c660d230edd0e630f890f520fab0ec20d060da30ca50c0c0d830d;
    inBuf[4622] = 256'hd50d1e0e5f0eaf0e2f0f9e0fbf0f940f080f460eb30d660d690dd30d6a0e020f;
    inBuf[4623] = 256'h9c0ffb0f0210d10f630fe30eae0ec40e140f950fef0ff90fe00fae0f860fa30f;
    inBuf[4624] = 256'hd50ff50f11100c10f90f1e106510b11006112011ea1098102410a30f540f220f;
    inBuf[4625] = 256'h0c0f390f760fa10fc60fb30f6b0f3f0f3b0f6f0ffd0f97100211511169116511;
    inBuf[4626] = 256'h9611da110e1238121512a7114311f210cb10fe104c119111e711201232124712;
    inBuf[4627] = 256'h2d12d81181111a11bc10ad10c410e51021113d11301138113b11371151115011;
    inBuf[4628] = 256'h23110411e410df103f11dc1195126e130b1442144114f5138513531351137813;
    inBuf[4629] = 256'hd9131d141114d61347137e12d6114811e510e710211184113012e1126d13e113;
    inBuf[4630] = 256'hf0138c13f7122f126211ee10bb10bf1017118411fa11ae1276133b1408157d15;
    inBuf[4631] = 256'h6b15f8141914021324127c110b11f510fb10161185112912f612f613b914f714;
    inBuf[4632] = 256'hb714d3137e1241114a10db0f3b1021113f126013fb13d91335132c121e118c10;
    inBuf[4633] = 256'h63107a10ba10c2108f108b10db10a211e7121114961450141d136311e40ff60e;
    inBuf[4634] = 256'hc90e6e0f6e106d115612dc12e6129412c01187105d0f790e280eb10ebe0fe410;
    inBuf[4635] = 256'he01145120d129a11091189104510f90f810ffa0e530eb40d700d780dcb0d7b0e;
    inBuf[4636] = 256'h3e0fe50f65107010f40f2c0f2d0e410dcd0cc50c0f0d920df00d070efe0dd30d;
    inBuf[4637] = 256'ha60daa0db80dc00dd70dd80dc50dba0d870d1a0d8c0ccf0b0d0b990a750aa70a;
    inBuf[4638] = 256'h300bbe0b1d0c480c180c970bfe0a4e0aa4093909050917098b09330ae60a840b;
    inBuf[4639] = 256'hb50b500b730a3409f0072007eb06550740083509e009270af2096909d5084608;
    inBuf[4640] = 256'hd5079f078e07a107de0716082d081c08cb074f07dc067906340618060506fb05;
    inBuf[4641] = 256'h0f062d0649064f060a067705ca043e041e049304600525068406330648052404;
    inBuf[4642] = 256'h24039902a1020c03a1033704a804f10418050805b70427045f038b02e0017201;
    inBuf[4643] = 256'h4d0164019301c801ff0130025c027d027f0262023002f601c3018d012d018000;
    inBuf[4644] = 256'h7aff43fe3afdcbfc39fd7afe1f0081011002830107002afe8afc9cfb84fb08fc;
    inBuf[4645] = 256'hd0fc9cfd4dfef5feacff5f00d800d4001d00c6fe27fda7fbaffa70fac7fa70fb;
    inBuf[4646] = 256'h18fc70fc63fcfffb5dfbb0fa27fad0f9baf9e0f91cfa5dfa99fab9fac9facefa;
    inBuf[4647] = 256'ha9fa54fac5f9edf8fff73cf7ccf6e1f67bf755f836f9e0f911fad0f93ef971f8;
    inBuf[4648] = 256'hacf71bf7b8f694f6a4f6b9f6d9f606f728f750f776f766f718f788f6a3f5a2f4;
    inBuf[4649] = 256'hb7f3e8f262f22cf223f258f2cbf253f3f2f389f4ccf4b7f44cf48ef3d4f266f2;
    inBuf[4650] = 256'h49f295f21ef373f36bf3edf2f3f1e8f038f00bf090f099f195f234f332f367f2;
    inBuf[4651] = 256'h36f109f013efa2eeb2eeeeee42ef96efbcefe6ef25f04df066f05af0eaef3def;
    inBuf[4652] = 256'h73ee8bedd8ec89ec8fec1bed20ee3def43f0d7f086f070efe3ed33ec18ebf4ea;
    inBuf[4653] = 256'h9febebec59ee3bef79ef1eef3cee4fed9eec15ecdcebe2ebe0ebeeeb08ecf8eb;
    inBuf[4654] = 256'heaebe9ebcaebbeebcbebbaebafebb0eb8feb87ebaaebcaeb0eec6eeca0ecc0ec;
    inBuf[4655] = 256'hc2ec68ecddeb2feb44ea6fe9e1e88ae8aae836e9d1e973eae9eaddea81eafbe9;
    inBuf[4656] = 256'h4ee9e1e8dbe80be988e932eab0ea20eb7beb84eb60eb08eb45ea67e9a8e816e8;
    inBuf[4657] = 256'h13e8abe87fe978ea4eeb92eb69ebeaea0cea3ae9ade857e87ae80be9a8e94dea;
    inBuf[4658] = 256'hcdead6eaa4ea56ead4e966e91be9c4e8a0e8c3e8fee879e917ea7fead0ea17eb;
    inBuf[4659] = 256'h35eb72ebccebebebdeeb9ceb06eb87ea54ea47ea82eae1ea1ceb6eebfbeb9bec;
    inBuf[4660] = 256'h68ed1dee37eebfedd1ec8eeb8cea0eeae5e916ea6bea92eac6ea27eb98eb3fec;
    inBuf[4661] = 256'hfbec6aeda6edb3ed72ed2eedfaecaeec8aec9eecc3ec26edaeed02ee38ee56ee;
    inBuf[4662] = 256'h46ee5ceea5eed2eedeeea1eeefed30edbdeca9ec31ed24eeffeea5eff2efbeef;
    inBuf[4663] = 256'h56efd8ee2aee88ed11edc2ecefeca5ed90ee8fef48f054f0ddef22ef53eef6ed;
    inBuf[4664] = 256'h3eee00ef33f084f16ff2d6f2a0f2c0f1aef0ceef46ef56efdaef5cf0bcf0e1f0;
    inBuf[4665] = 256'hc6f0d7f052f11bf223f30bf44df4def3d1f24df1e6ef06efd2ee82efeef098f2;
    inBuf[4666] = 256'h27f421f519f52ff4b9f224f12df03df040f107f304f583f641f72af753f63af5;
    inBuf[4667] = 256'h3df47df32af333f35ef3b0f31cf485f4fef477f5bef5dbf5d0f59bf580f5a3f5;
    inBuf[4668] = 256'hfdf598f645f7b5f7cef77af7aef6b0f5bdf402f4c3f313f4cff4e8f527f74cf8;
    inBuf[4669] = 256'h49f906fa61fa5ffaf0f90cf9ebf7d5f618f617f6e8f655f806fa78fb3cfc38fc;
    inBuf[4670] = 256'h86fb67fa43f95ef8daf7d1f73df805f915fa3afb33fcd5fc06fdcefc66fc06fc;
    inBuf[4671] = 256'hcefbcafbdffbebfbeefbfcfb3afcccfca4fd90fe51ffb2ffaeff72ff37ff29ff;
    inBuf[4672] = 256'h4fff7fff8aff56ffe6fe71fe36fe5ffefbfeecfff300d80168028b025402e901;
    inBuf[4673] = 256'h7f0151017a01f101a3025e03f7036a04ae04c704c504a10457040804c903b503;
    inBuf[4674] = 256'hee036204eb047905f4055c06d9066407e40741084608e5075007b40643062d06;
    inBuf[4675] = 256'h57069b06f5064f07b4074d080b09cd09830af40a090be80a9b0a400a0c0aff09;
    inBuf[4676] = 256'h1a0a7e0a130bc20b8c0c340d8d0da20d5f0ddc0c670c160c030c570ce70c890d;
    inBuf[4677] = 256'h340ea60ec50eb40e730e200e030e140e450e9f0ee10eea0ee20ec80ec00e180f;
    inBuf[4678] = 256'hbe0f951096116c12e3121013d4123b129311e51059104510a010571165125f13;
    inBuf[4679] = 256'hf1132214da134e13fb12f7124713f0137f14a2146314ad13b9121112da112b12;
    inBuf[4680] = 256'h1c133c142115ad159315e31411144c13cf12ec126f1329141d15fb15a2163917;
    inBuf[4681] = 256'h8f1798178f175617fb16c71698165c163216da154715c614541412145414e414;
    inBuf[4682] = 256'h9715721615175b1776174817e116971653161b162e1654167516bc16ee160717;
    inBuf[4683] = 256'h4f17a017e9174a18661814188d17c9160216bd15ed15821682176f18fd184119;
    inBuf[4684] = 256'h06196118c4173417d816fe165f17be1718180c1892171817b2169216fa168617;
    inBuf[4685] = 256'he51720180318b717b717ee173e189f1899180e186317be166e16d816b0179d18;
    inBuf[4686] = 256'h7e19da199519071934184e17b8164e1604160b1623163c169116e9162e178217;
    inBuf[4687] = 256'h93174817e0164e16c415b415021692165f17ea17f817be17321791164a163a16;
    inBuf[4688] = 256'h42166a165616f51593152215b81496148014631478149a14d4145f15ee154b16;
    inBuf[4689] = 256'h7e163d169115db141d147a1336131b131c136513c01318148614b41480141c14;
    inBuf[4690] = 256'h7913cc127e127612a3120b13551368137f1385138513a51395133313ac12f611;
    inBuf[4691] = 256'h4f111d1144119d110a121712a411fd104310c80fe40f5a10e6105b115311c710;
    inBuf[4692] = 256'h1010510fcb0ec50e020f530fa60fb30f790f3d0fff0edf0e040f2f0f360f170f;
    inBuf[4693] = 256'h970ec40deb0c1e0c990b9e0b080cae0c6a0dc80d920dde0cb80b7e0ab2097509;
    inBuf[4694] = 256'hce099f0a640bc50bb10b160b340a6d09d30872084d082908f907db07c107bc07;
    inBuf[4695] = 256'hdd07f507f607ee07d207bb07c907d607c7078c0700073f068f051005e8041a05;
    inBuf[4696] = 256'h5e057d055d05e8044e04d3038d038c03c003e503d7038f0305036502e5019801;
    inBuf[4697] = 256'h9901ed016902ec024b034c03e302200224014200c9ffdfff88008a016e02d502;
    inBuf[4698] = 256'h810273010b00c5fefffdecfd5efeecfe39ff10ff7cfed0fd57fd33fd5efd99fd;
    inBuf[4699] = 256'ha8fd7efd30fde8fcd9fcfdfc2cfd42fd19fdb7fc4efc00fcdcfbdbfbc2fb63fb;
    inBuf[4700] = 256'hc1faf1f93bf9f3f833f9e9f9dafa92fbc2fb57fb5ffa32f93df8b6f7b7f728f8;
    inBuf[4701] = 256'hacf8fef8f7f87ef8bef7fdf65ef607f605f621f63af63bf601f6aef57cf580f5;
    inBuf[4702] = 256'he0f59df66bf70bf84bf8edf712f706f6fbf43ff4fcf302f437f47af490f485f4;
    inBuf[4703] = 256'h74f449f414f4dbf373f3fbf29ff265f27ef2f2f276f3dcf3f8f390f3d6f21df2;
    inBuf[4704] = 256'h91f180f1f9f1a4f246f3a1f36bf3d1f222f283f140f16af1aff1eaf1fef1b8f1;
    inBuf[4705] = 256'h54f114f1f2f00ff15bf17ff175f146f1e1f08af06df061f070f084f053f0f3ef;
    inBuf[4706] = 256'h83effbeea1eea1eecdee2fefa9efdbefc9ef80eff1ee78ee5bee89ee17efdbef;
    inBuf[4707] = 256'h57f070f020f059ef8cee19eeffed5eee07ef79ef97ef57ef9ceec1ed09ed67ec;
    inBuf[4708] = 256'h0fec09ec16ec54ecc7ec31edaeed38ee8aeec2eee5eebfee7dee33eebaed48ed;
    inBuf[4709] = 256'hf9eca2ec73ec78ec7deca9ec01ed44ed87edc0eda9ed70ed36ede5ecc9ecf9ec;
    inBuf[4710] = 256'h39ed97edf8ed06eedaed7fedd6ec31ecc5eb80eb9beb0cec75ecd0ec01edd1ec;
    inBuf[4711] = 256'h89ec64ec55ec97ec1eed89edd4edeaed96ed21edb9ec4fec23ec3fec61eca3ec;
    inBuf[4712] = 256'hfaec28ed55ed84ed7ced67ed4ded02edc2eca5ec80ec7eec91ec70ec3becffeb;
    inBuf[4713] = 256'ha9eb92ebe6eb7aec5bed47eebbeea7ee09eee7ecd5eb40eb3cebf3eb22ed32ee;
    inBuf[4714] = 256'hf4ee44ef02ef92ee34eed9edaced9fed6ded41ed29ed0aed19ed5bed98edf4ed;
    inBuf[4715] = 256'h65eeb2eef6ee21effceebdee82ee47ee52eea7eefbee47ef60ef0def92ee29ee;
    inBuf[4716] = 256'he9ed26eee4eed6efe4f0cbf134f237f2e4f135f17cf0e1ef5def2eef5fefc4ef;
    inBuf[4717] = 256'h6bf028f1a6f1e5f1d8f16ff1fbf0b1f097f0e3f084f12ff2d4f242f340f3f8f2;
    inBuf[4718] = 256'h89f207f2c5f1dbf122f29cf216f349f345f314f3bcf28ef2aff216f3daf3ccf4;
    inBuf[4719] = 256'h92f512f627f6bdf521f589f40cf4d8f3daf3e1f3fbf329f45ff4bff430f575f5;
    inBuf[4720] = 256'h8ff57ef557f574f5f6f5bcf6a1f74bf864f8fdf73ff767f6dbf5c1f50bf6b4f6;
    inBuf[4721] = 256'h8df756f8fcf859f94bf9f2f86df8e6f7aaf7d2f74af8fef8b4f934fa80fa9afa;
    inBuf[4722] = 256'h8afa75fa5bfa31fa0ffaf6f9ecf90afa47fa86fac2faecfa01fb28fb6ffbd5fb;
    inBuf[4723] = 256'h5afcdbfc34fd64fd65fd3ffd0efdd9fca7fc90fc97fcb9fcf8fc39fd68fd91fd;
    inBuf[4724] = 256'hc7fd2bfed9feb7ff7f00e5009e00a8ff4efefbfc23fc13fcc1fceffd46ff6600;
    inBuf[4725] = 256'h190158013101d400750034002a005900a700ff004f018401a001a70197017a01;
    inBuf[4726] = 256'h5d01460146015b01680156011401aa005d007b0038019e025b04e305bc069c06;
    inBuf[4727] = 256'h8f050c049b02ab017401d30171020a036d039503b103e4033404ab0428059105;
    inBuf[4728] = 256'he905280647064f062f06dc0573050805b504a404d1042805aa053b06c9065b07;
    inBuf[4729] = 256'hd30711081108c2073207a5064606380698064107fb07a80816092f090f09bf08;
    inBuf[4730] = 256'h5208f607b2078c07a207e6074a08d5086109cc09180a270af709b5096f093b09;
    inBuf[4731] = 256'h45097d09c809220a570a4a0a120ab309500934097009020ae20ac00b4f0c7e0c;
    inBuf[4732] = 256'h350c950bf90a840a4e0a6b0aa60ad30af50af30ad50ad00ade0a020b570bba0b;
    inBuf[4733] = 256'h150c740cb10cb70ca00c590cef0b9f0b6f0b720bc90b450cb80c140d220ddb0c;
    inBuf[4734] = 256'h770c070cb00ba80bda0b310cb60c3b0da60d030e240ef60d950dfc0c4d0cdb0b;
    inBuf[4735] = 256'hb40be00b6d0c0f0d8b0ddc0ddf0dab0d8b0d8d0db60d160e6a0e7f0e620efe0d;
    inBuf[4736] = 256'h6b0df90cb10c9f0ce20c490db10d260e770e9a0eb30eb00e960e8a0e6c0e300e;
    inBuf[4737] = 256'hf50da90d5e0d4e0d680d9b0dec0d200e200e1a0e090efb0d110e150ee50d950d;
    inBuf[4738] = 256'h220dbc0cc10c350d030e100fea0f451025107f0f860ea40df60c970ca50ceb0c;
    inBuf[4739] = 256'h3f0da50deb0d030e130e080ee90de60dec0df70d1b0e290e060ec80d5d0dda0c;
    inBuf[4740] = 256'h820c590c670cca0c510dd90d600eac0ea30e610edf0d410dd70ca80cb50c010d;
    inBuf[4741] = 256'h490d660d6f0d5f0d500d730da40dbd0dbb0d760df80c8a0c3e0c2e0c7c0cf60c;
    inBuf[4742] = 256'h6c0dd30def0dab0d2e0d7c0cbb0b350bef0aed0a440bc30b470cd40c380d5e0d;
    inBuf[4743] = 256'h590d180dae0c600c3a0c490c9e0cf60c1b0d060d9d0cfa0b6e0b0f0bed0a1c0b;
    inBuf[4744] = 256'h680bae0bf40b1a0c1b0c100cdf0b810b1c0bb20a5f0a550a7f0abf0a050b1a0b;
    inBuf[4745] = 256'hf00abb0a890a760aa00ada0afa0a000bd70a920a6c0a650a7b0ab40ae40af30a;
    inBuf[4746] = 256'hf00ac80a7c0a2d0ad30976093b09160906091a0934094309550953093c092f09;
    inBuf[4747] = 256'h2409250948096e0975095209e6083e089e073207220788073208e1087109b209;
    inBuf[4748] = 256'ha00961090109940842080a08f0070308200823080408aa072607b60676067806;
    inBuf[4749] = 256'hc2061b074e074b0700078c0632060e063506a6062c079007bb0795072f07b706;
    inBuf[4750] = 256'h4306e0059c055f052405030506053c05ae0534069c06ca069f062b06a5053205;
    inBuf[4751] = 256'hf104ef0403050205d8047804ff03a6038c03bd032d04a304ee04fd04c8046a04;
    inBuf[4752] = 256'h0c04bf038b037a0381039e03d3030b0430043104fc0398032903c80291029302;
    inBuf[4753] = 256'hbc02fd0247038603b003bf03a7036503020387020d02ae01770170019401cc01;
    inBuf[4754] = 256'h02021f021502e801af017b015c01550158015e016c018e01d30139029a02c002;
    inBuf[4755] = 256'h7e02c801d000ecff72ff96ff45002c01e9012b02db0124015100acff62ff6bff;
    inBuf[4756] = 256'ha1ffdbfff7ffefffd1ffa5ff6fff33fff0feb6fea3fec9fe2bffaeff16003000;
    inBuf[4757] = 256'he6ff43ff7dfee0fd9bfdc0fd40fee0fe6affb9ffafff54ffc7fe23fe8afd1cfd;
    inBuf[4758] = 256'hd5fcb3fcabfca3fc97fc8dfc85fc91fcc0fc07fd5dfdadfdcbfd9ffd27fd66fc;
    inBuf[4759] = 256'h8afbcefa57fa45fa9ffa3efbfefbbdfc46fd83fd6bfdeffc2dfc56fb8dfa05fa;
    inBuf[4760] = 256'hdaf9f1f932fa7dfaabfabffad0fadbfaeefa05fbf7fab7fa44fa9bf9e5f854f8;
    inBuf[4761] = 256'hfff704f868f8faf898f91efa5bfa50fa0ffa98f90df98df81bf8d5f7d0f7f4f7;
    inBuf[4762] = 256'h36f87cf88ff86cf82df8e1f7bef7def71ef85ef870f81ff87cf7bff60df6a9f5;
    inBuf[4763] = 256'hb5f50af689f60af750f761f74ff712f7c2f669f6e9f557f5d6f477f46cf4c8f4;
    inBuf[4764] = 256'h53f5e7f552f65cf61ff6cff583f566f578f574f53ef5c9f410f45df3fbf200f3;
    inBuf[4765] = 256'h82f362f43cf5d9f510f6baf507f535f45ef3bdf26df251f274f2d0f239f3abf3;
    inBuf[4766] = 256'h11f42ff40af4aef31bf391f247f238f275f2e9f24ff399f3c0f3a9f379f349f3;
    inBuf[4767] = 256'h07f3c9f298f255f222f213f213f235f273f29af2aef2b1f28bf262f24bf228f2;
    inBuf[4768] = 256'h0df201f2e6f1dcf1f3f10ff23bf26df274f25ff240f208f2e2f1dff1dcf1e1f1;
    inBuf[4769] = 256'he6f1c5f1a3f19ef1aef1f7f16ff2cff201f3eaf26ef2caf140f1e2f0dbf021f1;
    inBuf[4770] = 256'h6df1b2f1ecf104f223f256f26ff26cf244f2dff179f141f134f169f1c7f10af2;
    inBuf[4771] = 256'h2ef236f215f201f217f23bf279f2bdf2caf2a3f24cf2bdf13df105f11df1a9f1;
    inBuf[4772] = 256'h8ef270f320f46df426f47bf3a7f2cdf13cf115f136f1a3f13df2caf24ff3c4f3;
    inBuf[4773] = 256'h04f41ef40ef4b9f348f3e0f28df286f2d3f23df3b4f312f42af41bf405f4ecf3;
    inBuf[4774] = 256'hf5f320f43df451f454f433f416f419f42cf466f4bdf401f537f556f547f52af5;
    inBuf[4775] = 256'h10f5e9f4d1f4cef4caf4e1f419f554f59ff5ebf512f627f635f635f642f65cf6;
    inBuf[4776] = 256'h61f658f63ef609f6e4f5e6f508f65df6dbf655f7c7f71ff83cf82ff801f8b1f7;
    inBuf[4777] = 256'h6cf749f740f765f7aaf7ebf728f857f867f86ff87df888f8a9f8daf8fdf80ff9;
    inBuf[4778] = 256'h07f9d7f8a4f889f891f8d6f84ff9d2f955fac1fa00fb20fb28fb0cfbdefaa3fa;
    inBuf[4779] = 256'h58fa21fa12fa31fa8ffa19fba6fb20fc69fc65fc2cfcd8fb85fb5ffb76fbbafb;
    inBuf[4780] = 256'h23fc8efcd7fcf9fcf5fcd6fcbefcc2fce2fc20fd63fd8afd8ffd74fd48fd35fd;
    inBuf[4781] = 256'h50fd9efd1cfeaafe26ff7fffa9ffa0ff74ff31ffe5feadfe94fea4fee0fe35ff;
    inBuf[4782] = 256'h8effe0ff1b003b00450038001400e8ffbeffacffcaff17008900060169019a01;
    inBuf[4783] = 256'h9601680131011101160147019901ee01320258025c024f02440245025f028f02;
    inBuf[4784] = 256'hc402fa02250339033e0334031c030703fd02ff0217033e036a039f03d8031004;
    inBuf[4785] = 256'h4b047c0490048a046c04490449047d04da045005ad05c6059c053e05cd048504;
    inBuf[4786] = 256'h7c04b3042705b4053906ad06fa0615070d07df0693064c061306f40506063b06;
    inBuf[4787] = 256'h7f06ce060e072c0737072d0714070d0710071407230728071a07170725075507;
    inBuf[4788] = 256'hbf074b08d1083d095d091e09aa081a08990761077007b5072b08a108fb084509;
    inBuf[4789] = 256'h7309840998099b097f0958091409ba08790858085e08a108fa0843097f099509;
    inBuf[4790] = 256'h8c099709b109d5090a0a260a160afe09e309dc090c0a540a900abe0aba0a880a;
    inBuf[4791] = 256'h5c0a3b0a280a380a440a380a320a2e0a3b0a850af10a600bca0bfb0bdd0b970b;
    inBuf[4792] = 256'h2e0bbf0a820a700a7d0ab50aeb0a090b240b250b120b1d0b3b0b6a0bc10b130c;
    inBuf[4793] = 256'h410c580c3f0c050ce70be60b010c450c750c670c2b0cb90b340bec0ae80a250b;
    inBuf[4794] = 256'ha60b240c720c990c860c4f0c320c2c0c350c5b0c6a0c500c350c140c010c290c;
    inBuf[4795] = 256'h660c960cb50c950c390ce10b990b7b0bb00b0d0c6d0cd00c030dfe0ce50cad0c;
    inBuf[4796] = 256'h620c340c110cf50bfb0bfe0bf10bf00be30bd00be40b0c0c400c940cda0cf80c;
    inBuf[4797] = 256'h010dd30c720c0e0ca30b460b260b2f0b550ba20be20bfe0b0f0c020ce20be00b;
    inBuf[4798] = 256'hea0bfa0b200c320c250c170cf50bc90bb80baa0b950b8e0b780b4d0b2e0b050b;
    inBuf[4799] = 256'hd40abc0aa30a880a8d0a9f0abe0a0a0b610bb50b0b0c320c170ccd0b440b940a;
    inBuf[4800] = 256'hfe09910965099609f409550aac0ac40a9b0a620a210af209f709100a280a470a;
    inBuf[4801] = 256'h4b0a340a220aff09c6098e094509fa08d808d508ee0824093f092509ee089c08;
    inBuf[4802] = 256'h560854088b08e7085409910983094009c7083c08d8079a078707a907d707fd07;
    inBuf[4803] = 256'h23082c081b080708e307b6079a078307750788079c07a107970760070107a206;
    inBuf[4804] = 256'h4e061f062e0658068606b506ce06d606e606ed06e106c4067d061f06db05c205;
    inBuf[4805] = 256'he3053d069106ab067906ed053605a2045a047204e3046a05cc05f105c7056d05;
    inBuf[4806] = 256'h1f05f304f1041705350530050b05c304710434040704eb03e103d603cc03d503;
    inBuf[4807] = 256'he503fd031c042c0429041b04ff03e303d203bc0399036f033403f402c902b402;
    inBuf[4808] = 256'hbc02d802e602d702ae026f023c02340257029702d802ed02c80276020d02b401;
    inBuf[4809] = 256'h84017501790179015e0132010c01fe0019015901a001d501e101b8016c011901;
    inBuf[4810] = 256'hd100a50094008c0086007e0072006d006e00650044000200a2ff43ff08ff0aff;
    inBuf[4811] = 256'h54ffcdff4900a300c100a2005a00feff9cff3dffddfe82fe3dfe1cfe2afe69fe;
    inBuf[4812] = 256'hc6fe21ff63ff73ff51ff0bffa8fe3bfed7fd86fd58fd61fda0fd0bfe87fee1fe;
    inBuf[4813] = 256'hf9fec3fe40fe97fdf8fc82fc49fc4efc77fcb1fcf1fc24fd4bfd6afd73fd66fd;
    inBuf[4814] = 256'h44fdfffca2fc3ffcddfb9afb8cfba7fbe1fb21fc3cfc2cfcfdfbbdfb94fb96fb;
    inBuf[4815] = 256'haefbc9fbcafb8ffb25fbb1fa4bfa1dfa38fa7dfad5fa20fb2efb00fbaafa39fa;
    inBuf[4816] = 256'he0f9c0f9ccf901fa46fa6cfa71fa5efa35fa12fafff9dff9aff96bf902f996f8;
    inBuf[4817] = 256'h49f825f843f89cf805f96df9bdf9ccf9a7f963f9fef89ef85bf82bf81ef836f8;
    inBuf[4818] = 256'h52f874f88ff87df847f8fcf79cf755f747f760f79ff7e9f708f800f8def7a8f7;
    inBuf[4819] = 256'h8cf79ff7bef7ddf7e2f7a3f73bf7cef66af642f666f6aaf6fff642f746f720f7;
    inBuf[4820] = 256'he6f69bf666f654f640f633f630f622f629f64cf66bf68ef6a4f687f64ef610f6;
    inBuf[4821] = 256'hc7f599f591f593f5acf5d7f5eff503f610f6f6f5ccf599f54cf509f5e1f4c3f4;
    inBuf[4822] = 256'hcdf404f542f58bf5c9f5caf5a3f55ff5faf4acf491f495f4c6f40ff53bf553f5;
    inBuf[4823] = 256'h54f528f5f8f4d9f4b9f4b8f4d1f4d6f4d0f4b7f474f438f425f437f48df40ff5;
    inBuf[4824] = 256'h76f5aff5a4f53cf5b3f43df4e5f3d7f307f43bf46ef494f494f49bf4bcf4dff4;
    inBuf[4825] = 256'h11f538f51ff5ddf48af42df408f431f481f4eff44ff564f541f5fbf495f44df4;
    inBuf[4826] = 256'h39f43af45df491f4adf4c7f4e3f4e9f4f9f414f51cf529f538f523f500f5d2f4;
    inBuf[4827] = 256'h89f453f447f459f4a2f412f56df5b3f5d1f5adf574f541f510f504f51cf530f5;
    inBuf[4828] = 256'h4cf565f560f55df567f567f578f594f595f58ff589f576f57df5a6f5d0f507f6;
    inBuf[4829] = 256'h3af641f638f62df615f615f62bf633f63bf63af61df60bf615f62ff674f6d9f6;
    inBuf[4830] = 256'h34f788f7bdf7aef771f717f7a4f654f641f665f6d0f666f7eaf74ff87bf855f8;
    inBuf[4831] = 256'h08f8b5f767f74ef773f7b7f71bf883f8c8f8f6f809f9f0f8caf8a0f86af84af8;
    inBuf[4832] = 256'h50f86ff8b7f811f953f97ff98af96cf953f957f977f9c3f921fa62fa81fa75fa;
    inBuf[4833] = 256'h39fafef9def9d9f902fa43fa72fa91fa97fa81fa73fa7ffa9dfad9fa1ffb51fb;
    inBuf[4834] = 256'h7afb99fba5fbbafbd7fbe8fbf3fbe9fbbffb91fb71fb6afb98fbf9fb6cfce1fc;
    inBuf[4835] = 256'h34fd47fd25fdd8fc75fc2afc11fc2ffc8dfc15fda2fd21fe6ffe74fe3efedbfd;
    inBuf[4836] = 256'h67fd10fdf0fc09fd5cfdcafd2dfe76fe99fe9efea9fec9fe03ff54ff9cffb7ff;
    inBuf[4837] = 256'h96ff3bffc1fe5afe2ffe58fedafe8fff4000c7000a010601d80097005b003000;
    inBuf[4838] = 256'h0f00f2ffdeffd9fff2ff350099000c017701bb01cf01b7017f0140011001ff00;
    inBuf[4839] = 256'h1c016701d0014302a602dd02e102b8027402360212020d022302410255026302;
    inBuf[4840] = 256'h76029d02e8025003b603fd030804ce036f031503ea020f037303eb0350047b04;
    inBuf[4841] = 256'h62042704ea03c603cf03f303190440045f047e04b7040705550592059f057305;
    inBuf[4842] = 256'h2f05f004d504f90442058405a80596055c0533053d0589050e068e06cb06b406;
    inBuf[4843] = 256'h4c06c10569056b05c905740620078d07a7076507e90678062e06180640068006;
    inBuf[4844] = 256'hb806ed0615073b078207d90727085f085908090899072307d106d5061e078c07;
    inBuf[4845] = 256'h09085b0864083c08ef07a3079207ba070e088408e1080009e9089a083208f007;
    inBuf[4846] = 256'hde07fc074b089808bf08c508a308700864087d08b10801093b09430931090a09;
    inBuf[4847] = 256'hea08fb0827095109730966092809ea08bb08ac08d7081509440966095d093209;
    inBuf[4848] = 256'h150906090d0945098c09c709fe09110afa09d6099f095c0935091a090e093209;
    inBuf[4849] = 256'h7309c209270a6d0a770a560a000a9109500946097609df09410a6a0a5e0a0a0a;
    inBuf[4850] = 256'h8e093709150933099a09080a4a0a560a140aa1094d0931095a09d4095c0ab80a;
    inBuf[4851] = 256'hdf0ab50a4e0ae909910952094109380928092a09340950099c09f909480a850a;
    inBuf[4852] = 256'h850a430ae9097f092109ff08060927096809a009bc09ce09be098d095e092609;
    inBuf[4853] = 256'hf108e108df08e308fe0812091e093e0966099109ce09f009df09a8093a09ac08;
    inBuf[4854] = 256'h3a08ef07da0712086f08d3083a097a098a0985095c091509d10884083c081e08;
    inBuf[4855] = 256'h1f083e088308c108db08d908a9085e0829080c080a082d084608430838081d08;
    inBuf[4856] = 256'h0608180842087308a308a60872082708c80770074e0754077507b107e007f407;
    inBuf[4857] = 256'hfe07f107d507c807b7079f078c076a073c071d070407f70609071d072a073407;
    inBuf[4858] = 256'h2307fa06d306a80688068f06ab06d006ff0616070e07f706cd06a00691068c06;
    inBuf[4859] = 256'h880682065a061106c605820561058005c205100657066d064d061006c1057e05;
    inBuf[4860] = 256'h68056d0581059f05a705970585056b05570554054c0536051805e704b504a204;
    inBuf[4861] = 256'ha904cb04050536054f05520533050405da04ad04820463043f041a040504fa03;
    inBuf[4862] = 256'h0304230442045a046e046e0462045a044b0436041b04eb03b0037f035f036303;
    inBuf[4863] = 256'h9203ce0304041d04fd03af034c03eb02ad02ab02d80226037703a2039b036603;
    inBuf[4864] = 256'h0e03b6027b0262026e029302b002b902ab0281024d021e02f401dc01d601d601;
    inBuf[4865] = 256'hdd01ea01f301fa01fe01f601e301c40193015d012b010001e800e400e800f500;
    inBuf[4866] = 256'h04010a010901fe00e900d200b9009900790056002a00feffdaffc3ffc4ffdaff;
    inBuf[4867] = 256'hf6ff11001600feffd6ffa8ff7bff5aff3dff1bfff7fed3febdfecafefafe3dff;
    inBuf[4868] = 256'h80ff9aff74ff13ff89fe01feaafd98fdc8fd25fe7cfea7fe9bfe5bfe05fec4fd;
    inBuf[4869] = 256'ha4fda8fdc5fdd5fdc2fd8dfd3cfdeafcb6fca3fcb3fcdffc06fd1cfd22fd11fd;
    inBuf[4870] = 256'hf3fcd6fcb1fc87fc5ffc30fc07fcf2fbecfbfafb1bfc34fc3bfc30fc01fcbafb;
    inBuf[4871] = 256'h6dfb1ffbe5facffad3faf2fa24fb44fb49fb34fbfcfab5fa77fa43fa2afa32fa;
    inBuf[4872] = 256'h43fa59fa70fa70fa5ffa44fa11fad6f99ff965f93bf92bf92af942f972f999f9;
    inBuf[4873] = 256'hb5f9bff99ff961f915f9bcf872f847f82ff833f855f876f898f8b9f8c0f8b4f8;
    inBuf[4874] = 256'h98f859f80cf8c6f77ff753f74bf750f768f78df7a6f7c2f7e7f7f7f7f9f7e7f7;
    inBuf[4875] = 256'ha7f74cf7edf68ef659f65df67df6b9f6fef622f72af71af7e4f6a8f679f64bf6;
    inBuf[4876] = 256'h34f634f629f621f61cf606f6fcf508f60df616f61ef606f6e0f5bcf58df573f5;
    inBuf[4877] = 256'h71f568f564f566f550f53ef53bf532f53cf559f568f574f577f550f51cf5e6f4;
    inBuf[4878] = 256'ha0f46ff460f455f462f481f490f4a4f4bcf4baf4b8f4b6f497f474f453f421f4;
    inBuf[4879] = 256'hfdf3f1f3e1f3e8f304f410f41cf428f419f40cf406f4eef3def3d8f3c1f3b9f3;
    inBuf[4880] = 256'hc5f3c9f3d9f3edf3e2f3cdf3b4f385f36af370f377f397f3c3f3cdf3c5f3a9f3;
    inBuf[4881] = 256'h66f327f304f3eef209f34bf384f3b8f3ddf3d0f3b2f392f35cf335f320f303f3;
    inBuf[4882] = 256'hfbf208f30ef327f351f368f386f3a7f3a7f3a1f397f36ff34af32df302f3eaf2;
    inBuf[4883] = 256'he5f2d8f2e2f207f32af360f39bf3b0f3b1f39ef363f32ef30ef3f0f2f6f21cf3;
    inBuf[4884] = 256'h3cf36af39cf3aef3b9f3bdf39ff382f36cf349f33af340f343f35ef38bf3a8f3;
    inBuf[4885] = 256'hcaf3ecf3f2f3fcf30cf409f40ff41af40ff40bf40ff402f403f40ef40af40ff4;
    inBuf[4886] = 256'h20f42af448f479f49ef4cff402f518f529f535f527f51cf516f504f506f51df5;
    inBuf[4887] = 256'h32f55cf591f5b3f5d7f5f8f5fff509f61af61ef62ef647f652f668f688f6a3f6;
    inBuf[4888] = 256'hd2f60df734f755f767f75cf752f755f75cf77ff7b2f7d6f7f7f712f81df837f8;
    inBuf[4889] = 256'h63f88ef8c3f8f5f809f910f914f912f927f952f97ff9b2f9dbf9e8f9f1f9fdf9;
    inBuf[4890] = 256'h0dfa39fa7bfabdfa01fb34fb43fb3efb2afb0cfb03fb15fb3bfb80fbd8fb2bfc;
    inBuf[4891] = 256'h77fcb1fcd0fce2fce6fcddfcdcfce3fcedfc0cfd3dfd7afdc6fd14fe57fe91fe;
    inBuf[4892] = 256'hb5febdfebbfeb2feabfeb6fed2fefbfe32ff6cffa7ffe7ff250060009a00c700;
    inBuf[4893] = 256'he300f200f300f100fc0014013f017901b301e70112022d024102580271029502;
    inBuf[4894] = 256'hc602f90232036e03a403d603fc030c0410040b040304110439047104bd040b05;
    inBuf[4895] = 256'h460572058a058d058f0594059c05ba05e605150653069506cc0602072a073c07;
    inBuf[4896] = 256'h4807450732072c07310740076f07b007f1073b0878089d08ba08c308b708b608;
    inBuf[4897] = 256'hb908c408f0082b0960099609b409b409bb09c309d309050a400a690a900a9f0a;
    inBuf[4898] = 256'h910a8f0a900a970abf0aef0a150b480b710b880bac0bc70bd20be60bee0be50b;
    inBuf[4899] = 256'hef0bff0b0e0c3c0c6b0c8c0cb60ccb0ccc0ce10cf70c050d2b0d4c0d5d0d7e0d;
    inBuf[4900] = 256'h920d900d9d0d9f0d930da50dc00ddd0d1c0e560e750e950e940e720e630e540e;
    inBuf[4901] = 256'h4a0e6f0e9b0ebc0ef00e110f160f2a0f360f330f490f540f4b0f570f5d0f5c0f;
    inBuf[4902] = 256'h800fa50fba0fe20ff20fe60fea0fe50fd70fed0ffd0ffd0f1810271024103d10;
    inBuf[4903] = 256'h501052106c107410661075107d107b109c10b610ba10ce10cb10b010b110ac10;
    inBuf[4904] = 256'h9d10b110c010be10d910ed10f61020113e11481163116311411131111211e910;
    inBuf[4905] = 256'hec10f81006113e116e118511a811a91187117611551127112311251127114f11;
    inBuf[4906] = 256'h6c11741193119c119011a011a311901192118011561149113a112e1153117a11;
    inBuf[4907] = 256'h9111b311ad117e115e1135110d111a11311141116911721158114d1130110411;
    inBuf[4908] = 256'hfb10ec10d110d310cb10ba10c810cb10be10ca10c0109d108b10671035102610;
    inBuf[4909] = 256'h1b1016103b10591061106d1050100a10ca0f800f3a0f2b0f2c0f360f630f800f;
    inBuf[4910] = 256'h7e0f7a0f540f140fe70eaf0e730e5d0e480e330e3f0e420e360e380e210ef60d;
    inBuf[4911] = 256'hdd0dba0d910d860d750d5a0d510d340d090df00ccd0c9f0c870c690c460c3c0c;
    inBuf[4912] = 256'h2d0c1d0c1f0c0e0ce80bc70b8f0b4a0b1d0bf30ad20acf0ac40aac0a9b0a760a;
    inBuf[4913] = 256'h480a300a180a040a010aea09ba0983093409de08a4087b086d0886089f08aa08;
    inBuf[4914] = 256'hac0886083f08f2079a0747071107e606cb06c806c606be06b606970667063306;
    inBuf[4915] = 256'hee05a6056e0538050f05f804e304d304c804ab047e044b040a04c80394036903;
    inBuf[4916] = 256'h4f0341032b030e03ed02bc02820249021102e201bf019c017e01640146012a01;
    inBuf[4917] = 256'h0d01e800bf008f0054001900dcffa0ff6dff3fff16fffdfef1feecfef1feedfe;
    inBuf[4918] = 256'hd2fe9ffe50fef1fd9cfd55fd26fd18fd17fd19fd1cfd0ffdf2fccefc9dfc66fc;
    inBuf[4919] = 256'h34fcf7fbb6fb7cfb44fb1ffb16fb15fb19fb1dfb03fbd2fa96fa49fa01fad4f9;
    inBuf[4920] = 256'hacf990f985f96ef953f93ef91af9f3f8d7f8b2f890f876f84df822f803f8d9f7;
    inBuf[4921] = 256'hbaf7aff79bf786f772f743f70bf7dbf69ef66ef659f643f63af642f630f614f6;
    inBuf[4922] = 256'hf3f5b4f576f54cf51cf5fff4fbf4eaf4dbf4d5f4b7f49af488f45ff436f415f4;
    inBuf[4923] = 256'hdbf3a6f387f361f34ff35af356f354f357f335f309f3e4f2a8f276f25ff23df2;
    inBuf[4924] = 256'h2bf22ff21ff215f214f2f3f1cff1b0f176f14af13ef129f129f141f13bf12df1;
    inBuf[4925] = 256'h1cf1dff0a1f077f03ef020f028f026f033f051f04ff04bf04af021f0f7efd5ef;
    inBuf[4926] = 256'h93ef60ef4cef2def29ef48ef50ef5cef6bef4def27ef08efceeea7ee9fee86ee;
    inBuf[4927] = 256'h81ee90ee80ee75ee7bee65ee5eee6dee5dee53ee4eee1deeeeedceed9bed8bed;
    inBuf[4928] = 256'ha7edb6edd6ed01eef6edd8edb7ed75ed50ed57ed5aed79eda9eda5ed90ed79ed;
    inBuf[4929] = 256'h3ced12ed0eed04ed16ed3ded3ced38ed3aed17ed06ed10ed04ed0aed1fed0aed;
    inBuf[4930] = 256'hfbecfeecebecf1ec13ed1bed2ced44ed30ed1fed19edf5ece7ecf4ece9ecf3ec;
    inBuf[4931] = 256'h12ed13ed23ed45ed49ed59ed73ed62ed51ed4bed28ed1aed29ed2ced4aed7ced;
    inBuf[4932] = 256'h8bed9eedb7edaaeda3edaaed97ed9aedb5edb7edcbedededebedf1ed06eeffed;
    inBuf[4933] = 256'h0aee29ee30ee46ee6cee70ee7cee93ee8cee91eea3ee9aeea3eec0eec6eedeee;
    inBuf[4934] = 256'h0bef21ef3fef62ef5def59ef5bef47ef51ef77ef8defb0efdeefecef03f024f0;
    inBuf[4935] = 256'h30f04ef079f085f096f0aaf09ff09ef0aff0b4f0d3f007f128f158f18df1a1f1;
    inBuf[4936] = 256'hb8f1d3f1d1f1dcf1f7f101f21bf246f261f288f2b6f2caf2e0f2faf201f31bf3;
    inBuf[4937] = 256'h46f361f38bf3bdf3d8f3f7f315f41cf432f453f465f489f4baf4d9f402f531f5;
    inBuf[4938] = 256'h4bf56df595f5adf5cff5f5f508f623f644f653f66ef695f6b2f6e0f618f743f7;
    inBuf[4939] = 256'h76f7a7f7c1f7d8f7ecf7f1f7fff718f82ef859f893f8caf809f946f96df98ff9;
    inBuf[4940] = 256'ha6f9a9f9b0f9bff9d0f9f8f92dfa5efa95fac9faebfa0dfb2efb4afb73fb9ffb;
    inBuf[4941] = 256'hc0fbe1fbf9fb00fc0cfc23fc43fc7afcbdfcfefc37fd5ffd70fd7bfd85fd98fd;
    inBuf[4942] = 256'hc2fdf7fd2cfe5efe7cfe85fe8bfe96feb5fef2fe44ff99ffe6ff140022001c00;
    inBuf[4943] = 256'h0b000200120038007000b000e8001a0149016f019901c601eb01090221022e02;
    inBuf[4944] = 256'h3a024d026a029a02d1020403380361037b039703b703d303f903210442046704;
    inBuf[4945] = 256'h85049804b604d804f904260556057c05a405c205d405ee050a0623064c067a06;
    inBuf[4946] = 256'ha206ce06ec06f60601070b0716073c077107ab07f3072b084308530852084408;
    inBuf[4947] = 256'h490858086e08a208dc080d094b097c099309aa09b509b009bb09c709d109f509;
    inBuf[4948] = 256'h180a320a5f0a850a9c0ac30ae40af90a1c0b360b3e0b530b610b630b790b8f0b;
    inBuf[4949] = 256'h9d0bbf0bda0bec0b140c380c520c7d0c980c990ca50ca50c9b0cb00ccd0ce70c;
    inBuf[4950] = 256'h1c0d440d530d6a0d6f0d630d770d910da70dd60dfa0d060e180e130efc0dfe0d;
    inBuf[4951] = 256'h020e050e2e0e590e770ea70ec40ec50ed10ecd0eba0ec40ecd0ece0eeb0eff0e;
    inBuf[4952] = 256'h030f1f0f330f390f590f6c0f6a0f790f780f670f700f740f6f0f8a0fa00fa30f;
    inBuf[4953] = 256'hbb0fc50fbf0fd30fdc0fd40fe90ff30fe70ff00ff00fdf0fe60fe50fda0fed0f;
    inBuf[4954] = 256'hf90ff80f1310231020102e102910111011100810f50f00100310f80f08100f10;
    inBuf[4955] = 256'h06101c102910231032102e1012100810f30fd60fda0fd90fce0fdf0fe30fd60f;
    inBuf[4956] = 256'he10fe50fdb0fea0feb0fd40fcd0fb20f850f750f670f580f6c0f7b0f7b0f8c0f;
    inBuf[4957] = 256'h880f6b0f5e0f440f240f240f1f0f0d0f130f090fea0edf0ecb0eae0eb00eac0e;
    inBuf[4958] = 256'h9c0ea10e960e770e6c0e570e380e380e310e190e140e030ee20dd70dc30da60d;
    inBuf[4959] = 256'ha00d910d730d690d550d360d300d240d0d0d080df30cce0cbc0ca30c820c7f0c;
    inBuf[4960] = 256'h780c660c650c540c2f0c150ced0bbc0ba60b900b740b700b660b550b560b490b;
    inBuf[4961] = 256'h2c0b1a0bf80ac80aac0a8d0a690a5d0a500a390a2d0a160af209dc09c0099f09;
    inBuf[4962] = 256'h9209800967095e09470923090809df08af0896087e0868086908640852084208;
    inBuf[4963] = 256'h2008ef07c907a007770765075107370728071407f706e606d006b506a5068b06;
    inBuf[4964] = 256'h640643061806eb05d005b8059f059205800565055105340515050105e804c804;
    inBuf[4965] = 256'haf048f0469044d04310417040604f103d603be039c0375035503350316030203;
    inBuf[4966] = 256'hed02d602c402ae0292027c02620245022c021202f301d601b801980179015a01;
    inBuf[4967] = 256'h410130011e010b01fa00e100c000a1008200680054004100310021000a00ecff;
    inBuf[4968] = 256'hcbffa8ff87ff6bff54ff44ff37ff2aff1aff05ffecfed1feb2fe92fe78fe64fe;
    inBuf[4969] = 256'h51fe3efe29fe14fefffde5fdcbfdb9fda8fd99fd8afd75fd5efd48fd2dfd14fd;
    inBuf[4970] = 256'h03fdf1fcdefccffcbbfca7fc93fc7cfc6afc5efc4cfc37fc25fc0dfcf2fbd9fb;
    inBuf[4971] = 256'hc0fbaffba8fb9efb96fb8efb7efb6cfb56fb37fb1efb11fb03fbfcfaf9faebfa;
    inBuf[4972] = 256'hdafac6faa6fa8afa7dfa71fa6efa74fa6ffa65fa56fa38fa1dfa0dfafef9faf9;
    inBuf[4973] = 256'h00fafaf9eff9e4f9cdf9b9f9aef99cf992f993f98af980f979f96af960f95cf9;
    inBuf[4974] = 256'h52f94cf94cf942f939f935f926f921f926f922f920f921f910f900f9f5f8e1f8;
    inBuf[4975] = 256'hd7f8dcf8def8e7f8f4f8edf8e3f8dbf8c6f8b8f8bbf8bdf8c6f8d3f8cef8c4f8;
    inBuf[4976] = 256'hbbf8a9f8a3f8acf8b0f8bbf8cbf8c8f8bff8b6f8a2f899f89bf897f8a0f8b5f8;
    inBuf[4977] = 256'hb8f8bbf8c2f8bef8bff8c6f8c0f8bbf8bbf8adf8a4f8a7f8a5f8b0f8c5f8ccf8;
    inBuf[4978] = 256'hd4f8ddf8d2f8c9f8c9f8c0f8bff8caf8cdf8d5f8e1f8ddf8dcf8e3f8e0f8e2f8;
    inBuf[4979] = 256'heef8f2f8faf804f9fff8fef802f9fbf8fef80bf90cf913f921f91ef91ff928f9;
    inBuf[4980] = 256'h26f92bf939f93af93df944f93cf93bf944f943f94bf95af95af95bf962f95ff9;
    inBuf[4981] = 256'h65f975f97cf989f99cf99bf995f990f97ff978f982f98af9a0f9bef9cbf9d5f9;
    inBuf[4982] = 256'hd9f9cbf9c1f9c2f9bef9c5f9d6f9dcf9e8f9f5f9f4f9f6f9fef9f9f9f9f9fef9;
    inBuf[4983] = 256'hf8f9f9f904fa06fa10fa24fa2efa37fa3ffa35fa2cfa2cfa28fa2ffa44fa53fa;
    inBuf[4984] = 256'h64fa73fa71fa6cfa66fa56fa4ffa51fa52fa60fa79fa84fa90fa9dfa9bfa96fa;
    inBuf[4985] = 256'h96fa8efa90fa9bfaa0faa8fab2faaefaaafaadfaa9faacfab9fac1facffadefa;
    inBuf[4986] = 256'hdefadffae4fadefadafae1fae4faebfafbfa05fb14fb23fb23fb20fb1dfb10fb;
    inBuf[4987] = 256'h08fb0dfb13fb22fb37fb44fb51fb59fb53fb4ffb50fb49fb4afb58fb63fb75fb;
    inBuf[4988] = 256'h8dfb9bfba5fba9fb9afb8afb82fb7cfb86fba0fbbafbd6fbeefbf1fbe6fbdbfb;
    inBuf[4989] = 256'hd0fbcffbdcfbecfb03fc18fc1dfc1dfc20fc1bfc1ffc2dfc39fc46fc55fc59fc;
    inBuf[4990] = 256'h5afc5afc55fc59fc66fc73fc83fc97fca1fca7fcaefcadfcaffcb7fcbcfcc2fc;
    inBuf[4991] = 256'hcafccefcd8fce8fcf0fcfbfc0efd1afd1ffd24fd23fd22fd25fd2dfd3cfd51fd;
    inBuf[4992] = 256'h5ffd6bfd72fd6bfd60fd5bfd5afd63fd79fd93fdaffdc7fdcffdd0fdcffdc7fd;
    inBuf[4993] = 256'hc2fdc7fdd0fdddfdedfdf8fd04fe13fe1bfe22fe29fe2afe29fe2cfe31fe3efe;
    inBuf[4994] = 256'h53fe65fe75fe83fe89fe87fe86fe86fe8bfe97fea6feb6fec5fecafecafecbfe;
    inBuf[4995] = 256'hccfed0fedafee9fef8fe06ff11ff18ff1eff21ff26ff30ff3bff49ff57ff60ff;
    inBuf[4996] = 256'h65ff6eff76ff7bff82ff87ff89ff8cff8fff95ffa5ffbaffccffdeffeaffeaff;
    inBuf[4997] = 256'he1ffd9ffd9ffe2fff4ff0d002a003e0045004100360029002200270036004e00;
    inBuf[4998] = 256'h66007a00890094009700960097009b00a300ab00b300bc00c500c900d000da00;
    inBuf[4999] = 256'he100e800f300fc0005010f01180122012d01330138014101460149014f015401;
    inBuf[5000] = 256'h590163016d017801830189018a018f0192019801a501b401c301d401e001e601;
    inBuf[5001] = 256'he801e501e301e701ef01fb010a02160222022d022c022702280229022d023c02;
    inBuf[5002] = 256'h4d02600276028202850285027f0277027b0283029002a202b002b802c002c002;
    inBuf[5003] = 256'hbc02c002c502cc02db02e902f40202030c030f03150319031c03220325032a03;
    inBuf[5004] = 256'h34033a0340034d03540356035c035e035e0366036e037703880393039a03a703;
    inBuf[5005] = 256'haa03a403a603a803aa03b603c303ce03de03e503e103df03d803d203dd03ed03;
    inBuf[5006] = 256'hff031a042c043004310427041704120413041d0430043c0441044b044c044704;
    inBuf[5007] = 256'h4d04540456045f04650467046f047304770486048d048e04950495048c048a04;
    inBuf[5008] = 256'h8604830490049c04a404b204b704b304b204ad04a704b104bd04c704d604dd04;
    inBuf[5009] = 256'hda04d604cc04c004c004c004c104cd04d204d104d904db04d804df04e204e004;
    inBuf[5010] = 256'he504e304db04de04df04dc04e204e404e404ea04e804e104e504e404df04e404;
    inBuf[5011] = 256'he504dd04da04d604d104d704d804d804e204e604de04dd04d704ca04c704c104;
    inBuf[5012] = 256'hb904bd04bf04bf04c804cb04c704c904c104af04a704a2049e04a904af04af04;
    inBuf[5013] = 256'hb304ab0497048c0483047a047f0483048204870485047a0476046f0464046204;
    inBuf[5014] = 256'h5f04570454044e0448044b0449044104400439042c04240417040a040b040b04;
    inBuf[5015] = 256'h08040e0412040d040704f903e903e403df03da03e003e103d903cf03bc03a303;
    inBuf[5016] = 256'h990391038c039603a103a103a003950380036e035f0356035d03640365036903;
    inBuf[5017] = 256'h630353034403320321031d031a0316031a0318030f030a030103f502f302ef02;
    inBuf[5018] = 256'he702e402dd02d002cc02c702c002c202c102b902b202a5029302870281028002;
    inBuf[5019] = 256'h8a029302950290027f026602530244023f024c025a02620266025d0247023202;
    inBuf[5020] = 256'h1f02130216021e022302290228021f0214020502f901f701f701f601f701f401;
    inBuf[5021] = 256'hed01ea01e201d501d001cd01c901cb01cb01c501c001b901b401b501b501b501;
    inBuf[5022] = 256'hb801b601ae01a7019f0198019601940195019901950188017a016d0165016701;
    inBuf[5023] = 256'h6f017d0191019b019501860171015a014c0147014b015b016c01760175016a01;
    inBuf[5024] = 256'h570146013a0135013c01490155015b0157014d01410135013101380143014a01;
    inBuf[5025] = 256'h4d014a013d012b011e0118011c0124012d0133013101290122011d011c012101;
    inBuf[5026] = 256'h2601280126011c010e0104010101010106010f011801190111010601fc00f400;
    inBuf[5027] = 256'hf400fb000601100111010701f800e500d300cc00d200de00ec00f600f700ec00;
    inBuf[5028] = 256'hd900c600bc00ba00bd00c900d600dc00da00d200c500b800b000af00af00af00;
    inBuf[5029] = 256'hb100b100ab00a00095008c0088008b0091009600950091008c00860080007e00;
    inBuf[5030] = 256'h7e007c00790076006d00620059005300500054005a005b0057004e0041003500;
    inBuf[5031] = 256'h2c0028002f003a004000400037002a001e0012000b000c000e00120015000e00;
    inBuf[5032] = 256'h0100f4ffe8ffdfffdeffe2ffe9ffeffff1ffedffe5ffd8ffc8ffbaffb0ffacff;
    inBuf[5033] = 256'hb0ffb4ffb5ffb4ffacffa2ff9aff95ff94ff98ff99ff96ff8fff86ff7aff6fff;
    inBuf[5034] = 256'h69ff67ff67ff65ff61ff59ff4dff45ff41ff3fff42ff47ff49ff45ff3cff2fff;
    inBuf[5035] = 256'h22ff19ff0fff0dff12ff13ff11ff11ff0afffdfeeffee3fedcfedcfedefee2fe;
    inBuf[5036] = 256'he4fedffed4fec7febafeb4feb6febcfec4fecafec6febcfeacfe97fe86fe7ffe;
    inBuf[5037] = 256'h7bfe7dfe85fe88fe87fe82fe77fe6efe67fe60fe5dfe5dfe57fe53fe52fe4bfe;
    inBuf[5038] = 256'h45fe41fe3bfe37fe35fe2ffe29fe26fe1ffe18fe14fe0ffe09fe09fe06fefffd;
    inBuf[5039] = 256'hf8fdeffdeafde8fde5fde5fde8fde5fdddfdd4fdc4fdb4fdabfda5fda6fdadfd;
    inBuf[5040] = 256'hb0fdb0fdaffda6fd98fd8dfd83fd7bfd7afd7afd7bfd7afd70fd63fd57fd48fd;
    inBuf[5041] = 256'h40fd40fd41fd47fd50fd4ffd47fd3efd2cfd1cfd14fd0dfd0dfd14fd14fd0ffd;
    inBuf[5042] = 256'h0afdfdfcf0fce8fce0fcdcfcdcfcd7fcd2fccefcc3fcbefcbffcbcfcbbfcbdfc;
    inBuf[5043] = 256'hb4fcabfca2fc92fc89fc8bfc8afc8cfc93fc8dfc7ffc72fc60fc50fc4efc4ffc;
    inBuf[5044] = 256'h54fc5cfc5dfc59fc53fc44fc37fc30fc27fc24fc27fc23fc20fc1efc12fc06fc;
    inBuf[5045] = 256'h00fcf7fbf5fbfafbf6fbf4fbf6fbedfbe1fbd7fbc9fbc3fbc5fbc0fbc1fbc7fb;
    inBuf[5046] = 256'hc3fbbefbbdfbaffba2fb9cfb93fb8dfb8cfb86fb86fb89fb82fb7efb7ffb77fb;
    inBuf[5047] = 256'h70fb6dfb60fb54fb4ffb46fb46fb4cfb49fb49fb4afb3cfb30fb2bfb1ffb17fb;
    inBuf[5048] = 256'h1cfb1cfb23fb2efb2afb21fb16fbfffaeefaebfae8faebfaf6faf8faf8faf6fa;
    inBuf[5049] = 256'he6fad9fad4faccfacdfad8fad8fad4fad2fac7fabefabdfab4fab5fac0fabefa;
    inBuf[5050] = 256'hbafabafaaffaa5faa2fa9afa99fa9ffa9efaa1faa8faa3faa1faa3fa9bfa98fa;
    inBuf[5051] = 256'h9efa98fa93fa95fa8efa8bfa90fa8efa8ffa96fa95fa93fa93fa88fa82fa86fa;
    inBuf[5052] = 256'h86fa8dfa9afa9efaa1faa2fa95fa8bfa8afa83fa85fa93fa9afaa2faadfaadfa;
    inBuf[5053] = 256'haafaa9faa2faa2faabfaacfab0fabafab9fabafac0fabefac2facdfacefad1fa;
    inBuf[5054] = 256'hd8fad5fad3fad8fad7fadefaedfaf0faf6fa00fbfffafffa06fb08fb11fb1efb;
    inBuf[5055] = 256'h20fb23fb29fb27fb29fb32fb35fb3efb4bfb4ffb56fb5ffb5efb63fb70fb73fb;
    inBuf[5056] = 256'h7bfb8bfb91fb98fba1fba3fba7fbaefbabfbacfbb6fbc0fbcffbe0fbe8fbf2fb;
    inBuf[5057] = 256'hfdfbfbfbfafbfdfbfffb09fc19fc26fc35fc46fc4bfc4efc56fc58fc5dfc66fc;
    inBuf[5058] = 256'h6cfc75fc80fc84fc8dfc9bfca5fcb3fcc4fccafccefcd6fcdafce1fcebfceefc;
    inBuf[5059] = 256'hf8fc07fd0dfd12fd1bfd20fd27fd37fd45fd53fd62fd6afd71fd77fd79fd80fd;
    inBuf[5060] = 256'h8bfd92fd9cfda9fdb2fdbafdc4fdcafdd4fddffde5fdeffdfcfd04fe0cfe18fe;
    inBuf[5061] = 256'h22fe2dfe3afe42fe49fe50fe54fe59fe63fe6dfe79fe89fe94fe9afe9dfe9ffe;
    inBuf[5062] = 256'ha5feb0febbfec7fed6fee4fef1fefcfefffe00ff06ff10ff1cff29ff32ff39ff;
    inBuf[5063] = 256'h40ff46ff4cff53ff5eff69ff71ff78ff80ff89ff90ff9affa7ffb2ffbaffc2ff;
    inBuf[5064] = 256'hc6ffc9ffceffd5ffddffe7fff4ff000008000e00120016001d0025002c003800;
    inBuf[5065] = 256'h4600500058005e00610066006a006c00760084008f009a00a300a500a400a500;
    inBuf[5066] = 256'ha900b100bb00c600d500e200eb00f200f400f200f400fa00ff0006010e011301;
    inBuf[5067] = 256'h1a0121012c013b01450148014c01510153015801610169017101780182018a01;
    inBuf[5068] = 256'h8b018c01910193019601a101ac01b501c201ca01ca01ca01cb01cd01d501df01;
    inBuf[5069] = 256'he801f601010204020802080204020802100219022602320236023a023a023902;
    inBuf[5070] = 256'h3d0242024902580265026d02760279027502770278027802800287028b029502;
    inBuf[5071] = 256'h9e02a002a602ab02ac02b102ba02c002c502c702ca02cf02d102d602e202eb02;
    inBuf[5072] = 256'hed02ef02ee02ec02ed02ee02f40202030c0313031b031a031203110311031303;
    inBuf[5073] = 256'h1d032a033403400341033803350332032c0330033b0344034f03550352035003;
    inBuf[5074] = 256'h4b034903500359035e0369036d036903680364035e0364036b036d0372037203;
    inBuf[5075] = 256'h6d036d036e036f0377037c037d0383038203790377037603730377037e038003;
    inBuf[5076] = 256'h8603860381037f037b03750377037b03800388038a0383037f03790370036f03;
    inBuf[5077] = 256'h720374037e0386038403800379036c036503640365036c037303750376037103;
    inBuf[5078] = 256'h65035e035c035d0364036703640362035d0352034a034603440347034b034d03;
    inBuf[5079] = 256'h52035003470341033b033503350335033403360333032b032603220320032603;
    inBuf[5080] = 256'h2703240323031a030d030403fc02f902010308030d0313030e030203fb02f202;
    inBuf[5081] = 256'he902eb02f002f202f502f302eb02e302d802cf02d002d102d202d902dd02d702;
    inBuf[5082] = 256'hd102cc02c402c302c402c302c602c702c202be02b602ad02ab02ab02ac02b202;
    inBuf[5083] = 256'hb702b602b402ab029e029a02990299029c029e029d029e029902930290028d02;
    inBuf[5084] = 256'h8e02940292028d028e028b0282027d027b027b0283028702860285027f027502;
    inBuf[5085] = 256'h6f026b026c027202750277027b0276026d02690263025f02640269026d027202;
    inBuf[5086] = 256'h6f026602600257024e025002530254025a025d025902570253024d024c024d02;
    inBuf[5087] = 256'h4c024b024a02480245023e0239023c023f0240024302450240023b0232022c02;
    inBuf[5088] = 256'h2c022b0229022c022d02290224021e02170217021c0222022602260224022002;
    inBuf[5089] = 256'h130205020002fe01000209020f020f020a02ff01f601f001e901ea01f401fa01;
    inBuf[5090] = 256'hfb01f601ed01e201d601cc01cc01d301d801dc01de01d801cd01c301b901b501;
    inBuf[5091] = 256'hb601b501b401b401ad01a301a0019d0199019b019d019d019b01920186017c01;
    inBuf[5092] = 256'h7401700170017101740175016d0163015c0152014c014d014c014a0148014001;
    inBuf[5093] = 256'h3601310128011f011b011a011a011c011b0115010d010101f600ee00e700e500;
    inBuf[5094] = 256'he600e500e000d900d100ca00c400bd00ba00ba00b600af00a7009c0092008700;
    inBuf[5095] = 256'h7e007d007e007d007c0078006f00630057004f004b004800450043003b002f00;
    inBuf[5096] = 256'h2300180010000f00110010000e000a000000f4ffe8ffdeffdaffdaffd6ffd3ff;
    inBuf[5097] = 256'hceffc3ffb6ffacffa5ffa2ffa2ffa1ff9fff9dff94ff88ff7dff72ff68ff61ff;
    inBuf[5098] = 256'h61ff61ff5eff5bff57ff4eff43ff3bff33ff2dff2cff2aff25ff21ff19ff0dff;
    inBuf[5099] = 256'h03fffefefffe00fffefefffefcfeeffee1fed7fecdfec9fec9fec7fec6fec4fe;
    inBuf[5100] = 256'hbcfeb5feb1fea9fea7feaafea7fea4fea3fe99fe8dfe87fe7ffe77fe76fe77fe;
    inBuf[5101] = 256'h77fe78fe75fe6efe69fe62fe5bfe59fe59fe58fe56fe50fe48fe40fe37fe32fe;
    inBuf[5102] = 256'h34fe37fe3afe3ffe3efe35fe2cfe22fe18fe14fe11fe11fe15fe16fe13fe0ffe;
    inBuf[5103] = 256'h08fe02fe01fe00fe02fe07fe07fe01fefafdf2fdeafde4fddffde3fdeafdecfd;
    inBuf[5104] = 256'hebfdeafde5fde0fdd9fdd2fdd3fdd8fdd6fdd5fdd6fdcefdc5fdc2fdc1fdc3fd;
    inBuf[5105] = 256'hc9fdcdfdcffdcefdc8fdc1fdbbfdb6fdb7fdbafdb9fdbcfdbefdb9fdb6fdb7fd;
    inBuf[5106] = 256'hb6fdb7fdbbfdbdfdbefdbefdb6fdaffdabfda7fda8fdb0fdb5fdb8fdbdfdbefd;
    inBuf[5107] = 256'hbdfdbbfdb8fdb6fdb7fdb7fdbafdbcfdb7fdb3fdb5fdb4fdb4fdb8fdbdfdc6fd;
    inBuf[5108] = 256'hcffdd0fdd0fdd0fdc9fdc4fdc7fdc8fdccfdd5fddbfddefde0fdddfddcfddcfd;
    inBuf[5109] = 256'hddfde6fdedfdeffdf4fdf8fdf4fdf2fdf3fdf3fdf8fd03fe0cfe14fe18fe16fe;
    inBuf[5110] = 256'h17fe1afe1bfe1ffe25fe29fe2ffe31fe2ffe32fe36fe3afe42fe4dfe56fe60fe;
    inBuf[5111] = 256'h65fe63fe63fe65fe63fe66fe70fe7afe84fe8efe91fe91fe94fe96fe9bfea6fe;
    inBuf[5112] = 256'haefeb5febdfebefebcfebffec2fec7fed1fedefeebfef5fef9fefdfe02ff02ff;
    inBuf[5113] = 256'h03ff0aff12ff1bff26ff2dff2fff33ff37ff3cff44ff51ff5eff6bff74ff7bff;
    inBuf[5114] = 256'h7dff7dff7dff80ff85ff8eff9affa7ffaeffb2ffb8ffc1ffc8ffd2ffe0ffeaff;
    inBuf[5115] = 256'hf2fff8fff9fff9fff9fffdff0600130020002e0039003f004200450049004d00;
    inBuf[5116] = 256'h560062006c00730078007c00800086008f009a00a800b300bb00c000c000bf00;
    inBuf[5117] = 256'hc200c700cf00d900e200ec00f600fc00000106010d0114011e012a0131013301;
    inBuf[5118] = 256'h360138013801390140014a0155015e016701700173017401760178017b018301;
    inBuf[5119] = 256'h8e019401970198019a019e01a201a801b501c001c501c701c701c701c701c701;
    inBuf[5120] = 256'hc801cf01d901e001e601e901eb01ed01f101f701fc01fd01000203020102fe01;
    inBuf[5121] = 256'hfd01fc01fc0102020b0214021b021d021e021f021e021b021b021d021f022102;
    inBuf[5122] = 256'h23022302240221021e021d022102290231023302320231022c02270226022802;
    inBuf[5123] = 256'h2b022f0230022f022e022b0227022802290228022902260222021e0219021702;
    inBuf[5124] = 256'h1802180217021d0220021e021d021b02160212020d020b02090204020002ff01;
    inBuf[5125] = 256'hfa01f501f401f501f701f801f401f201f001e801df01dc01d801d401d401d201;
    inBuf[5126] = 256'hce01cd01c901bf01b901b601b301b101af01ab01a601a1019a0193018c018501;
    inBuf[5127] = 256'h820180017f017f017e017b017301690160015a0153014c014b0147013f013801;
    inBuf[5128] = 256'h34012f012d012f012e01290122011a0110010701ff00f700ee00e900e600e200;
    inBuf[5129] = 256'he100df00da00d500d200ce00c900c300ba00b300ad00a5009f009a0093008c00;
    inBuf[5130] = 256'h8a00880084007e0075006d00650060005d005b00590057005100490041003b00;
    inBuf[5131] = 256'h3800360033002d00270021001a0013000c000500fffffafff8fff6fff2fff1ff;
    inBuf[5132] = 256'hefffebffe9ffe7ffe1ffd8ffd0ffc9ffc5ffc0ffbaffb7ffb4ffafffadffabff;
    inBuf[5133] = 256'ha6ffa1ffa0ff9bff96ff93ff8fff89ff86ff82ff7cff77ff76ff74ff71ff6dff;
    inBuf[5134] = 256'h6aff67ff63ff5cff58ff54ff51ff4eff4aff44ff40ff3cff3aff3bff3bff3aff;
    inBuf[5135] = 256'h38ff31ff27ff23ff21ff1fff1cff1aff19ff16ff0fff0bff0aff08ff09ff0bff;
    inBuf[5136] = 256'h0cff0aff06ff00fffcfef7feeffeebfeecfeeefeeffeeffeecfee9fee7fee5fe;
    inBuf[5137] = 256'he5fee2fedefedffee0fedffedcfed8fed4fed3fed5fed6fed7fed7fed5fed4fe;
    inBuf[5138] = 256'hd2fecdfecafecbfeccfecbfecbfec8fec7fec9fecafec9fecbfecefecffecffe;
    inBuf[5139] = 256'hcefecefecbfec5fec6fec8fec5fec6fecbfecbfecafecbfecafecafec9fec8fe;
    inBuf[5140] = 256'hcffed6fed5fed4fed4fecffeccfec9fec8fecdfed4fed6fed8fedafed7fed5fe;
    inBuf[5141] = 256'hd3fed1fed2fed5fed7fed9fedcfedbfedbfedafed5fed6feddfee1fee2fee2fe;
    inBuf[5142] = 256'hdffedcfedbfed7fed6fedbfee1fee7feeafee6fee2fee3fee3fee3fee4fee6fe;
    inBuf[5143] = 256'heafeebfee5fee2fee2fedffeddfee1fee5fee7fee9fee9fee9fee6fee2fee2fe;
    inBuf[5144] = 256'he4fee3fee6feebfeeafee9fee8fee2fee0fee3fee5fee7fee9feeafee9fee4fe;
    inBuf[5145] = 256'hdffedefedffedefee3fee9feeafee9fee7fee3fee1fee3fee3fee3fee2fee4fe;
    inBuf[5146] = 256'he5fee3fedffedefedffedffee0fee3fee4fee3fee3fee3fee3fee1fedffee3fe;
    inBuf[5147] = 256'he7fee8fee9fee9fee5fee1fedffee0fee4fee8feebfeeefeedfee9fee9feecfe;
    inBuf[5148] = 256'hebfeeafeecfeeefef0feeffeeffef1feeffeebfeedfef0fef0fef5fefafef9fe;
    inBuf[5149] = 256'hf9fef8fef5fef3fef5fef9fe00ff06ff06ff06ff05ff00fffbfefbfefffe05ff;
    inBuf[5150] = 256'h08ff09ff09ff08ff06ff06ff06ff09ff10ff15ff13ff12ff14ff14ff13ff13ff;
    inBuf[5151] = 256'h13ff14ff17ff18ff18ff18ff15ff15ff14ff13ff17ff1fff22ff23ff23ff20ff;
    inBuf[5152] = 256'h1dff1dff1dff1fff22ff27ff2cff2bff25ff22ff20ff1fff22ff28ff2bff2dff;
    inBuf[5153] = 256'h2fff2bff29ff2aff2aff2aff2fff31ff33ff37ff37ff34ff34ff35ff34ff35ff;
    inBuf[5154] = 256'h36ff37ff3aff3dff3bff39ff39ff3aff3cff41ff46ff48ff4aff4bff46ff41ff;
    inBuf[5155] = 256'h42ff45ff48ff4dff53ff53ff51ff51ff52ff53ff55ff58ff5bff5fff64ff64ff;
    inBuf[5156] = 256'h63ff66ff68ff66ff67ff6cff6fff70ff73ff74ff72ff73ff76ff77ff79ff7eff;
    inBuf[5157] = 256'h83ff8aff8eff8cff8bff8cff8cff90ff98ff9cff9effa0ffa2ff9fff9cff9eff;
    inBuf[5158] = 256'ha3ffa8ffacffb1ffb3ffb4ffb6ffb8ffbcffc2ffc7ffc9ffcdffcfffcfffcfff;
    inBuf[5159] = 256'hd1ffd3ffd8ffdcffe0ffe4ffe7ffeaffebffebffedfff0fff2fff8ff01000600;
    inBuf[5160] = 256'h09000a0009000a000d00130018001d002200270028002600280028002a003000;
    inBuf[5161] = 256'h38003e004300470049004b004d005000550059005e006400670068006a006e00;
    inBuf[5162] = 256'h7100730076007b00830089008e009300970098009b009d009e00a300aa00ae00;
    inBuf[5163] = 256'hb000b200b400b800be00c100c700ce00d100d500da00dc00dd00e100e900f100;
    inBuf[5164] = 256'hf500f900fe0000010201060109010c011201160119011e012101240129012d01;
    inBuf[5165] = 256'h32013b01430149014e0150015101540152015201560159015f0168016d017201;
    inBuf[5166] = 256'h7801780176017c0185018b018f0192019501980199019b01a001a401a701ad01;
    inBuf[5167] = 256'hb201b401b801bb01bc01c101c601c801cc01d001d201d601d801d901de01e201;
    inBuf[5168] = 256'he401eb01ef01ef01f201f301f201f501f801f901fd01020206020a020a020a02;
    inBuf[5169] = 256'h0e021002120219021c021b021d021d021d021f021f021d022002230227022b02;
    inBuf[5170] = 256'h2b022c02300231022e022e023002330236023802380238023702340235023702;
    inBuf[5171] = 256'h3b023e023e023c023d023b0237023602370238023d0240023d023d023e023d02;
    inBuf[5172] = 256'h3c023a0238023b023b023502320230022d022c022b022b023002310232023202;
    inBuf[5173] = 256'h2d02270226022402220224022302220223021f021602120210020f020f020e02;
    inBuf[5174] = 256'h0d020d0208020202ff01fd01fb01fb01f901f701f601f201ed01e801e301df01;
    inBuf[5175] = 256'hde01db01d801d701d201ce01cd01c801c301c101bf01bd01be01bb01b501b101;
    inBuf[5176] = 256'hab01a501a1019a019601970193018c01880181017a017a017b017a017a017501;
    inBuf[5177] = 256'h70016c0160015601550152014b014901450140013c0133012d012c0127012401;
    inBuf[5178] = 256'h25012101190115010e0106010201fe00fc00fa00f500ee00e900e200da00d300;
    inBuf[5179] = 256'hce00ca00c600c100bc00b800b100a800a2009f009f009d009a0095008d008500;
    inBuf[5180] = 256'h80007a00740070006b0064005e0056004c00460043003e003b00390035003000;
    inBuf[5181] = 256'h2a0023001e0017000f000d000b0007000300fbfff2ffecffe5ffdcffd6ffd1ff;
    inBuf[5182] = 256'hceffcdffc9ffc2ffbeffb9ffafffaaffa8ffa2ff9dff9aff94ff8eff88ff80ff;
    inBuf[5183] = 256'h7aff75ff70ff6bff66ff5fff5aff56ff51ff4fff4cff47ff42ff39ff32ff2fff;
    inBuf[5184] = 256'h29ff21ff1cff18ff13ff12ff0fff0aff04fffefefafef7fef0feeafee8fee3fe;
    inBuf[5185] = 256'hddfed7fed2fecffec9fec1febefebdfeb7feb3feb1feacfea7fea2fe9bfe96fe;
    inBuf[5186] = 256'h96fe93fe8efe8bfe86fe81fe7efe78fe74fe73fe6ffe69fe68fe63fe5dfe5afe;
    inBuf[5187] = 256'h57fe50fe4bfe49fe48fe46fe43fe42fe43fe3efe38fe35fe31fe2dfe2bfe26fe;
    inBuf[5188] = 256'h23fe23fe1ffe1bfe1bfe16fe12fe12fe0efe0bfe0cfe07fe04fe05fe06fe07fe;
    inBuf[5189] = 256'h05fe00fefdfdfbfdf5fdf4fdf4fdf1fdf0fdeffdeafde9fde9fde4fde4fde6fd;
    inBuf[5190] = 256'he1fddffde4fde3fde0fde1fde2fde2fde3fde1fddefddefdddfdddfdddfddafd;
    inBuf[5191] = 256'hd8fdd7fdd6fdd6fdd6fdd6fdd9fddcfddafddafddefddafdd7fddbfddbfdd9fd;
    inBuf[5192] = 256'hdafdd9fddafddefddefddcfddefdddfdddfde1fde0fde1fde6fde5fde6fdeafd;
    inBuf[5193] = 256'he8fde9fdeefdeefdf1fdf6fdf3fdf3fdf9fdf8fdf8fdfdfdfcfdfcfd01fe01fe;
    inBuf[5194] = 256'h04fe0afe0bfe0dfe12fe14fe17fe1afe18fe19fe1cfe1efe22fe26fe25fe26fe;
    inBuf[5195] = 256'h2bfe2ffe35fe3cfe3ffe41fe46fe48fe4afe50fe54fe59fe5efe5ffe64fe69fe;
    inBuf[5196] = 256'h68fe68fe6cfe6ffe76fe7ffe80fe84fe89fe89fe8efe99fe9cfea1fea9fea9fe;
    inBuf[5197] = 256'haefeb9febafebbfec2fec6fecbfed3fed5fedbfee1fee0fee4feeffef1fef4fe;
    inBuf[5198] = 256'hfefe04ff09ff11ff16ff1bff21ff24ff2bff31ff35ff39ff3eff40ff42ff49ff;
    inBuf[5199] = 256'h50ff56ff5cff62ff69ff6eff73ff7aff7fff84ff8bff91ff95ff98ff9dffa3ff;
    inBuf[5200] = 256'ha8ffaeffb3ffb9ffbcffc1ffc8ffceffd0ffd4ffd8ffdbffe1ffe7ffecfff4ff;
    inBuf[5201] = 256'hfbfffdff030009000b000f0016001a001e002300230025002b00300035003a00;
    inBuf[5202] = 256'h3d0043004b005000530057005b0060006300620065006b006e00700076007c00;
    inBuf[5203] = 256'h7f00800085008a008f00930097009a009b009c009f00a300a700a900ad00b200;
    inBuf[5204] = 256'hb600b900bc00bf00c100c500c900cb00cc00cf00d200d500da00de00e000e300;
    inBuf[5205] = 256'he600e800ec00ef00f000f100f300f300f400f700fb00ff00010105010a010c01;
    inBuf[5206] = 256'h0b010d0110011101140118011a011c0120012201230125012401250129012901;
    inBuf[5207] = 256'h29012d012f012e01310135013601360139013b013c013d013f01410143014501;
    inBuf[5208] = 256'h48014601450148014a0148014801480149014c014f014f01500151014f015101;
    inBuf[5209] = 256'h5201510154015601550155015601540152015201530155015601560155015101;
    inBuf[5210] = 256'h4f01500150014f01500151015101530151014c014a014b014a01490147014601;
    inBuf[5211] = 256'h4701470144014301430141013e013c013b013a0138013401310130012e012d01;
    inBuf[5212] = 256'h2c01290128012801240120011e011c011b011b01190117011501110110010e01;
    inBuf[5213] = 256'h0a0109010901050102010001fc00fb00fa00f600f600f400ef00ed00eb00e700;
    inBuf[5214] = 256'he600e300df00de00da00d500d500d500d200d100ce00cb00ca00c700c500c300;
    inBuf[5215] = 256'hbf00bc00bc00b700b200b100b100af00b000af00ac00aa00a600a2009e009a00;
    inBuf[5216] = 256'h99009a009a009700960093008e008d008c008700850082007f00800080007a00;
    inBuf[5217] = 256'h780077007400740074006f006e006d006900660062005c005d005e005a005800;
    inBuf[5218] = 256'h5700550053004d004a004b004a004700460043003f003d003900360035003300;
    inBuf[5219] = 256'h320030002e002d002c002a002b0029002400210021001e001b00160013001500;
    inBuf[5220] = 256'h14001000100010000d000c000a000700030002000100ffffffff00000000fdff;
    inBuf[5221] = 256'hfbfff8fff6fff6fff7fff7fff5fff4fff5fff1ffebffebffecffe9ffe6ffe6ff;
    inBuf[5222] = 256'he9ffecffebffebffedffecffe8ffe7ffe9ffe9ffe8ffe8ffe7ffe4ffe1ffe1ff;
    inBuf[5223] = 256'he0ffe0ffe4ffe5ffe4ffe6ffe5ffe0ffe2ffe6ffe6ffe9ffebffecffedffebff;
    inBuf[5224] = 256'he6ffe6ffebffebffe8ffe9ffedffefffeeffefffefffeefff1fff3fff3fff4ff;
    inBuf[5225] = 256'hf4fff3fff5fff8fffafff8fff7fff8fffafffcfffefffffffdfffeff00000200;
    inBuf[5226] = 256'h04000600060005000500060009000c000c000a000e0013001300110012001200;
    inBuf[5227] = 256'h0f0011001300120015001900190019001b001d001f0020001f00200022002400;
    inBuf[5228] = 256'h230023002300240023002400280029002a002e0030002c002b002c002c002e00;
    inBuf[5229] = 256'h3200330034003600340033003300320033003800390037003700380037003600;
    inBuf[5230] = 256'h370039003b003c003e003e003c003d003e003d003f0042004100400040003f00;
    inBuf[5231] = 256'h400041003f0040004400460047004700470049004a0048004600460046004900;
    inBuf[5232] = 256'h4900450044004500430044004a004d004c004c004b004b004d004e004c004c00;
    inBuf[5233] = 256'h4c004c004c004d004e004d004a004b004c004c004d004a0048004a004c004b00;
    inBuf[5234] = 256'h4c004c0049004a004b004b004b004a0048004600440044004600460047004900;
    inBuf[5235] = 256'h480047004600440042004100410041004100400040004100420041003e003c00;
    inBuf[5236] = 256'h3c003c003b003a00380038003800370036003700360033003200340032002d00;
    inBuf[5237] = 256'h2d0030002e002b002b0029002800290029002900280025002300250025002100;
    inBuf[5238] = 256'h1f00200020002000210020001a00170017001500140014001200110012001400;
    inBuf[5239] = 256'h150012000f000f000e000f000f000c000b000c000800060005000000fdfffeff;
    inBuf[5240] = 256'hfafff8fffbfffafff7fff7fff7fff8fff6fff2fff3fff5fff2ffefffeeffedff;
    inBuf[5241] = 256'hecffe9ffe4ffe3ffe3ffe1ffdeffdbffd8ffd7ffd6ffd5ffd2ffceffd0ffd2ff;
    inBuf[5242] = 256'hd2ffcfffccffcaffc8ffc6ffc3ffc2ffc0ffbbffb6ffb6ffb5ffb0ffadffaeff;
    inBuf[5243] = 256'hadffaaffa9ffa6ffa4ffa5ffa4ffa1ffa1ffa1ff9fff9eff99ff93ff91ff90ff;
    inBuf[5244] = 256'h91ff92ff90ff8cff8aff88ff86ff83ff81ff80ff7fff7dff7cff7cff7bff7aff;
    inBuf[5245] = 256'h79ff7aff7aff76ff74ff74ff71ff6fff6fff6bff69ff6bff6aff69ff6aff68ff;
    inBuf[5246] = 256'h66ff65ff63ff64ff67ff69ff68ff65ff65ff65ff63ff5fff5dff5cff5cff5cff;
    inBuf[5247] = 256'h5aff5aff5cff5dff5cff5bff5cff5dff5fff61ff61ff5fff5eff5fff5eff5eff;
    inBuf[5248] = 256'h60ff5eff58ff58ff5cff5eff5eff5cff5aff5cff5eff5dff5dff5fff5fff5fff;
    inBuf[5249] = 256'h61ff61ff60ff61ff61ff5fff5eff5dff5cff5dff5eff5fff61ff61ff60ff60ff;
    inBuf[5250] = 256'h60ff62ff65ff63ff60ff62ff64ff65ff65ff66ff65ff63ff62ff65ff67ff65ff;
    inBuf[5251] = 256'h65ff68ff6cff6eff6eff6dff6eff6dff6cff70ff71ff6fff70ff74ff74ff76ff;
    inBuf[5252] = 256'h76ff74ff76ff7cff7dff7bff7cff7eff80ff82ff83ff86ff8aff8aff8aff8eff;
    inBuf[5253] = 256'h91ff8fff8fff93ff94ff93ff94ff95ff98ff9cffa0ffa4ffa7ffa8ffaaffadff;
    inBuf[5254] = 256'hafffafffb1ffb5ffb9ffbaffbbffbbffbcffbdffc0ffc4ffc7ffc9ffceffd3ff;
    inBuf[5255] = 256'hd6ffdaffdbffdbffdeffe0ffe2ffe5ffe6ffe5ffe8ffecffedffeffff4fff8ff;
    inBuf[5256] = 256'hfafffdfffeffffff00000300050007000a000e00110013001300150018001b00;
    inBuf[5257] = 256'h1c001c001d001d001e001e001f00220026002a002b002a002b002f0030003200;
    inBuf[5258] = 256'h360037003600340033003200350039003800350038003d003e003e003d003d00;
    inBuf[5259] = 256'h400040003e003e003e003c003d00410043004300430045004500440044004200;
    inBuf[5260] = 256'h3e004000430040003f0040003f0041004300420045004a004a00470045004200;
    inBuf[5261] = 256'h410041003f003e003f004000410040003f003e003d003d004100440045004300;
    inBuf[5262] = 256'h40003f003e004000420043004400450046004700470045004500460044004300;
    inBuf[5263] = 256'h430041004000400040004400470048004b004d004e0050004e004a004c004e00;
    inBuf[5264] = 256'h4d004d004d004d004f0050004f00500052005100510053005300540056005500;
    inBuf[5265] = 256'h5300540055005500560057005600570056005500540053005200550055005300;
    inBuf[5266] = 256'h530052005300560057005900590057005700580053004f004d004c004d005000;
    inBuf[5267] = 256'h4e004e004e004a00480049004700450044004300430040003b0039003a003a00;
    inBuf[5268] = 256'h3a0038003600390039003600340031002f0030002d002600240022001d001b00;
    inBuf[5269] = 256'h1a00180019001b001b001a001900150010000c00070006000800060003000300;
    inBuf[5270] = 256'h030001000000fdfffbfffcfffcfffcfffcfff8fff4fff0ffecffecffecffebff;
    inBuf[5271] = 256'heaffeaffe7ffe5ffe5ffe7ffeaffebffe9ffe9ffe7ffe3ffe2ffdeffd6ffd6ff;
    inBuf[5272] = 256'hd8ffdaffddffe0ffddffdcffdeffdeffddffdbffd8ffd8ffdaffd8ffd6ffd4ff;
    inBuf[5273] = 256'hd2ffd2ffd8ffdcffd9ffd6ffd6ffd5ffd4ffd4ffd4ffd4ffd5ffd4ffd5ffd3ff;
    inBuf[5274] = 256'hceffcdffd1ffd3ffd3ffd3ffd4ffd6ffd6ffd3ffd2ffd3ffd1ffd0ffd0ffceff;
    inBuf[5275] = 256'hceffceffceffcfffceffccffccffceffcdffcbffc9ffc7ffc6ffc6ffc4ffc2ff;
    inBuf[5276] = 256'hc2ffc4ffc5ffc6ffc7ffc7ffc7ffc5ffc2ffc2ffc2ffc2ffc2ffc2ffc2ffbfff;
    inBuf[5277] = 256'hbbffb9ffb5ffb1ffb0ffb1ffb0ffb1ffb4ffb5ffb7ffb6ffb4ffb5ffb5ffb4ff;
    inBuf[5278] = 256'hb4ffb4ffb1ffb0ffb1ffb0ffb1ffb2ffafffabffaaffa9ffa7ffa6ffa6ffa8ff;
    inBuf[5279] = 256'haaffaaffaaffacffabffaaffaaffaaffa9ffaaffabffabffaaffaaffacffacff;
    inBuf[5280] = 256'hacffb0ffb3ffb2ffb1ffb3ffb3ffb3ffb3ffb2ffb3ffb2ffb0ffb1ffb1ffafff;
    inBuf[5281] = 256'hb1ffb4ffb3ffb3ffb6ffb8ffbaffbcffbeffc0ffc2ffc1ffc3ffc4ffc2ffc3ff;
    inBuf[5282] = 256'hc9ffccffcbffcbffcdffccffcaffc8ffc8ffc9ffcaffcdffd3ffd6ffd6ffd9ff;
    inBuf[5283] = 256'hdbffdbffdcffdcffdbffdcffdaffdaffdeffdeffdfffe4ffe7ffe8ffedffedff;
    inBuf[5284] = 256'he9ffeaffeaffe8ffe9ffe9ffeaffeefff0ffeffff0fff1fff1fff3fff4fff4ff;
    inBuf[5285] = 256'hf3fff3fff4fff5fff5fff7fff8fff8fffafffdfffcfffbfffcfffdfffbfffcff;
    inBuf[5286] = 256'hfdfffefffdfffcfffcfffefffffffdffffff0300060008000800070007000600;
    inBuf[5287] = 256'h0300030005000600090008000700080006000000ffff00000200060007000800;
    inBuf[5288] = 256'h0c00100013001500120011001200100010000f000c000d001000110015001b00;
    inBuf[5289] = 256'h1b001b001e001e001e0020001d001b001c001c001c001d001e001e001f002000;
    inBuf[5290] = 256'h22002200240028002c00300032003200340038003b003a003b003e003f003d00;
    inBuf[5291] = 256'h3c003b003d003f003e003e00420043004100420042004300470049004d005300;
    inBuf[5292] = 256'h5600570059005a005a005b005c005e005f005d005b005d005f00620064006300;
    inBuf[5293] = 256'h640068006a0069006700660065006400650068006800680069006b006d007000;
    inBuf[5294] = 256'h720077007a007800760077007400720071006f006f0070007200740076007600;
    inBuf[5295] = 256'h7700770076007600760074007300740074007400730072007400740071007000;
    inBuf[5296] = 256'h730074007100710073007300740074007100700070007000700071006f006d00;
    inBuf[5297] = 256'h6c006c006b006b006b00690069006a00690069006c006e006c006d006f007000;
    inBuf[5298] = 256'h6f006d006900680068006600660064005f005e00600061006100620064006600;
    inBuf[5299] = 256'h67006600660066006600650065006600670068006a006a006800670065006200;
    inBuf[5300] = 256'h61005f005c005d006000600060005f005d005c005d005f0060005f005e005f00;
    inBuf[5301] = 256'h6300640060005f005f005e005c005d005f006100620064006600660065006500;
    inBuf[5302] = 256'h63005e005a00570053004f004d004d004e005000520056005a005c005e006100;
    inBuf[5303] = 256'h61005f005c005b005900550050004d004c004b004a004a0049004a004d004c00;
    inBuf[5304] = 256'h4c0050005300510050004d004a00470043004000400040003e003c003c003d00;
    inBuf[5305] = 256'h3a0038003700340034003800380037003a003900330030002d00290029002900;
    inBuf[5306] = 256'h29002b002d002e002e002c00270021001d001c001b00180018001a001a001a00;
    inBuf[5307] = 256'h1a001800150011000c0008000600040003000500060005000400060007000700;
    inBuf[5308] = 256'h06000500060004000100fffffbfffafffafff8fff5fff6fff4fff0fff1ffefff;
    inBuf[5309] = 256'he9ffe7ffe5ffe4ffe6ffe8ffe9ffebffedffecffecffebffe9ffe6ffe1ffdfff;
    inBuf[5310] = 256'hdeffdbffdaffdaffd8ffd8ffdaffd9ffd9ffdcffdcffdcffdcffd8ffd4ffd1ff;
    inBuf[5311] = 256'hcdffcaffc9ffcaffccffcdffcfffd2ffd3ffd3ffd1ffcfffcbffc9ffc8ffc7ff;
    inBuf[5312] = 256'hc7ffc7ffc7ffc5ffc5ffc3ffc1ffc0ffc0ffbfffc1ffc3ffc4ffc3ffc1ffbfff;
    inBuf[5313] = 256'hbcffb8ffb6ffb6ffb5ffb7ffb8ffb8ffbcffbfffbcffbbffbcffb9ffb6ffb5ff;
    inBuf[5314] = 256'hb2ffafffaeffacffaaffa8ffa8ffaaffacffaeffb2ffb3ffb2ffb3ffb2ffafff;
    inBuf[5315] = 256'hb0ffadffaaffabffabffa9ffaaffaaffa6ffa4ffa2ffa0ff9eff9cff9aff99ff;
    inBuf[5316] = 256'h99ff9aff99ff9aff9dffa1ffa3ffa5ffa7ffa7ffa6ffa4ffa2ffa0ff9dff9aff;
    inBuf[5317] = 256'h99ff99ff9aff9bff9dff9fff9dff98ff95ff93ff91ff8fff8eff8fff91ff94ff;
    inBuf[5318] = 256'h97ff97ff95ff95ff94ff93ff96ff98ff99ff9effa1ffa1ffa1ffa1ff9eff9bff;
    inBuf[5319] = 256'h9aff97ff97ff9aff9dff9eff9eff9fff9eff9bff99ff96ff94ff94ff94ff93ff;
    inBuf[5320] = 256'h97ff9bff9effa3ffa9ffafffb4ffb9ffbcffbeffbfffbdffb7ffafffaaffa6ff;
    inBuf[5321] = 256'ha4ffa3ffa5ffabffb0ffb6ffbdffc2ffc6ffc8ffc9ffc8ffc6ffc2ffc0ffc0ff;
    inBuf[5322] = 256'hc0ffc1ffc5ffcaffceffd4ffdaffddffdfffdfffdfffdcffd6ffd1ffceffcaff;
    inBuf[5323] = 256'hc6ffc8ffcfffd7ffdeffe3ffe7ffecfff0fff1fff2fff2fff0ffefffefffedff;
    inBuf[5324] = 256'heaffe8ffe6ffe5ffe8ffecfff0fff6fffafffcfffcfff9fff3ffebffe4ffe0ff;
    inBuf[5325] = 256'hdeffdfffe4ffecfff6ffffff05000c00110011000d0008000100fafff6fff3ff;
    inBuf[5326] = 256'hf2fff3fff5fffaff010005000600070006000100fcfff8fff3fff1fff0fff2ff;
    inBuf[5327] = 256'hf5fffcff030009000f00150018001b001e001c00180014000f000a0007000300;
    inBuf[5328] = 256'hfdfffcfffeff010006000f00190023002b002f002f002d0025001c0014000e00;
    inBuf[5329] = 256'h09000a000d0013001b0023002b003100350036003500320030002f002e002f00;
    inBuf[5330] = 256'h34003a004100460049004a0047003f0036002d0024001d001b001e0024002f00;
    inBuf[5331] = 256'h3e0050005f006a007100730072006d00630058004c0042003b00360033003500;
    inBuf[5332] = 256'h38003c0044004d00560060006a0072007b0080007f007e007b00720067005d00;
    inBuf[5333] = 256'h54004e004a0048004b00520057005c00610064006500630060005f0060006400;
    inBuf[5334] = 256'h6a0072007c0087008f00930093008e0083007500640051004100370033003900;
    inBuf[5335] = 256'h470058006d00830092009b009c00930085007400630058005300510054005b00;
    inBuf[5336] = 256'h62006b00720074007500730070006e006c006a006c006f007100730072006e00;
    inBuf[5337] = 256'h6900610059005300520054005b0063006c0075007900780074006e0067005f00;
    inBuf[5338] = 256'h580054005300540056005c006200660069006a0066005e0056004d0047004800;
    inBuf[5339] = 256'h4f005b006a00790085008900840076005f004300290014000800070011002400;
    inBuf[5340] = 256'h40005c0076008c009a009c00960087006f0054003a00230013000a0008000d00;
    inBuf[5341] = 256'h14001d0028003100380040004900510058005c005d0058004f00430037002b00;
    inBuf[5342] = 256'h2000190017001400120010000e000a0006000100fbfff4ffeeffecfff1fffaff;
    inBuf[5343] = 256'h0b002500400059006b006f00630047001e00eeffbeff95ff78ff6dff70ff82ff;
    inBuf[5344] = 256'ha0ffc4ffe9ff090021002d002d0022000e00f7ffdfffccffc0ffbaffbbffbfff;
    inBuf[5345] = 256'hc1ffc1ffbbffafffa1ff91ff84ff7fff80ff88ff95ffa6ffb7ffc5ffcfffd1ff;
    inBuf[5346] = 256'hceffc6ffbaffabff9dff8fff84ff7bff74ff70ff6eff6bff67ff64ff61ff61ff;
    inBuf[5347] = 256'h66ff71ff81ff95ffaaffbbffc3ffbeffaeff92ff6eff49ff29ff12ff09ff0dff;
    inBuf[5348] = 256'h1fff3aff5bff7bff95ffa5ffa8ff9dff85ff64ff41ff23ff0fff07ff0eff22ff;
    inBuf[5349] = 256'h3eff5bff72ff80ff82ff76ff62ff4bff32ff1cff0fff0aff0dff15ff1fff2bff;
    inBuf[5350] = 256'h36ff3cff3bff37ff31ff2aff26ff25ff2aff33ff3dff47ff4eff4bff40ff30ff;
    inBuf[5351] = 256'h1cff06fff3fee5fedefedffee8fef5fe03ff10ff18ff1dff20ff1eff1cff1bff;
    inBuf[5352] = 256'h1cff22ff2eff3aff46ff50ff52ff4aff38ff1cfff7fed1feb0fe98fe90fe98fe;
    inBuf[5353] = 256'haffed1fef8fe1dff3bff4eff54ff50ff45ff39ff30ff2eff34ff40ff4bff51ff;
    inBuf[5354] = 256'h4cff3aff1affeffebffe92fe73fe67fe73fe98fecffe13ff59ff96ffc2ffd8ff;
    inBuf[5355] = 256'hd4ffbcff94ff63ff31ff08ffe8fed2fecafecbfed1fedcfee8fef4fe03ff15ff;
    inBuf[5356] = 256'h2aff42ff5dff79ff93ffa7ffb1ffaeff9fff84ff61ff3aff17fffdfeeefeeefe;
    inBuf[5357] = 256'hfcfe14ff32ff50ff68ff78ff7eff7aff71ff68ff62ff64ff6eff7fff95ffabff;
    inBuf[5358] = 256'hbbffc3ffbfffadff92ff70ff4dff2fff1aff12ff18ff2cff4bff72ff9bffc2ff;
    inBuf[5359] = 256'he3fffcff080009000000edffd4ffb9ffa0ff8bff7fff7bff7fff8bff9cffafff;
    inBuf[5360] = 256'hc2ffd0ffdaffe0ffe1ffddffd7ffd0ffc9ffc5ffc3ffc5ffccffd9ffeaff0200;
    inBuf[5361] = 256'h1d003b0058006f007c007c006a0049001c00e7ffb5ff8dff76ff76ff8fffbcff;
    inBuf[5362] = 256'hf8ff380073009f00b600b700a3008000590037002200210036005c008d00be00;
    inBuf[5363] = 256'he200f300e900c5008a004200f9ffbdff96ff8effa7ffdeff2c008700e0002f01;
    inBuf[5364] = 256'h6b018c0192017f0159012501ec00b3007d004f002b0011000100fdff06001d00;
    inBuf[5365] = 256'h40007200af00f3003a017a01ae01d001d801c401960155010701b80071003b00;
    inBuf[5366] = 256'h1c0017002b0052008600bf00f50020013e014e01530152015001500157016401;
    inBuf[5367] = 256'h74018201870181016a0144011301dd00aa0082006900640074009500c500fd00;
    inBuf[5368] = 256'h37016d019b01bd01d301dc01db01d201c001a8018901630137010701d700ab00;
    inBuf[5369] = 256'h8b007b0080009d00cf0011015b01a501e4011102260221020402d40198015a01;
    inBuf[5370] = 256'h2201f600da00cf00d400e400fc001601300149015f01740188019a01ab01b901;
    inBuf[5371] = 256'hc101c101b701a40187016501430124010f0106010a0119013001490160017101;
    inBuf[5372] = 256'h7a017a0172016501560147013b01320130013501400150016301770188019601;
    inBuf[5373] = 256'h9e01a0019b01910181016e0155013a011c01ff00e500d100c400bf00c300cd00;
    inBuf[5374] = 256'hdd00f000070121013d015c017c019901b101c101c601bf01ac018f016b014001;
    inBuf[5375] = 256'h1101e000ae007d0051002c0012000500090020004a008600d20027017e01ce01;
    inBuf[5376] = 256'h0e02320236021502d3017401040190002500cfff97ff82ff8fffbafffaff4600;
    inBuf[5377] = 256'h9200d50009012a013801340123010a01ec00cc00ae0092007900630050003e00;
    inBuf[5378] = 256'h2d001f0013000c000c001500280045006a009200b900db00f30000010001f100;
    inBuf[5379] = 256'hd400a9006f002800d8ff87ff3bfffefedafed5fef1fe2fff8afff9ff7200e900;
    inBuf[5380] = 256'h5201a201d001d401ae015f01f0006c00e3ff64fffbfeb3fe8efe8efeacfee2fe;
    inBuf[5381] = 256'h26ff6fffb6fff2ff1e00390043003e00310024001b001c0029003f0058006d00;
    inBuf[5382] = 256'h76006d0050001e00dbff91ff47ff07ffd9fec2fec4feddfe08ff3dff74ffa4ff;
    inBuf[5383] = 256'hc7ffd8ffd5ffc3ffa5ff83ff66ff54ff56ff6cff97ffd0ff0f00490072008400;
    inBuf[5384] = 256'h77004d000900b0ff4effeafe8efe45fe14fe02fe0ffe3afe7efed2fe2bff80ff;
    inBuf[5385] = 256'hc7fffbff1900220019000300e4ffc2ffa0ff84ff70ff65ff64ff6aff73ff78ff;
    inBuf[5386] = 256'h74ff62ff41ff13ffdcfea5fe76fe55fe49fe52fe71fea2fee1fe28ff71ffb4ff;
    inBuf[5387] = 256'hebff0f001a000b00e4ffacff6bff2efffefee5fee6fe02ff35ff75ffb7fff0ff;
    inBuf[5388] = 256'h12001500f2ffaaff42ffc6fe42fecafd6cfd37fd34fd67fdcefd60fe0fffc8ff;
    inBuf[5389] = 256'h78000c017301a4019a015901e8005600b4ff12ff82fe11fecafdb0fdc2fdf9fd;
    inBuf[5390] = 256'h49fea3fef9fe3eff6cff7fff7cff68ff4cff2eff14ff04ff01ff0cff27ff50ff;
    inBuf[5391] = 256'h84ffbdfff4ff2200400049003d001f00f1ffb9ff7dff3fff05ffd2fea7fe87fe;
    inBuf[5392] = 256'h74fe6efe75fe84fe99feb0fec5fed7fee8fefafe0fff2cff51ff7effb4ffeeff;
    inBuf[5393] = 256'h2b0067009d00c900e700ef00dd00ae005f00f3ff6fffdcfe43feb0fd31fdd0fc;
    inBuf[5394] = 256'h98fc91fcbffc23fdb7fd74fe4bff2c000401bf014b029902a3026702eb013d01;
    inBuf[5395] = 256'h6f0096ffc8fe18fe94fd46fd31fd52fd9ffd0afe82fef5fe52ff8fffa5ff98ff;
    inBuf[5396] = 256'h71ff3cff0dfff1fef8fe27ff7ffff8ff83000e018401d101e601ba014c01a500;
    inBuf[5397] = 256'hd6fff7fe21fe70fdf8fcc9fce7fc49fde1fd95fe4efff2ff6f00b800cb00ab00;
    inBuf[5398] = 256'h630003009cff43ff08fff6fe15ff62ffd4ff5900dd004a018c0197016601fb00;
    inBuf[5399] = 256'h6300adfff0fe42feb7fd60fd45fd69fdc4fd49fee4fe7fff08006f00ad00bf00;
    inBuf[5400] = 256'had00820049001100e6ffd1ffd7fff7ff2d007100b600f2001b0128011501e000;
    inBuf[5401] = 256'h8d002000a1ff18ff90fe13feadfd65fd44fd4efd86fde9fd75fe21ffe4ffb000;
    inBuf[5402] = 256'h76012802b4020d032a030603a202070243016a0090ffcbfe2bfebdfd86fd86fd;
    inBuf[5403] = 256'hb4fd08fe73fee7fe54ffaeffecff0b000d00fcffe5ffd7ffe0ff09005400bd00;
    inBuf[5404] = 256'h3901b70123026a027c024e02db012901450045ff46fe63fdb8fc5afc54fca7fc;
    inBuf[5405] = 256'h4bfd2dfe34ff41003801fd017c02ab02890220028301cb00120074ff04ffd2fe;
    inBuf[5406] = 256'he4fe34ffb4ff4e00e7006101a501a0014c01ae00d8ffe4fef1fd22fd94fc5dfc;
    inBuf[5407] = 256'h89fc19fdfffd25ff6a00a801bc028503ed03e8037b03b702b7019e008fffaafe;
    inBuf[5408] = 256'h07feb7fdbafd08fe8ffe34ffdbff6700c400e100bc005a00cbff26ff85fe04fe;
    inBuf[5409] = 256'hbbfdb9fd07fea0fe75ff6e0070015c0216038703a1035d03bf02d801c00099ff;
    inBuf[5410] = 256'h85fea6fd19fdebfc20fdabfd74fe5bff3b00f200660188015701de0035007bff;
    inBuf[5411] = 256'hd2fe57fe1ffe38fe9efe45ff1800f900cc017702e4020a03e3027702d2010601;
    inBuf[5412] = 256'h290051ff91fef9fd96fd6efd82fdcdfd45fedcfe81ff2200ae0015014f015801;
    inBuf[5413] = 256'h3501f1009b0046000200ddffddff03004800a000fc004b017d0185015901fa00;
    inBuf[5414] = 256'h6f00c7ff17ff77fefdfdb7fdaefde0fd46fed2fe76ff2200c9006001de013f02;
    inBuf[5415] = 256'h7f029b029102600208028a01ec00350073ffb4fe0afe86fd39fd2ffd6efdf3fd;
    inBuf[5416] = 256'hb2fe96ff83005b0100025e026a022902a90104015b00cdff75ff63ff99ff0e00;
    inBuf[5417] = 256'haa005101e2013d024b02fd0153015c0035ff06fefbfc3ffcf3fb2afce4fc0dfe;
    inBuf[5418] = 256'h83ff17019702d203a304f004b004eb03bc024901c0ff54fe33fd81fc54fcb0fc;
    inBuf[5419] = 256'h87fdbafe1f008601c102a7031e04170492039e025901e8ff7afe3dfd5efcfcfb;
    inBuf[5420] = 256'h29fce1fc0bfe7dff020160026403ec03e8035c0362022301d0ff9efebafd49fd;
    inBuf[5421] = 256'h5dfdf6fdfffe5300c30118031f04af04ad041104e802540184ffb3fd1dfcf5fa;
    inBuf[5422] = 256'h63fa79fa35fb7ffc2ffe1300f2019403cd047a058f050d050d04b2022b01a7ff;
    inBuf[5423] = 256'h55fe5bfdd3fcc8fc37fd0cfe25ff5a007b015d02dd02e402700292016e0036ff;
    inBuf[5424] = 256'h1ffe5bfd0ffd49fd01fe1aff6600b101c6027f03c0038503d902d601a20066ff;
    inBuf[5425] = 256'h49fe6efdeefcd3fc1efdc2fda7feafffba00ab016b02ed022b032903ee028302;
    inBuf[5426] = 256'hf5014f019d00eaff41ffaefe39feeafdc7fdd0fd07fe67fee7fe7dff1700a600;
    inBuf[5427] = 256'h190164018201750147010801c7009400770074008800ab00d400f8000d010b01;
    inBuf[5428] = 256'hec00af005700ecff79ff0affabfe66fe43fe47fe75fecdfe4dffecff9f005301;
    inBuf[5429] = 256'hf6017202b602b7027102e80125013b0040ff4dfe7afde2fc99fcb0fc2efd0efe;
    inBuf[5430] = 256'h40ffa400110258034d04ce04c70438043403da015800dcfe94fda8fc31fc3afc;
    inBuf[5431] = 256'hbafc98fdadfecbffc6007b01d501ce017301dc002b0083ff02ffc0fec6fe14ff;
    inBuf[5432] = 256'h9dff4e000d01c1015002a902c002920224028301c000eeff20ff68fed7fd7bfd;
    inBuf[5433] = 256'h5dfd83fde9fd85fe45ff1200d2006c01cf01ed01c5015f01cd00280089ff0cff;
    inBuf[5434] = 256'hc4febdfef8fe6afffeff9a0023018201a90195014e01e2006500ebff85ff40ff;
    inBuf[5435] = 256'h26ff38ff74ffcfff37009700dc00f400da008f002000a0ff23ffbcfe77fe5bfe;
    inBuf[5436] = 256'h65fe90fed4fe29ff89fff1ff5e00ce003d01a501ff014202680269024302f301;
    inBuf[5437] = 256'h7a01dd00270065ffabfe0dfe9afd60fd63fd9ffd0cfe9cfe3effe2ff7800f300;
    inBuf[5438] = 256'h4b017e018d017b014e010d01bf0068001100beff78ff43ff25ff23ff3dff71ff;
    inBuf[5439] = 256'hbaff0f006300ac00de00f300e700bf0080003700eeffb1ff89ff7eff8fffb7ff;
    inBuf[5440] = 256'hebff1d003e0044002a00f3ffaaff5cff15ffe1fec4febefecffef4fe2dff79ff;
    inBuf[5441] = 256'hdaff4c00c6003d019f01e001f501de01a1014b01e80083002200caff7bff37ff;
    inBuf[5442] = 256'h00ffdafec8feccfee4fe0dff3eff70ff98ffafffb1ff9dff78ff4bff22ff0bff;
    inBuf[5443] = 256'h11ff40ff9bff2200cc0086013a02cc0223032a03d90231024201290006fffffd;
    inBuf[5444] = 256'h39fdcefccdfc36fdf7fdf5fe0a000f01e20166028d025202be01e700ecfff1fe;
    inBuf[5445] = 256'h1cfe89fd4afd63fdc9fd67fe24ffeaffa7005101e3015902b102e402e802b602;
    inBuf[5446] = 256'h4902a701e0000c0046ffa7fe41fe18fe27fe61feb5fe10ff65ffa9ffd7ffecff;
    inBuf[5447] = 256'he7ffceffa9ff85ff6eff73ff9efff1ff6800f600860105025c027d025e02fe01;
    inBuf[5448] = 256'h62019800b4ffd1fe0cfe81fd49fd6ffdf6fdccfed8fff300f801c00232033f03;
    inBuf[5449] = 256'he70237024901390028ff30fe66fddafc93fc97fce5fc79fd4afe48ff5e007001;
    inBuf[5450] = 256'h640220039003ac037303f10238025e017c00a7fff1fe6bfe1ffe13fe4bfebdfe;
    inBuf[5451] = 256'h59ff0600a50019014c013401d700440094ffe2fe47fed8fda5fdb8fd15feb6fe;
    inBuf[5452] = 256'h90ff8c008e017602250380037a0310034f025001320019ff27fe75fd16fd15fd;
    inBuf[5453] = 256'h72fd25fe1bff3a005e015f021603650337038d0278011b00a3fe45fd2ffc89fb;
    inBuf[5454] = 256'h68fbd3fbbcfc07fe8bff17017c028c0327043c04ca03e702b501620021ff20fe;
    inBuf[5455] = 256'h84fd60fdb7fd74fe73ff86007a0125026a023b02a101b1008cff57fe3bfd5dfc;
    inBuf[5456] = 256'hdcfbcffb40fc27fd6dfeeeff7701d802e3037804870414042f03f301840007ff;
    inBuf[5457] = 256'ha4fd81fcc1fb82fbd4fbb2fc04fe9cff3f01ae02b503310419047b0377023501;
    inBuf[5458] = 256'he3ffaafeaefd07fdc3fce2fc54fd01fec6fe81ff1100630070004000e5ff7bff;
    inBuf[5459] = 256'h20ffedfef4fe3affbbff69002d01f0019802100346032f03ca021b022e011800;
    inBuf[5460] = 256'hf0fed1fdd3fc0efc91fb69fb97fb17fcdcfcd4fdecfe0d0024011d02e5026a03;
    inBuf[5461] = 256'h9e037703f1021602fa00bfff8efe8ffde4fca2fccdfc58fd2dfe2bff33002601;
    inBuf[5462] = 256'hec016e029e027502f701330144004bff6afebefd57fd34fd4bfd8afde0fd3ffe;
    inBuf[5463] = 256'ha0fe01ff64ffc9ff2e008e00e30026015101620158013201f2009a002f00baff;
    inBuf[5464] = 256'h47ffe7fea8fe94feadfee9fe39ff87ffc1ffdcffd4ffadff73ff37ff09fff6fe;
    inBuf[5465] = 256'h07ff3cff8effecff43007d008b0064000a008bfff9fe6bfef9fdb6fdb0fdeffd;
    inBuf[5466] = 256'h72fe2fff12000201de018602dc02cd02550280016d0044ff30fe5afddcfcc2fc;
    inBuf[5467] = 256'h07fd9bfd66fe4cff3100f9008901cd01b6014001770072ff58fe50fd85fc14fc;
    inBuf[5468] = 256'h12fc83fc5dfd8afeecff5e01b702cd037c04a60443045b030f028e000fffc7fd;
    inBuf[5469] = 256'hddfc64fc5cfcb1fc44fdf2fd9bfe27ff86ffb4ffb4ff92ff5fff2cff0dff13ff;
    inBuf[5470] = 256'h47ffacff3700d7007401f20138023502e4014c018200a1ffcdfe26fec7fdbdfd;
    inBuf[5471] = 256'h06fe92fe43fff5ff8a00ea000a01ee009d0028009cff09ff7ffe10fecdfdc4fd;
    inBuf[5472] = 256'hfefd78fe24ffeaffaf005901d40116021b02e6017f01f1004a009cfffafe7cfe;
    inBuf[5473] = 256'h31fe22fe4dfea5fe12ff80ffdbff1c0044005b006a007700810085007d006700;
    inBuf[5474] = 256'h45001e00faffdeffccffbdffa9ff87ff54ff13ffcefe95fe78fe85fec5fe37ff;
    inBuf[5475] = 256'hd1ff81003101c7012d0254023702de015701b9001b0090ff26ffe2fec1febffe;
    inBuf[5476] = 256'hd2fef4fe1eff4eff81ffb6ffedff25005a008900af00c600cc00bc0095005900;
    inBuf[5477] = 256'h0d00b9ff6cff32ff18ff27ff5fffbaff2c00a50016017301b501d901db01bc01;
    inBuf[5478] = 256'h7d012101b1003700c3ff61ff17ffe4fec3feaafe94fe80fe76fe81feaefe04ff;
    inBuf[5479] = 256'h83ff2300d300810118028702bf02ba02790203026a01c3002500a6ff56ff39ff;
    inBuf[5480] = 256'h4bff81ffc8ff0b00390048003100f8ffaaff57ff13fff3fe06ff52ffd4ff7c00;
    inBuf[5481] = 256'h3301dc015a02970289023202a001e70023006effe0fe8bfe7bfeb3fe2cffd5ff;
    inBuf[5482] = 256'h93004701cf0114020902b20126018400eeff83ff52ff61ffa4ff09007a00e300;
    inBuf[5483] = 256'h35016601720157011801bb004a00d4ff69ff1cfffbfe0aff47ffa8ff1e009b00;
    inBuf[5484] = 256'h14018101dc01210249024e022902d9016501d8004200b5ff3effe8feb7feb1fe;
    inBuf[5485] = 256'hd6fe27ff9fff3400d5006d01e10120021c02d8015d01c200210093ff31ff0aff;
    inBuf[5486] = 256'h25ff7dff0400a1003601a901e601e801b50160010001a800650038001a000000;
    inBuf[5487] = 256'he3ffc3ffa5ff93ff97ffb5ffeaff2c006e00a600cc00e000e300dc00cf00bf00;
    inBuf[5488] = 256'hb100a500a100a900bc00d700f100fa00e400a7004200c2ff3cffc8fe7efe6efe;
    inBuf[5489] = 256'h9efe0fffb4ff80005d013102df024f03690325038702a201940080ff8afecdfd;
    inBuf[5490] = 256'h59fd35fd5afdbdfd4bfef0fe9aff3900c1002d018101c001f2011a0238024402;
    inBuf[5491] = 256'h35020302ac013601ad002400aaff49ff02ffcffea7fe83fe63fe4bfe47fe60fe;
    inBuf[5492] = 256'h9afef5fe69ffeaff6d00e9005a01be0110024b02650256021602a30106014d00;
    inBuf[5493] = 256'h8effe2fe5afe06feeafd04fe4cfeb5fe32ffb3ff2b008c00cf00ef00f200e100;
    inBuf[5494] = 256'hca00b900b400b800b900a6006f000c0080ffdffe44fed0fd9dfdbcfd2ffee7fe;
    inBuf[5495] = 256'hcbffbb009301370292029a025302ce0123016c00bfff2effc0fe76fe50fe4afe;
    inBuf[5496] = 256'h61fe8efecafe06ff34ff4bff48ff33ff20ff24ff54ffb8ff4a00f600a0012702;
    inBuf[5497] = 256'h71026d0219027e01b100cbffe7fe1ffe85fd27fd08fd26fd75fde7fd6bfef3fe;
    inBuf[5498] = 256'h77fff2ff6600d60040019f01e4010102e6018b01f60037006cffb2fe26fed8fd;
    inBuf[5499] = 256'hcbfdf4fd40fe98fee8fe24ff45ff4dff42ff2bff0efff6feecfefdfe34ff9bff;
    inBuf[5500] = 256'h3300f600d001a6025303b303a403130300027f00bbfeedfc57fb30faa1f9b7f9;
    inBuf[5501] = 256'h65fa89fbf5fc78feeaff3001390200038103bd03b5036c03e802350263018300;
    inBuf[5502] = 256'ha3ffd1fe17fe7efd10fdd6fcd5fc0dfd75fdfcfd8bfe11ff82ffdcff23006000;
    inBuf[5503] = 256'h9500c000d700d100a80061000700b0ff6fff52ff5cff85ffbbffe9fffbffe7ff;
    inBuf[5504] = 256'hb0ff65ff1bffe9fee3fe0cff5dffc3ff240067007c005f001600b3ff4bfff2fe;
    inBuf[5505] = 256'hb5fe99fe9bfeb3fedcfe12ff57ffafff1b00970015018201c701d00192010c01;
    inBuf[5506] = 256'h4b0066ff78fea1fdfefca8fcadfc14fdd3fdd3feeffffe00d501570279024202;
    inBuf[5507] = 256'hd0014301be0055000f00e1ffb9ff86ff3bffd9fe68fefafd9ffd67fd5bfd7ffd;
    inBuf[5508] = 256'hd5fd5afe0bffdfffc800ae017402fa022303e00235023c01200017ff52fef6fd;
    inBuf[5509] = 256'h11fe96fe60ff3d00f5005d015701e300130011ff0efe3bfdc1fcb6fc20fdedfd;
    inBuf[5510] = 256'h00ff300050013902cc02f802bd022d0263018300afff02ff8ffe5bfe64fea3fe;
    inBuf[5511] = 256'h10ffa2ff51000d01c201510299027c02e601de0081ff04fea9fcacfb3afb61fb;
    inBuf[5512] = 256'h15fc32fd8afef1ff460173026b0324049504b3047204d303e002b10169002fff;
    inBuf[5513] = 256'h24fe5ffde9fcc1fcdafc27fd97fd1bfea4fe2bffa7ff15007700d00024017701;
    inBuf[5514] = 256'hcb011e026c02aa02cd02c7028d021d027901af00d6ff04ff4dfec1fd67fd41fd;
    inBuf[5515] = 256'h4dfd89fdf4fd8afe42ff0f00da008901060240023402f4019a014a0123013401;
    inBuf[5516] = 256'h7901d801290244020d027f01aa00b3ffc5fe03fe82fd45fd44fd6cfdaffd04fe;
    inBuf[5517] = 256'h6cfeebfe83ff3300f200b0015b02e6024a0386039c038e035803f30259028d01;
    inBuf[5518] = 256'h990097ffa6fee2fd5ffd22fd25fd5afdb4fd27feadfe43ffe4ff88002201a201;
    inBuf[5519] = 256'hfc01290229020502cc018a014e011c01f200ca009e006c0036000800eefff5ff;
    inBuf[5520] = 256'h1d005f00a800e000ed00c1005c00cdff31ffa6fe48fe23fe37fe74fecafe2bff;
    inBuf[5521] = 256'h92ff04008d003201ed01ae025603c703e803ad031b0348024e014a0053ff7bfe;
    inBuf[5522] = 256'hccfd52fd13fd17fd60fde8fd9bfe61ff1800a500f7000e01fa00d600bb00bc00;
    inBuf[5523] = 256'he10020016b01b401f1011f023f0250024b022202c6012b0153004bff32fe2ffd;
    inBuf[5524] = 256'h67fcf7fbeefb46fceefccbfdc2febdffb100950167022203bd032a045c044704;
    inBuf[5525] = 256'heb0353038c02aa01c100ddff01ff31fe6dfdbbfc27fcc6fbb0fbf8fba5fcacfd;
    inBuf[5526] = 256'hf4fe5400a201bb028503f8031804ed038303e6021c0234013d004fff86fefcfd;
    inBuf[5527] = 256'hbffdd2fd2afeacfe40ffcfff4b00af00fc002c013a011e01cf004e00abff02ff;
    inBuf[5528] = 256'h75fe25fe26fe78fe0bffbfff73000d017f01cc01fd011e0235023e022a02e801;
    inBuf[5529] = 256'h7101c300edff08ff31fe83fd13fde7fcfcfc4cfdc7fd62fe11ffccff8c004701;
    inBuf[5530] = 256'hf2018002e70218030b03c20242029801d5000a0042ff88fee3fd5ffd08fdeefc;
    inBuf[5531] = 256'h1efd9efd62fe53ff50003501e301490263023702d20140019000d1ff12ff65fe;
    inBuf[5532] = 256'he5fda9fdc4fd3dfe08ff090018010402a902ee02cf025902a701d200efff0fff;
    inBuf[5533] = 256'h3afe79fdd8fc69fc41fc73fc06fdf0fd18ff58008501790218035b034803f102;
    inBuf[5534] = 256'h6b02ce012a018a00f5ff6efff8fe94fe41fe00fed2fdb7fdb3fdccfd07fe68fe;
    inBuf[5535] = 256'hf0fe94ff4300e9006b01b701c30192013701cb006900250008000a0018001d00;
    inBuf[5536] = 256'h0400c5ff66fffbfe9ffe6dfe77febdfe32ffbcff3e009f00ce00c80095004000;
    inBuf[5537] = 256'hd7ff68fffffeaafe7afe7ffec4fe48fff8ffb8006001cc01e301a00114015c00;
    inBuf[5538] = 256'h9efffffe96fe6efe82fec3fe1bff75ffbdffe8ffefffd6ffa5ff6cff3cff2bff;
    inBuf[5539] = 256'h48ff9bff1b00b4004201a201b7017501e400210051ff9dfe22feeefd01fe4cfe;
    inBuf[5540] = 256'hbafe36ffb1ff1e007800be00ed000201f700c7007100f8ff69ffd9fe63fe20fe;
    inBuf[5541] = 256'h25fe79fe12ffd9ffaa005d01cf01e901a5010d013f005dff8efef3fda3fdaafd;
    inBuf[5542] = 256'h03fe9efe63ff3200ea0069019e01830120018e00edff5ffffdfed0fed5fe01ff;
    inBuf[5543] = 256'h41ff84ffbdffe6fffeff0300f7ffe0ffc4ffb3ffb6ffd9ff1c007300c9000201;
    inBuf[5544] = 256'h0301c0003b0089ffcafe27fec2fdb2fdfcfd92fe5fff3e000d01ae010b021802;
    inBuf[5545] = 256'hd6015301a500edff43ffbefe6afe47fe4efe73feaefef6fe48ffa2ffffff5a00;
    inBuf[5546] = 256'haa00e60008011001fc00d3009d005f002200eaffb9ff91ff6fff51ff32ff11ff;
    inBuf[5547] = 256'hedfeccfeb5feb2fed1fe1bff8fff2400c9006601df011d021302c00131017600;
    inBuf[5548] = 256'haaffe9fe48fedafda8fdb4fdfdfd78fe12ffbaff5f00f0006301b201d801da01;
    inBuf[5549] = 256'hb6016c0101017c00e6ff4dffc2fe53fe0efef7fd0ffe50feb3fe2affadff3000;
    inBuf[5550] = 256'hab0017016c01a301b801a80171011701a5002600a5ff2dffc6fe78fe48fe39fe;
    inBuf[5551] = 256'h52fe95fefffe88ff2400c4005501c901120227020602ac011d0164008fffb3fe;
    inBuf[5552] = 256'hebfd50fd00fd0ffd7efd43fe47ff63006d014302cb02fd02dd027902e5013701;
    inBuf[5553] = 256'h8100d1ff35ffb6fe5bfe2bfe24fe45fe85fedafe35ff8cffd6ff110040006800;
    inBuf[5554] = 256'h9400ca000c0151018c01af01a901710106017100c8ff1eff90fe34fe1afe48fe;
    inBuf[5555] = 256'hbafe5dff1800cc005801a501a7015e01dc003b009aff1affcffec1fee9fe38ff;
    inBuf[5556] = 256'h96fff1ff40007f00b400e60016014301630169014c010801a1002400a4ff30ff;
    inBuf[5557] = 256'hd8fea3fe8ffe97feb6fee8fe2aff7cffdeff4a00ba001f017201ab01c901ce01;
    inBuf[5558] = 256'hbc0192014f01f1007600e5ff4dffc0fe51fe12fe0ffe49feb9fe50fff9ffa000;
    inBuf[5559] = 256'h2c018801ab0190013f01c6003e00beff5eff2fff3eff8aff07009f003701ac01;
    inBuf[5560] = 256'he201ca016401c100fdff3dffa3fe4afe39fe6cfecffe48ffbbff180056007800;
    inBuf[5561] = 256'h8b009900a900bf00d600e600ee00ea00dd00ca00b4009d00840069004d003300;
    inBuf[5562] = 256'h1c000600eeffcfff9fff5eff11ffc4fe89fe73fe92feeffe84ff3f000701bd01;
    inBuf[5563] = 256'h4302880284023e02c70135019a0008008bff29ffe6fec2febefed8fe0fff5dff;
    inBuf[5564] = 256'hbcff24008800df001f01410144012b01f700ab004a00d8ff5cffe2fe7cfe41fe;
    inBuf[5565] = 256'h43fe8afe17ffdcffbe009e015d02e40224031a03ca023d028201a300b2ffc4fe;
    inBuf[5566] = 256'hecfd43fddefcc9fc08fd93fd56fe3bff27000101b7013c028a029e027a022402;
    inBuf[5567] = 256'ha70112017600eeff8eff61ff69ff9cffe2ff20003f003000f4ff98ff32ffe0fe;
    inBuf[5568] = 256'hb6febffefafe5effd6ff4e00b600040132013e012a01fc00c0007c003f001200;
    inBuf[5569] = 256'hfcfffbff0d00270040004f004d003d0025000d00fffffdff02000500f7ffccff;
    inBuf[5570] = 256'h80ff1fffbbfe6dfe51fe75fedffe85ff53002c01f8019f0213034a033e03f102;
    inBuf[5571] = 256'h6802a501b400a6ff8dfe81fd99fceefb95fb9bfb05fcd2fcf6fd5bffe4007102;
    inBuf[5572] = 256'hd903f3049c05b50536052804ab02ee0029ff93fd55fc8efb46fb79fb17fc06fd;
    inBuf[5573] = 256'h26fe5aff810083014e02d4020e030103b20230028c01d800260087ff00ff96fe;
    inBuf[5574] = 256'h4dfe23fe1afe35fe74fed6fe52ffdfff6c00ec0050018d01a301930162011c01;
    inBuf[5575] = 256'hca0072001700baff5eff05ffb5fe75fe51fe52fe77fec2fe2affa5ff25009d00;
    inBuf[5576] = 256'h000146016901660142010701bf0079004200200011000f000b00f8ffc8ff77ff;
    inBuf[5577] = 256'h0cff9afe37fefefd07fe56fee2fe98ff580003017e01ba01b7017f011f01ab00;
    inBuf[5578] = 256'h3800d1ff84ff55ff46ff56ff80ffb8fff5ff2b0051005e004f002400e3ff97ff;
    inBuf[5579] = 256'h46ff00ffcdfeb5febcfee6fe2fff95ff0f008e0003015f019101920164010a01;
    inBuf[5580] = 256'h96001a00a4ff41fffcfed2febffebefec8fedcfef9fe21ff59ffa1fff1ff4200;
    inBuf[5581] = 256'h8e00cd00fe002201360138012401ed008e00090066ffb5fe10fe93fd57fd6afd;
    inBuf[5582] = 256'hcdfd77fe52ff3c001501c301350263024f0201028901f3004d00a8ff16ffa2fe;
    inBuf[5583] = 256'h56fe36fe39fe57fe88febffef9fe36ff75ffb6fff5ff2b0058007b009700b000;
    inBuf[5584] = 256'hd300010137016c01910193016101ee00400069ff86feb8fd23fddcfcebfc4afd;
    inBuf[5585] = 256'he5fda5fe75ff3c00e7006e01cb01fd010b02fa01d0018f013501c1003900a5ff;
    inBuf[5586] = 256'h0eff85fe16fecafdaafdb7fdf3fd5cfeeafe8cff3400cd0044018c01a2018a01;
    inBuf[5587] = 256'h54010b01bb0070002900e2ff97ff47fff6feb0fe7cfe65fe71fe9dfee1fe38ff;
    inBuf[5588] = 256'h9bff06007800e70048019001b1019f015901e8005e00cdff48ffdefe9dfe84fe;
    inBuf[5589] = 256'h8bfeaefee1fe1bff57ff94ffd3ff1b006800b500fd003101460138010101a700;
    inBuf[5590] = 256'h3700bcff47ffebfeb6feaefed5fe1fff7dffdfff3100680081007e0064003f00;
    inBuf[5591] = 256'h1c0006000300150035005a00740075005c002c00eeffafff7bff57ff45ff42ff;
    inBuf[5592] = 256'h48ff5aff75ff97ffc6ff02004a009b00ea0029014b0144010e01af003300acff;
    inBuf[5593] = 256'h30ffccfe8bfe7afe9bfee9fe60fff3ff900020018a01c001ba017501fa005f00;
    inBuf[5594] = 256'hbcff29ffbbfe82fe7ffeadfefcfe5cffbdff15005e009800c300e100f200f800;
    inBuf[5595] = 256'hf200e500d400c000a700850052000a00adff47ffeafea9fe93feb1fefdfe66ff;
    inBuf[5596] = 256'hd9ff4700a000e00004010e010201e300b700850051001f00f1ffc7ffa6ff92ff;
    inBuf[5597] = 256'h92ffa8ffd6ff120050008300a100a50093006e003c000300caff98ff75ff66ff;
    inBuf[5598] = 256'h72ff97ffcfff0c0043006b007d007400540029000000e7ffecff15005b00ac00;
    inBuf[5599] = 256'hf3001f0127010701cc007f002600c7ff66ff0affbbfe87fe7dfea4fefafe73ff;
    inBuf[5600] = 256'h00008e0009016601a101b901b20192015b010f01b0004000c7ff51ffeefeadfe;
    inBuf[5601] = 256'h96fea7fed9fe23ff78ffd2ff2e008b00e6003a017d01a501ad018f014e01ef00;
    inBuf[5602] = 256'h7b0000008bff25ffddfebafebbfedbfe12ff57ffa3fff1ff3c008600ce000d01;
    inBuf[5603] = 256'h3e015e01660155012f01f600b60073002a00dcff8dff3dfff6fec7febdfeddfe;
    inBuf[5604] = 256'h20ff7affddff3e009000d700150144015f015f013e01fe00a3003900cfff73ff;
    inBuf[5605] = 256'h2aff00fffafe15ff4cff99ffedff3f008a00cb0001012b0144014a0136010301;
    inBuf[5606] = 256'hb90062000600acff5cff1bffeafecbfebefec7fee7fe19ff60ffbdff3000b500;
    inBuf[5607] = 256'h4101c101250258024c020402900100016900dbff61ff04ffc9feaffeb8fee0fe;
    inBuf[5608] = 256'h17ff52ff85ffa9ffbfffcfffe0ffffff32007900ce0025016c01930191016301;
    inBuf[5609] = 256'h1501b8005600fdffb3ff74ff42ff21ff13ff1aff3aff6cffadfff8ff43008b00;
    inBuf[5610] = 256'hc600e800f100e100bc0090006b0050003b0025000700e1ffb2ff7fff58ff46ff;
    inBuf[5611] = 256'h46ff57ff7dffafffe7ff23006400ac00fc0048018901b201af017b011b019a00;
    inBuf[5612] = 256'h0c0080ff00ff92fe3dfe07fefffd30fe9afe37fff2ffab004801b601ed01f201;
    inBuf[5613] = 256'hd20196014f010601b70067001500bbff59fff3fe93fe49fe27fe38fe85fe0bff;
    inBuf[5614] = 256'hb6ff71002501b8011c0249023b02f5018401f2005200b7ff2cffc0fe7bfe5ffe;
    inBuf[5615] = 256'h6cfe9ffeeafe45ffa4fffbff46008a00c400f4001801270124010f01ea00c000;
    inBuf[5616] = 256'h99007400510031000f00eaffbeff8bff55ff25ff07ff09ff2dff66ffa6ffddff;
    inBuf[5617] = 256'h000015002b004e007d00a900bf00b800950060002e0012000b00120022003400;
    inBuf[5618] = 256'h4a0060006e006a004e001300c8ff80ff4dff38ff41ff60ff89ffb7ffe4ff0f00;
    inBuf[5619] = 256'h300040003b0028000c00f4ffebfff2ff05001e003b005b007c00920096008100;
    inBuf[5620] = 256'h52001800e7ffd0ffd5ffe9fff7fff0ffd2ffa9ff8bff83ff90ffa7ffb7ffb7ff;
    inBuf[5621] = 256'habffa0ffa2ffb6ffd7ffffff27004c0071009600b300c000b7009b006f003f00;
    inBuf[5622] = 256'h1300ebffbfff8dff59ff2dff10ff09ff18ff38ff60ff8dffbffff7ff30006300;
    inBuf[5623] = 256'h880096008f00770054002a00fdffd4ffb4ffa3ffa6ffbaffd8ffeffff4ffe5ff;
    inBuf[5624] = 256'hc9ffa7ff88ff74ff6eff77ff8bffa8ffccffedff020008000600010000000300;
    inBuf[5625] = 256'h07000400f2ffd6ffbeffb6ffc0ffd8ffeffff4ffe1ffbbff8eff66ff49ff36ff;
    inBuf[5626] = 256'h2dff2eff3fff6affaefffeff4c0086009f0098007e005c0037001000e5ffb8ff;
    inBuf[5627] = 256'h8aff5eff3eff2bff1fff1aff1dff27ff3aff53ff6bff81ff93ffa6ffbeffdbff;
    inBuf[5628] = 256'hf7ff0d001a00220035005e009100bd00c40093002e00a9ff26ffc5fe93fe86fe;
    inBuf[5629] = 256'h94feb3fedcfe13ff56ff9bffd9ff020010000b00fcffe9ffd8ffc9ffb9ffb0ff;
    inBuf[5630] = 256'hb0ffb9ffccffddffe3ffdfffd0ffb9ffa1ff8bff70ff57ff44ff3eff4cff69ff;
    inBuf[5631] = 256'h8cffabffbbffb8ffacff9dff88ff72ff5aff3fff29ff20ff2bff4aff70ff92ff;
    inBuf[5632] = 256'hafffc6ffd9fff5ff1b00410061006e0061003a00fbffa5ff44ffe1fe8afe56fe;
    inBuf[5633] = 256'h4ffe6ffeb1fefdfe3dff6fff97ffc1fff5ff2e005c00730069003c000000c2ff;
    inBuf[5634] = 256'h85ff49ff0cffccfe9afe83fe93fed2fe37ffaeff2b009f00f7002b012e01f500;
    inBuf[5635] = 256'h8600ebff39ff8dfefafd8cfd51fd4ffd86fdf6fd91fe3effe7ff7700e3003201;
    inBuf[5636] = 256'h600167014301ef007000e2ff61ff01ffc7fea4fe81fe57fe2cfe19fe3bfe96fe;
    inBuf[5637] = 256'h19ffafff39009c00d500e600d00096003b00c6ff4dffe2fe90fe63fe56fe63fe;
    inBuf[5638] = 256'h8bfecefe24ff86ffe7ff3200620079008000810073004800feff94ff1cffbbfe;
    inBuf[5639] = 256'h87fe83fea6fedbfe18ff5effb0ff09005c00880072002000aeff44ff09ff06ff;
    inBuf[5640] = 256'h29ff5aff83ffa0ffc1ffeeff1a0035002500e4ff86ff28ffe3fec7feccfee6fe;
    inBuf[5641] = 256'h19ff6affdcff6a00f10041014001ec005e00c4ff3effd9fe90fe52fe20fe11fe;
    inBuf[5642] = 256'h38fe98fe23ffb7ff32008400b200cf00ea00ff00fd00d7008d002d00d1ff8cff;
    inBuf[5643] = 256'h61ff4bff3bff29ff1cff1aff26ff39ff47ff49ff43ff3cff41ff5cff89ffbeff;
    inBuf[5644] = 256'hf6ff2f0068009c00be00c200a20067002500fbfff2ffffff0a00f8ffbfff6eff;
    inBuf[5645] = 256'h21fff3feeffe07ff29ff46ff5fff81ffc0ff1e008d00f9004d01790176014401;
    inBuf[5646] = 256'hed007900f1ff6afffbfeb2fe91fe96febcfe00ff5cffc7ff35009500d000da00;
    inBuf[5647] = 256'hc1009a0076005d004e0044003c003a0049006a008b00950079003800ecffb4ff;
    inBuf[5648] = 256'ha3ffb1ffc4ffc4ffabff88ff75ff8affc6ff150060009d00ce00f9001c012d01;
    inBuf[5649] = 256'h2001f000a9006c00500056006d0077005f002a00edffbfffb0ffb7ffbfffbcff;
    inBuf[5650] = 256'hadffa3ffb4ffe7ff35008f00e2001e0145015b0163015c0145012201fc00d200;
    inBuf[5651] = 256'ha600770043000900d5ffb4ffb3ffd3ff06003b006e009800bd00e4000d012e01;
    inBuf[5652] = 256'h420141012f011501f400c50085002c00c4ff6cff3fff4dff9aff0d008700f000;
    inBuf[5653] = 256'h41018501cd011702590283027d023c02cb013e01a8001c00a2ff48ff19ff14ff;
    inBuf[5654] = 256'h39ff84ffe5ff5100c8004401bb011d024f024402ff0195012501d00095006800;
    inBuf[5655] = 256'h41001c000c002e008a000f019c0103022a021802e10199014601db005300c4ff;
    inBuf[5656] = 256'h50ff23ff5affe5ff99004901ce0123025c028202970291026002060298012501;
    inBuf[5657] = 256'hbc0066001c00e0ffc3ffd3ff18008700fe005d019c01bf01d501ee010202fa01;
    inBuf[5658] = 256'hc8016a01fc00aa0089009c00d50013014301670184019c01ab019d016e012901;
    inBuf[5659] = 256'hdf00ab00a000b500da000b0144018901da012702560254021902bc0169013701;
    inBuf[5660] = 256'h28013101340124010f01050112012e013a011d01dd00900066007e00cf003001;
    inBuf[5661] = 256'h79018d01780163016c019d01e901290246024602360225021602f401ad014501;
    inBuf[5662] = 256'hca005b001600fbff000022005e00c10055010302a20205030703ae0224029501;
    inBuf[5663] = 256'h2101cf008a0046000c00f4ff1a00860015019801eb010102f101e001e001ee01;
    inBuf[5664] = 256'hf801e301b0017a015901520156014001fb008c001900d6ffe7ff4500ca004d01;
    inBuf[5665] = 256'ha901d901f001ff010d0215020602dc01a20162012d010701e300bc0096007700;
    inBuf[5666] = 256'h690073009100bb00e900150142017501a301c301cb01b00173011e01bd006000;
    inBuf[5667] = 256'h1800edffe5ff000035007b00d2003701aa0126029802e502f602bd024302a401;
    inBuf[5668] = 256'hfa005b00d3ff63ff0cffd7feccfef3fe49ffbfff4400cc004d01c50131028202;
    inBuf[5669] = 256'ha8029e025f02f5017101e2005500d5ff6bff28ff15ff2fff69ffb2fff5ff3100;
    inBuf[5670] = 256'h6e00b40009016501b001d801d501af018001570132010501bc004e00c6ff48ff;
    inBuf[5671] = 256'hf8feeefe23ff7affd6ff24006500ac0007016801b401c4018001f000380084ff;
    inBuf[5672] = 256'hf9fea6fe8afea3feeffe6cff1700d4007b01e401f601b7014301bc003d00d3ff;
    inBuf[5673] = 256'h7eff3eff1aff12ff25ff48ff6bff82ff94ffa8ffc6fff1ff1a00310038003700;
    inBuf[5674] = 256'h41005e0083009a0090005d001100c7ff8dff61ff37fffcfeb0fe69fe3dfe3dfe;
    inBuf[5675] = 256'h6bfeb5fe0dff6bffc7ff21007300a400a800830045000700d6ffabff73ff23ff;
    inBuf[5676] = 256'hbffe68fe46fe68fec1fe2fff82ffa4ff9eff81ff5eff39ff07ffc8fe8cfe71fe;
    inBuf[5677] = 256'h95fefefe88ff020044003900f0ff89ff16ffa1fe2bfeb3fd50fd22fd37fd8efd;
    inBuf[5678] = 256'h0bfe85feeafe3dff8bffdfff3700700073003a00d5ff67ff0affb9fe66fe01fe;
    inBuf[5679] = 256'h8afd23fdf7fc18fd7cfdfbfd60fe95fea2fea3feb7fee9fe1fff3cff2efff9fe;
    inBuf[5680] = 256'hb9fe8bfe75fe71fe6ffe5afe39fe22fe1dfe2afe36fe26fef5fdb4fd7dfd71fd;
    inBuf[5681] = 256'h99fddffd28fe60fe77fe7bfe7afe6ffe57fe2ffefbfdd5fdd4fdfefd4bfe9efe;
    inBuf[5682] = 256'hd2fedffed3feb8fe9bfe74fe34fed8fd6efd0dfdd4fccdfce3fcfcfc09fd08fd;
    inBuf[5683] = 256'h13fd3ffd8cfdf4fd61febefe07ff3eff5eff60ff3affe6fe75fefffd93fd38fd;
    inBuf[5684] = 256'he4fc83fc1cfcc6fb9afbb9fb27fccbfc87fd3dfed9fe5bffc1ff03001a00fbff;
    inBuf[5685] = 256'h99ff04ff52fe9afdf8fc7efc2cfc01fcf4fbfafb1afc59fcb2fc21fd92fde9fd;
    inBuf[5686] = 256'h1dfe2dfe26fe23fe2efe3dfe46fe44fe3dfe40fe54fe6efe7bfe61fe12fea5fd;
    inBuf[5687] = 256'h3afde4fca9fc81fc61fc54fc6afcaffc21fd9ffdfcfd2cfe3bfe4afe7dfecffe;
    inBuf[5688] = 256'h12ff1affd0fe46feb6fd56fd35fd43fd51fd3efd13fdeffcedfc16fd4ffd6afd;
    inBuf[5689] = 256'h56fd21fdf4fc00fd59fde7fd7ffef3fe29ff29ff06ffd1fe97fe4ffeeefd82fd;
    inBuf[5690] = 256'h1efdd5fcbefcdafc15fd58fd8dfdaffdc8fde1fd00fe2afe56fe78fe91fea5fe;
    inBuf[5691] = 256'hb3fec2fec9feb9fe8efe4afefafdb2fd79fd4efd2cfd05fdd6fcb7fcc3fc09fd;
    inBuf[5692] = 256'h8efd38fedafe50ff89ff8cff73ff55ff35ff07ffb6fe40fec1fd5cfd2cfd41fd;
    inBuf[5693] = 256'h85fdcffd04fe24fe40fe6dfeaffef5fe29ff35ff1bfff2fecefeacfe86fe50fe;
    inBuf[5694] = 256'h0afed2fdc4fdecfd3cfe91fec7fed7fed3fed5feebfe03fffcfec9fe75fe25fe;
    inBuf[5695] = 256'h0dfe42fea7fe0dff4dff5bff52ff53ff6fff94ff95ff53ffd7fe51fefbfd01fe;
    inBuf[5696] = 256'h5dfee1fe58ffa0ffb6ffb1ffa7ff9cff83ff4afff6fea2fe6ffe73feb2fe14ff;
    inBuf[5697] = 256'h77ffc8ffffff17000f00e6ffa0ff49fffefed7fedbfef9fe16ff27ff38ff60ff;
    inBuf[5698] = 256'hb6ff3300a900e900e0009e004e001400ecffb0ff3cff97fefcfdbafd00febefe;
    inBuf[5699] = 256'hadff7a00ff0052019e01f001280203025701400021ff62fe33fe74fed3fe13ff;
    inBuf[5700] = 256'h36ff7aff1c000f01f4015602f001e500b3ffe2feacfef1fe60ffb5fff2ff4e00;
    inBuf[5701] = 256'hfc00ed01c9022403cf02ec01d900fbff7fff4bff2bff05ffedfe18ffa4ff7700;
    inBuf[5702] = 256'h4f01e1010d02ee01c001b101c201c901920111016d00deff99ffafffffff5900;
    inBuf[5703] = 256'h9c00c800f8004301a201fa011f02f0017d01fb009f008b00b600f30017011301;
    inBuf[5704] = 256'hff000f016301e801650295025302c0012801cc00ca00050135012e01fa00c900;
    inBuf[5705] = 256'hd40028019a01e601e1019101360114014101a70112024f025d025a0260026e02;
    inBuf[5706] = 256'h68022702a6010c018e005a007300b100ec0017013a017501db015402b602e502;
    inBuf[5707] = 256'hd702a80283027d029502b302b10284023502ce0166010d01c3008d0074007700;
    inBuf[5708] = 256'ha000f4006e010602ae024603af03d803b7036103f90290023402ea01a1015901;
    inBuf[5709] = 256'h210104010a01300161019101bd01e4010d023f026c028e02a802b702c302cd02;
    inBuf[5710] = 256'hc702aa028002520236023f0263029002b302b6029d0273023502e80193013b01;
    inBuf[5711] = 256'hf500dc00f6003c01a00106026802ca02250370039c0391034d03ea0286024002;
    inBuf[5712] = 256'h240219020502e001ab0186018f01c5010e0241023d020702cd01bd01f6016f02;
    inBuf[5713] = 256'he90224030803aa0253024a029c0219036f034d03ad02d8012f01f9003901a701;
    inBuf[5714] = 256'hf001f401c601ad01e6016802f5024a033c03e0027a023b0234024b0251023202;
    inBuf[5715] = 256'h0402e501ea01160249026e0287029b02b102c502b5026a02f3017a0134014701;
    inBuf[5716] = 256'ha50120028902bc02c102bf02c902e002f302e2029f023c02d9019b019d01d101;
    inBuf[5717] = 256'h16024c02560236020b02f201fd0129024e0245020a02b2016c016b01b8013602;
    inBuf[5718] = 256'hb402040326033a0358037f038f034c03970292018700cfffa2fff1ff80000f01;
    inBuf[5719] = 256'h7d01dc015802ff02b30333043d04c203fd024102d001b901cb01bf017e012a01;
    inBuf[5720] = 256'h0d015d010102a602e7028d02c001f0007e008400d1000d010b01f2001a01c701;
    inBuf[5721] = 256'he6020904a9048804cd03f5027402620275024a02a401a400bbff49ff65ffd8ff;
    inBuf[5722] = 256'h4e009c00d7003801e701d202a4030f04fa038803f80286023a02fa01b1016001;
    inBuf[5723] = 256'h270129016901c90117022602e8017601f40089005300530072009800b300c500;
    inBuf[5724] = 256'hed004e01f901d802ab032c043604d3034003c40275022e02b201df00d3ffe6fe;
    inBuf[5725] = 256'h6ffe8ffe22ffd8ff79000601a801820287036504bc045f0463031402d100d6ff;
    inBuf[5726] = 256'h31ffddfeddfe46ff26005c019f029403ec039803ce02dc01fd004800b0ff26ff;
    inBuf[5727] = 256'hb8fe93fee3feb1ffc700cb016a02860250021e022f027c02c502ad020602f900;
    inBuf[5728] = 256'hecff42ff1eff52ff8fffa0ff91ffadff38002c013502e402ee0263029a01f600;
    inBuf[5729] = 256'ha3008c007c004f001700feff22007300b800c20091004f002e003f0057003700;
    inBuf[5730] = 256'hc5ff2fffd5fe13fff9ff3e016402ff02f5028102fc019f015d01f700350025ff;
    inBuf[5731] = 256'h1bfe86fda8fd67fe5cff1200530048004a00a0003c01c501d6014e016e00acff;
    inBuf[5732] = 256'h5cff7affb4ffaaff4fff06ff5bff8a002c025a034703d401b8ff0afe76fdc1fd;
    inBuf[5733] = 256'hf8fd3cfd8efbf9f9ecf921fcfbffc603d0058905d40353021f02f70276033802;
    inBuf[5734] = 256'h09ff32fba8f8aff8eefabafd4fff16fffffdabfd0fffa401b803b3034f01defd;
    inBuf[5735] = 256'h5cfb10fbb4fccbfed6ff6aff6dfe3efe84ff9f011903ce02ce0054fed5fce6fc;
    inBuf[5736] = 256'hd6fd49fe60fd72fbd9f9e3f9ccfb8afe8c00e700fcff1aff66ffe9007b02ac02;
    inBuf[5737] = 256'heb000cfebffb51fbc0fcb9fea0ffc7feeefcacfb30fc4ffe9b006b011c0080fd;
    inBuf[5738] = 256'h47fbbefae5fb89fd40fe88fd2bfc96fbb9fc3cffb701b702cc01ccff2bfed8fd;
    inBuf[5739] = 256'h94fe35ff9dfea6fc4cfaf3f861f92ffb20fd13fed1fd20fd15fd2dfee9ff3001;
    inBuf[5740] = 256'h3301f8ff4cfe22fdd6fcf7fcbdfcc2fb68fa95f906faaefbbcfd26ff60ffb2fe;
    inBuf[5741] = 256'heffdb9fd0efe50fed4fd85fc08fb47fac8fa3cfca9fd26fe7ffd53fca2fb0ffc;
    inBuf[5742] = 256'h5bfd9ffef4fe14fe8cfc52fb07fb99fb5ffc9afc1dfc63fb1efbb5fbedfc0bfe;
    inBuf[5743] = 256'h6ffe01fe37fdbbfce4fc67fdabfd3dfd24fcf4fa57fa85fa3afbe5fb13fcd0fb;
    inBuf[5744] = 256'h8efbb0fb49fcfbfc42fdf0fc4ffcd9fbf6fb94fc2cfd40fdb5fce4fb71fbc7fb;
    inBuf[5745] = 256'hbcfcc0fd3afee5fd0cfd39fcc1fba7fb90fb12fb27fa2ff9a2f8d8f8c5f905fb;
    inBuf[5746] = 256'h3dfc40fd12feddfe9eff1000f0ff21ffc3fd44fc0dfb45fae3f9baf9a0f9a4f9;
    inBuf[5747] = 256'he9f977fa3cfbf7fb5efc6efc55fc4bfc83fcf6fc56fd61fdf5fc2dfc66fbf8fa;
    inBuf[5748] = 256'h02fb74fb0cfc8efcf7fc58fdabfde3fdd7fd5dfd84fc7efb80fab7f930f9e1f8;
    inBuf[5749] = 256'he1f847f919fa4dfba3fcb5fd49fe5cfe1efedafdacfd78fd18fd77fcb3fb27fb;
    inBuf[5750] = 256'h19fb7ffb16fc71fc47fcb6fb1ffbd9fa0cfb84fbddfbe2fb9afb4efb5efbdefb;
    inBuf[5751] = 256'h91fc24fd5afd36fd09fd1cfd82fd0cfe5bfe20fe63fd64fc77fbe4faaefaaefa;
    inBuf[5752] = 256'hc6faecfa30fbb7fb81fc63fd23fe84fe69fee9fd28fd58fcb1fb56fb52fbacfb;
    inBuf[5753] = 256'h50fc1afde6fd8efef4fe12ffdffe5bfe9bfdbdfcedfb60fb2ffb4dfba2fb0bfc;
    inBuf[5754] = 256'h71fce8fc88fd54fe26ffb2ffb8ff2fff46fe56fdb7fc7dfc7bfc73fc41fc05fc;
    inBuf[5755] = 256'h12fca9fcc9fd21ff2900780002000fff15fe76fd3efd36fd23fdf1fcc3fce0fc;
    inBuf[5756] = 256'h72fd66fe64ff05001500a5fff7fe55feebfdabfd72fd2dfdeafcd0fc0bfda2fd;
    inBuf[5757] = 256'h75fe4dfffbff6c00a500ad008c004000c0ff12ff59febffd63fd50fd7bfdd2fd;
    inBuf[5758] = 256'h3efeb1fe2cffa6ff09003d003300ebff86ff2bfff8fef9fe25ff65ffabfff5ff;
    inBuf[5759] = 256'h4700a000e800ff00cf006100d8ff67ff33ff3cff5eff6eff5fff4fff67ffc0ff;
    inBuf[5760] = 256'h4800c500f600c7005d000100f8ff4c00ca002f014a012401f600eb000f014701;
    inBuf[5761] = 256'h5b012e01e200b400ce002b018f01b3017201e3005000070022008300f6004c01;
    inBuf[5762] = 256'h7f01ad01e6012702590259021f02cf0193018b01bc01090253029302c302e402;
    inBuf[5763] = 256'hec02bd0243029301df0062004b008d00fa006001a901ee015b02fc02b7035404;
    inBuf[5764] = 256'h8c045004ce034003d902af02a002800245020202d901ee014702c9025403c203;
    inBuf[5765] = 256'h080423040804b30331038e02e801710140015801b7014d021603130428052706;
    inBuf[5766] = 256'hd406e40640061d05cc03a702f001a0018e019c01c5012a02f20208042405eb05;
    inBuf[5767] = 256'h0d068e05cb042c04f6032e0483049b045a04e2037e037503c10330048e04b504;
    inBuf[5768] = 256'hb804d2041f058905e105e4058405ef045104d20391037c038003ae030b049004;
    inBuf[5769] = 256'h2d05b105f6050206eb05d705de05e405c20577050805a2048304ac04f6043205;
    inBuf[5770] = 256'h33050705f2042205a8057106290784077207f8063d067c05c304180495034b03;
    inBuf[5771] = 256'h5203c603930490059706700701085708660824089707bd06b705ce042d04f803;
    inBuf[5772] = 256'h3a04ba044305ca053d06a0060507490751072407c60658060d06e405c0059005;
    inBuf[5773] = 256'h4a0515052f05a1055b062a07b007cd07b30791078b07a5079707200747063c05;
    inBuf[5774] = 256'h670429047f042a05d805390657067806c0063d07d6072e080f089107de063a06;
    inBuf[5775] = 256'he105c805d405ef05fd050a063e069a061807a7070f0832080d089407e4062e06;
    inBuf[5776] = 256'h8005fa04c404d6043005d30590064007cc070f080008bc074907c2064906e005;
    inBuf[5777] = 256'h9d059c05d1053106ab060b0738073c071d07f706e106be067e062506ba056505;
    inBuf[5778] = 256'h56057d05bb05f3050106fe05290694062e07c407ff07c007340792061b06e705;
    inBuf[5779] = 256'hc10579050f05aa049c0421050d060607a907ac0726077106cb055305fa048c04;
    inBuf[5780] = 256'h0904b303c7036f049805d306b5070a08cf074507b6062f06a5050b055b04c103;
    inBuf[5781] = 256'h7f03a7032c04de047005bf05d705c505a5058e0568052a05e804a90479046104;
    inBuf[5782] = 256'h49042204f003c603d7034304ec04a5053b066a0622069505e0041a045903a302;
    inBuf[5783] = 256'h0202a101a901360236035c045605e605ed058e0509057604dd0341039102e201;
    inBuf[5784] = 256'h790183010b02ef02d8037404a40470040b04b303790350032603da026d02fe01;
    inBuf[5785] = 256'ha3016f017301a401f5015802b202f10210030603dc02a6025e02fe018d011001;
    inBuf[5786] = 256'ha5008000bf0061013d020703800397035503e1026702e7014a0186009effbefe;
    inBuf[5787] = 256'h29fe0dfe79fe57ff71008b017e022c0389038d032e03790290018f0099ffcffe;
    inBuf[5788] = 256'h38fecefd97fda7fd10fed8fee0fff800df0153023c02b301dd00e0ffe2fef9fd;
    inBuf[5789] = 256'h36fdb1fc87fcd1fc92fdabfee5ffff00be01ff01ba01fe00efffbbfe90fd98fc;
    inBuf[5790] = 256'heffba1fbb0fb10fcaefc7afd5efe30ffc4fff7ffb6ff0dff31fe64fdd7fc96fc;
    inBuf[5791] = 256'h93fcaefcbffcc2fccffcf4fc38fd91fdddfdf5fdcafd5afdbbfc10fc79fb18fb;
    inBuf[5792] = 256'h03fb34fb9ffb29fcabfc11fd55fd72fd6ffd4bfdf7fc79fce4fb51fbe0faa8fa;
    inBuf[5793] = 256'h95fa8ffa85fa78fa8ffaebfa7bfb13fc75fc68fcf8fb6bfbf9fac6fabefaa2fa;
    inBuf[5794] = 256'h5afa01facff9fbf980fafefa22fbcdfa27faa5f9a8f928facafa08fb93faa8f9;
    inBuf[5795] = 256'hd0f877f8d2f89ff947fa78fa44faf7f9f3f94dfaacfaadfa17fafff8e6f747f7;
    inBuf[5796] = 256'h3bf7a3f72ef886f8b0f8e2f833f9a8f912fa23facbf92cf973f8e6f797f75df7;
    inBuf[5797] = 256'h33f71ff722f767f7ecf76af8b9f8caf89df875f883f8a8f8b5f86ff8aff7b8f6;
    inBuf[5798] = 256'hf2f59cf5d9f575f607f76bf7aaf7d5f723f885f89bf838f863f75af6acf5b2f5;
    inBuf[5799] = 256'h46f613f796f76ff7d9f649f602f626f675f677f619f69cf555f5a9f58df67ef7;
    inBuf[5800] = 256'h0ff807f875f7d5f679f647f615f6a4f5d5f40ef4cdf33af44df59cf695f70ff8;
    inBuf[5801] = 256'h1af8d6f786f72bf78bf6b1f5caf40cf4d9f341f4ebf495f504f616f611f62ef6;
    inBuf[5802] = 256'h5af688f68ff642f6d5f57df54af553f577f577f566f564f57af5c9f52ef656f6;
    inBuf[5803] = 256'h3bf6eef587f559f57bf5aef5c7f59df525f5c1f4c3f430f5f4f5b9f60cf7e6f6;
    inBuf[5804] = 256'h72f6ebf5a4f5a5f5a2f57cf52bf5c4f4a2f4faf4aef58ff63af753f7f3f651f6;
    inBuf[5805] = 256'h99f51bf5ebf4e0f4f9f42bf55cf5a0f5fbf54ff6aaf606f746f769f752f7ddf6;
    inBuf[5806] = 256'h2ff67ef5f7f4e7f451f5ebf584f6e9f6fcf6f6f6fdf603f704f7dbf66df6f6f5;
    inBuf[5807] = 256'hbcf5dcf56ff634f7bbf7e1f7adf745f701f709f735f75ff75af714f7cff6c2f6;
    inBuf[5808] = 256'hecf645f795f799f76af73bf735f785f70cf875f895f863f8fef7c2f7def738f8;
    inBuf[5809] = 256'ha6f8e0f8b8f863f82bf83af8a6f83af995f98ef928f98bf811f8e5f7f6f737f8;
    inBuf[5810] = 256'h85f8c5f814f988f918fab3fa2cfb5bfb45fbf3fa7cfa0efab4f963f929f9fff8;
    inBuf[5811] = 256'hd9f8d0f8f1f83ef9c9f984fa45fbf1fb61fc7efc68fc34fcecfba7fb5afbf8fa;
    inBuf[5812] = 256'ha0fa74fa8cfaf6fa85fbf6fb30fc3afc36fc64fccdfc3bfd75fd47fdb1fc03fc;
    inBuf[5813] = 256'h92fb80fbc3fb22fc69fc98fccffc32fdd7fd90fe13ff37fffcfe8afe26feeffd;
    inBuf[5814] = 256'hd2fdb7fd84fd3ffd12fd22fd80fd1ffecafe55ffb7ffecfff9ffe9ffb9ff6fff;
    inBuf[5815] = 256'h26fff5fef9fe44ffbcff3a00a500ec00120127012e011a01dc006800d8ff5dff;
    inBuf[5816] = 256'h22ff4bffdbffa300710117027c02b102c902ca02b80289023202ce0186017501;
    inBuf[5817] = 256'hb1012b02b6022803680372036703610363036e036b0347030d03d602c102f002;
    inBuf[5818] = 256'h5f03f403a3044505b805fc050b06e10596052d05ad043a04e303b003bd030f04;
    inBuf[5819] = 256'h97044e051006b406290752073407f906a9064f060c06d605a1058d05a005e205;
    inBuf[5820] = 256'h6e062807db076a08ae089f086a082508e807d107c407ae07a907b107c407fc07;
    inBuf[5821] = 256'h3d0866087c0878086d088c08d20829098e09d609ec09f109e709d509d009bd09;
    inBuf[5822] = 256'h94097c0974098009b709f009090a140a0c0a090a3d0a8e0ad90a170b240b090b;
    inBuf[5823] = 256'hfe0a0a0b2e0b720b990b8b0b6b0b430b2e0b590ba20be60b1f0c1e0ced0bc70b;
    inBuf[5824] = 256'ha80b960bb30be20b0e0c4f0c8d0cc40c080d350d360d1e0dd20c600c080cd40b;
    inBuf[5825] = 256'hd30b200c870ce50c3d0d750d980dd20d040e1b0e1a0ed80d5f0dfa0cb70ca70c;
    inBuf[5826] = 256'hda0c0d0d1a0d200d190d210d760df00d5c0eac0eb70e8b0e740e7a0e9b0ed10e;
    inBuf[5827] = 256'hcc0e6b0ed80d290d960c6b0c890cc90c2e0d940dfc0d990e4e0ff00f61104d10;
    inBuf[5828] = 256'ha40fb20eaa0dcd0c600c400c500c9b0c080da30d8b0e810f4210b0108e10e40f;
    inBuf[5829] = 256'h0d0f2f0e620dc40c300cac0b770b9c0b2e0c360d580e4b0f031059105e104310;
    inBuf[5830] = 256'he80f380f4f0e260df60b280bd00aec0a770b290ce70cc50d9d0e530fd80fdb0f;
    inBuf[5831] = 256'h440f540e320d260c840b350b200b490b8b0be90b8e0c4e0d010e8e0eaf0e570e;
    inBuf[5832] = 256'hc00df90c2c0c960b2a0be50add0aeb0a050b480b8d0bc70b080c2c0c2c0c260c;
    inBuf[5833] = 256'h080cdf0bd30bc60bad0b960b630b150bd90aa60a7d0a670a3f0a0c0af309e509;
    inBuf[5834] = 256'hec091b0a3a0a320a1d0a000af6091d0a4d0a680a680a310ad8098f0950091a09;
    inBuf[5835] = 256'hef08ab085c08360835085a08a308d608da08be08800840081a08f407c607a107;
    inBuf[5836] = 256'h6d073c07320738073f0752075807500751074f0746073e071d07de0695063c06;
    inBuf[5837] = 256'hdb058905470516050105fd040d0536056c05af05f40517060c06d4056c05f604;
    inBuf[5838] = 256'h9a04570428040304d503a003750365037d03aa03c603c2039b0358031c03fb02;
    inBuf[5839] = 256'he702d502b5027c0245022202130215021a0212020502fc01fc010b0219020502;
    inBuf[5840] = 256'hcb016f01fa008b002c00ddffa4ff81ff78ff9affe3ff3d009500cd00d600bb00;
    inBuf[5841] = 256'h81002e00d5ff71ff01ff9efe5bfe3ffe4ffe72fe8afe84fe54fe09fec1fd88fd;
    inBuf[5842] = 256'h68fd67fd73fd85fda5fdc5fde1fdf0fdd7fd93fd3afdd8fc87fc5afc3efc26fc;
    inBuf[5843] = 256'h08fcd5fba1fb8bfb8afb9ffbc2fbd3fbcdfbbdfb97fb6cfb4afb1bfbdffaa3fa;
    inBuf[5844] = 256'h5cfa18faecf9d3f9d6f9fcf92cfa61fa91fa94fa6efa36fae6f996f958f910f9;
    inBuf[5845] = 256'hbff879f83ef828f847f876f89cf8a6f87af836f803f8e2f7ddf7edf7e7f7d1f7;
    inBuf[5846] = 256'hcef7e4f724f879f89bf86ef8eff729f761f6d1f572f54cf54ff553f56bf5b4f5;
    inBuf[5847] = 256'h21f6b5f653f7b0f7c1f78df70af767f6d0f53ef5c5f46df420f4f6f303f430f4;
    inBuf[5848] = 256'h8df410f584f5e3f526f62cf607f6c6f554f5c7f437f49ff324f3e3f2d0f2fbf2;
    inBuf[5849] = 256'h57f3aff306f45cf491f4b2f4b8f487f440f4faf3b4f392f38df370f33bf3f2f2;
    inBuf[5850] = 256'h8ef251f25ef295f2edf23bf347f332f31af3f9f2eef2ecf2bdf276f233f2fcf1;
    inBuf[5851] = 256'h03f24ef29ff2e8f216f315f317f32bf327f30cf3c8f23ef2a5f12ff1e2f0e1f0;
    inBuf[5852] = 256'h17f14bf186f1caf1fef142f295f2c9f2e9f2eff2c0f289f25af21af2edf1d2f1;
    inBuf[5853] = 256'ha5f17ef158f110f1d1f0adf09cf0cef045f1c8f158f2dbf21cf339f334f3edf2;
    inBuf[5854] = 256'h89f20ef265f1c8f05cf01bf030f097f016f1b0f14bf2b7f20ff34ef34bf32cf3;
    inBuf[5855] = 256'hf0f272f2e8f16cf1f1f0b1f0b1f0c4f0fff058f1a0f1f7f165f2c2f222f376f3;
    inBuf[5856] = 256'h86f36cf331f3c6f262f21bf2d8f1bef1c8f1c6f1d6f1f9f107f224f254f273f2;
    inBuf[5857] = 256'ha1f2daf2f7f21bf34bf367f38cf3b4f3b3f3a8f398f369f342f327f3f2f2baf2;
    inBuf[5858] = 256'h8af257f259f29af2f8f27bf3fef34bf47bf494f484f474f45ef425f4eef3c6f3;
    inBuf[5859] = 256'ha4f3bbf306f44df498f4d3f4e2f4eaf4ecf4d1f4b3f489f446f425f434f45cf4;
    inBuf[5860] = 256'hb3f41df564f5a7f5e8f511f647f67cf67af651f607f699f543f51af506f51ef5;
    inBuf[5861] = 256'h5af59df508f698f622f79ff7edf7dff795f72bf7aef659f635f623f62ef651f6;
    inBuf[5862] = 256'h7cf6cff647f7c7f751f8c3f8f3f8f9f8ddf89ef86ef85af845f832f81af8eef7;
    inBuf[5863] = 256'hccf7bef7c1f7ecf737f885f8e0f843f9a0f904fa5dfa89fa8dfa6afa23fae9f9;
    inBuf[5864] = 256'hd4f9d6f9ebf9fcf9f4f9e4f9d9f9ddf90cfa5afaa5fae5fa0ffb1ffb38fb61fb;
    inBuf[5865] = 256'h8efbc4fbeffbfafbfcfbfffb02fc14fc2bfc32fc31fc2bfc23fc2cfc44fc5cfc;
    inBuf[5866] = 256'h78fc95fcb2fce8fc37fd87fdcefdfcfd09fe0dfe1bfe2ffe48fe55fe44fe1dfe;
    inBuf[5867] = 256'hf3fdd9fde6fd15fe4ffe8efed0fe18ff73ffd7ff2c005f00660043000c00d6ff;
    inBuf[5868] = 256'haeff96ff88ff86ff95ffbbff06007100e7005501ad01e401ff010402f301d301;
    inBuf[5869] = 256'ha9017b015f015b0167018e01c90103023a026e029702c002ed0213033a035e03;
    inBuf[5870] = 256'h730384039203a203c203ed030b0416040504d603a1037f038203bc031d048704;
    inBuf[5871] = 256'hee043b0560057505800586059605ac05bb05cd05d605d305d805de05dc05e405;
    inBuf[5872] = 256'heb05ea05f805110637067806bb06ef06270752076e079a07c907e9070208fb07;
    inBuf[5873] = 256'hd807bf07b207b007cf07ec07f107f907fa07fd0728086708a808f90834095209;
    inBuf[5874] = 256'h790994099b09b009b809a5099e098d0968095909540956098509c909070a510a;
    inBuf[5875] = 256'h890a9f0abd0ad70adf0aee0aea0ac70ab50ab10ab90ae40a0b0b150b200b230b;
    inBuf[5876] = 256'h260b550b900bb60bd90bdc0bc40bc90be10bfb0b280c400c350c2d0c220c160c;
    inBuf[5877] = 256'h220c1f0c000cf40bee0bf30b270c690ca20cea0c210d440d7a0d9e0d940d760d;
    inBuf[5878] = 256'h2e0dc50c7b0c500c450c760cb60cea0c2c0d5b0d6d0d870d8e0d7e0d840d910d;
    inBuf[5879] = 256'ha50dde0d100e1b0e160eea0d9b0d620d360d110d160d210d290d560d900dc60d;
    inBuf[5880] = 256'h110e480e530e520e380e0e0e010efc0df70d0f0e230e260e320e240ef60dc90d;
    inBuf[5881] = 256'h8c0d4c0d3d0d470d600da50dea0d1f0e640e960eaa0ec30ec30ea20e830e4d0e;
    inBuf[5882] = 256'h030ecc0d8e0d4d0d3a0d3b0d480d7c0daf0dd10d020e210e2a0e430e510e480e;
    inBuf[5883] = 256'h4a0e380e0d0eeb0db60d6e0d420d220d0c0d250d4a0d6a0d9f0dc40dd30ded0d;
    inBuf[5884] = 256'hf20ddc0dcc0daa0d750d570d360d110d090d000df30c030d0c0d010d000dee0c;
    inBuf[5885] = 256'hd00cd60ced0c0f0d4a0d6e0d6b0d5e0d350dfa0ccd0c940c510c260cff0be50b;
    inBuf[5886] = 256'hf80b0d0c170c290c230c120c220c380c500c7a0c8a0c7f0c7e0c670c3d0c1f0c;
    inBuf[5887] = 256'he90b9a0b5b0b1e0bec0ae40ae30ae80a0e0b340b540b870ba20b910b760b450b;
    inBuf[5888] = 256'h0b0bef0adb0ac60abd0a9e0a700a590a450a340a3d0a3f0a310a260a0b0ae709;
    inBuf[5889] = 256'hd709c409b109b909c609d409ec09ec09cf09ac0971092f090809e608c508b308;
    inBuf[5890] = 256'h94087208670863086d089408b208c008ce08c408aa08990875083808f1079307;
    inBuf[5891] = 256'h3407f906d406ca06e70602071007260738074b076d077c0768074107fa06a506;
    inBuf[5892] = 256'h650633060f060106ec05c6059f05700540052e052e053e05650589059d05a905;
    inBuf[5893] = 256'ha10584055f052f05f404b70477043e041904fa03e203d003b50395037b036303;
    inBuf[5894] = 256'h56035c0368037f03a603cd03ea03ed03c2036e03fc027802fc019b0154012e01;
    inBuf[5895] = 256'h30014e018e01e30133026c027f0266023102e60185012101bf005c000b00dcff;
    inBuf[5896] = 256'hcfffedff280067009f00c000bb0096005400fbffa3ff56ff18ffeffed5febffe;
    inBuf[5897] = 256'hb3feadfeacfeb8feccfedafedefecbfe9ffe64fe1afec5fd76fd37fd14fd13fd;
    inBuf[5898] = 256'h2cfd5efd99fdbefdccfdc2fd90fd44fdf2fc92fc31fce0fb9afb6dfb67fb7cfb;
    inBuf[5899] = 256'habfbeefb25fc44fc49fc20fcd7fb8bfb42fb09fbe7fac8faaffa9efa89fa78fa;
    inBuf[5900] = 256'h72fa6afa65fa61fa4bfa2cfa10fae7f9c0f9a0f97af95df953f94cf94ff95ff9;
    inBuf[5901] = 256'h69f975f982f97af964f93cf9f4f89ef84df8fcf7cbf7c1f7c5f7dcf701f81df8;
    inBuf[5902] = 256'h3ff868f87bf880f873f83bf8eef79ef746f701f7d5f6abf693f695f69ff6c6f6;
    inBuf[5903] = 256'h0af749f77ff7a2f792f76af739f7f0f6acf677f639f603f6ddf5b3f59df5a4f5;
    inBuf[5904] = 256'hadf5c9f5fcf528f657f687f697f68cf66af61ff6cef58ff557f540f54bf557f5;
    inBuf[5905] = 256'h6ef58cf593f598f59df587f56bf553f52bf50ef504f5f2f4eef4fdf401f511f5;
    inBuf[5906] = 256'h34f546f550f54ff528f5fcf4def4c0f4c1f4def4ecf4f4f4f8f4e1f4ccf4c6f4;
    inBuf[5907] = 256'hb3f4a8f4aaf49ef49cf4aaf4acf4b7f4ccf4c8f4c8f4d3f4c8f4c0f4c1f4a7f4;
    inBuf[5908] = 256'h8ff48bf483f48ef4a7f4a7f4a8f4aff4a0f4a4f4c4f4d0f4d9f4e1f4c6f4a5f4;
    inBuf[5909] = 256'h96f480f478f480f477f479f491f49ff4bcf4e9f4faf405f515f510f510f51cf5;
    inBuf[5910] = 256'h0ff501f5f3f4caf4abf4a1f48af486f49af4a5f4c2f4f4f413f531f547f539f5;
    inBuf[5911] = 256'h31f539f531f53af554f550f549f54df541f543f556f54ff544f539f512f5f3f4;
    inBuf[5912] = 256'hedf4e7f401f53bf56af5a5f5ebf511f62af63bf627f607f6e1f59ef561f535f5;
    inBuf[5913] = 256'h06f5f9f416f53bf57af5cff515f65df6a2f6c0f6caf6bdf678f621f6cdf573f5;
    inBuf[5914] = 256'h3ef53ef557f595f5eef53df68df6d8f609f72ff73ef71af7e1f69bf63df6f7f5;
    inBuf[5915] = 256'hddf5d8f5f6f530f663f69df6daf605f72ef74cf748f736f719f7e6f6c2f6b5f6;
    inBuf[5916] = 256'hadf6c2f6ecf611f745f77ff7a5f7c2f7d1f7bcf79bf771f735f709f7f2f6e0f6;
    inBuf[5917] = 256'hecf611f73af779f7c8f70bf84ff88af89ff89ef88af855f81bf8e7f7b0f799f7;
    inBuf[5918] = 256'haaf7ccf70df85cf890f8b4f8c7f8b7f8a4f89cf888f876f86bf857f858f881f8;
    inBuf[5919] = 256'hbbf808f959f98af9a1f9a9f99cf98df980f963f944f928f909f904f91bf937f9;
    inBuf[5920] = 256'h5af982f99ef9c0f9eef917fa3cfa57fa59fa52fa49fa39fa34fa38fa32fa36fa;
    inBuf[5921] = 256'h49fa63fa91facbfaf8fa1efb3bfb43fb44fb3ffb26fb08fbe6fabffaabfaadfa;
    inBuf[5922] = 256'hb7fad7fa09fb3cfb7cfbc8fb0efc50fc87fca3fcaafca2fc8cfc75fc5bfc38fc;
    inBuf[5923] = 256'h20fc10fc00fc00fc14fc2afc4afc72fc96fcc1fcf1fc1cfd4efd82fda5fdbcfd;
    inBuf[5924] = 256'hc6fdb9fda5fd97fd8cfd8cfd98fda1fdacfdbdfdd2fdf2fd18fe3afe56fe6afe;
    inBuf[5925] = 256'h77fe84fe8ffe92fe91fe8afe7cfe78fe8cfeb9fef6fe33ff65ff8dffa8ffbdff;
    inBuf[5926] = 256'hd2ffdfffddffcbffacff89ff72ff70ff86ffafffdcff0800320054006b007b00;
    inBuf[5927] = 256'h81007d007e0087009900b600d900ff0022013e01580172018101870185017a01;
    inBuf[5928] = 256'h6a0160015e0164016b016e0174017f019501bc01ef01250258027e029502a802;
    inBuf[5929] = 256'hb902c602ce02cc02c102b402a702a302b302c802d702e602f102f50202031503;
    inBuf[5930] = 256'h2803400354035e036e0385039f03c503f003130435044804430434041604eb03;
    inBuf[5931] = 256'hca03b503aa03b703d503fa0331046f04a804e00409051b0524051f050905f604;
    inBuf[5932] = 256'he204c604b204a1049604a604c604ec0428056b059f05ce05ee05f305e905d205;
    inBuf[5933] = 256'hac058c056f0552054805500562058e05c905ff053706660682069b06ab06a906;
    inBuf[5934] = 256'ha40696067e06730670066e06740676066e0671067e069406be06e70602071e07;
    inBuf[5935] = 256'h32073a074d0761076907710772076b077107750774077f07870788079907ab07;
    inBuf[5936] = 256'hb207c307d107d607ec070a08230840084e084b084f084f084f0862086c086508;
    inBuf[5937] = 256'h660860085708690881089708c008e508fe08220939093a09400937091a091109;
    inBuf[5938] = 256'h0b09020915092c093a0954096509650972097a0979099009a809b209cd09e109;
    inBuf[5939] = 256'he509f609040a070a170a200a1f0a320a440a480a5a0a670a600a610a5a0a420a;
    inBuf[5940] = 256'h380a2c0a1a0a210a350a500a830ab60ae10a1b0b490b620b7d0b7c0b5a0b390b;
    inBuf[5941] = 256'h110beb0ae80aee0af40a0d0b1d0b220b3a0b500b5d0b720b730b600b600b620b;
    inBuf[5942] = 256'h6c0b950bb40bc10bdc0be80be70bfe0b0e0c090c0f0c060cf00bf60b010c070c;
    inBuf[5943] = 256'h230c2c0c1a0c170c080ce70bdd0bd60bc60bce0bdb0bea0b180c470c6c0ca60c;
    inBuf[5944] = 256'hd40cec0c0a0d100df50cdd0cb20c740c4a0c1f0cec0bd80bc80bbb0bd50bfc0b;
    inBuf[5945] = 256'h230c640c950ca70cbb0cbd0cb00cbb0cc50cc50cd10cc90ca80c950c790c560c;
    inBuf[5946] = 256'h4e0c3d0c1b0c0d0cfa0be60bf70b0b0c150c2d0c330c260c280c230c180c250c;
    inBuf[5947] = 256'h260c190c240c2b0c2b0c440c520c4b0c4d0c370c080ce60bb60b790b570b330b;
    inBuf[5948] = 256'h0c0b070b060b010b1a0b350b480b700b8e0b9b0bb30bb90baa0ba30b890b560b;
    inBuf[5949] = 256'h2a0bf40ab70a940a780a5a0a4f0a410a2a0a260a230a1c0a250a240a160a160a;
    inBuf[5950] = 256'h120a080a130a1d0a1f0a2b0a2f0a220a140af209bc0986094209f908c4089808;
    inBuf[5951] = 256'h700860085f086808820896089d089f088d086d0854083e08290822081b081108;
    inBuf[5952] = 256'h0d080808fe07f307d4079f0765071e07d306970665063b0621060d0601060506;
    inBuf[5953] = 256'h0f0620063f065b066c067406680649062006e605a1055e051705d1049c047504;
    inBuf[5954] = 256'h5d04580457045704580450043f042d041004e903c1039403670346032b031903;
    inBuf[5955] = 256'h0f030403fb02fa02f602eb02da02ba0287024a020502bd0175012c01eb00be00;
    inBuf[5956] = 256'ha500a100af00c800e400f90003010001ef00cd009c005a001100ceff93ff61ff;
    inBuf[5957] = 256'h3eff24ff0efffcfeeafed4febefe9ffe77fe4dfe20fef3fdcffdaefd93fd84fd;
    inBuf[5958] = 256'h7afd73fd70fd64fd4dfd34fd15fdf4fcdafcb7fc8bfc5bfc1cfcd8fb9ffb6efb;
    inBuf[5959] = 256'h44fb26fb0bfbf8faf6faf6fafefa11fb13fb00fbdafa95fa43faf9f9b3f97df9;
    inBuf[5960] = 256'h61f94cf946f952f95af962f96df963f944f913f9c2f869f81cf8d4f7a1f78bf7;
    inBuf[5961] = 256'h7af77bf78df796f7a5f7b9f7b1f798f76ff724f7d4f691f648f614f600f6f2f5;
    inBuf[5962] = 256'hf9f514f620f628f632f618f6f3f5cdf58cf543f501f5b1f472f455f43ff445f4;
    inBuf[5963] = 256'h67f478f486f497f48ef486f483f45df428f4f4f3a6f362f343f328f322f330f3;
    inBuf[5964] = 256'h27f31ef323f312f305f304f3e4f2b9f293f255f227f215f2faf1f0f1fff1f9f1;
    inBuf[5965] = 256'hf9f10df208f207f212f2fef1e7f1d9f1b1f18ef17af14ff12ef126f10af1f7f0;
    inBuf[5966] = 256'hf9f0e1f0d1f0d3f0bbf0a9f0a8f090f083f089f07cf07ff09df0a4f0b1f0cbf0;
    inBuf[5967] = 256'hbff0aef0a7f07ff05bf046f015f0e8efcfefa6ef97efaeefbbefd5effbeffeef;
    inBuf[5968] = 256'h01f013f00ef014f028f01ef017f01af003f0fcef0cf0ffeff2efecefc8efaeef;
    inBuf[5969] = 256'haaef95ef8fef9aef91ef9aefb8efbeefd0efeeefebefebeff8eff1effcef19f0;
    inBuf[5970] = 256'h1cf029f043f041f043f04cf036f028f023f000f0ebefe7efd0efceefe7eff1ef;
    inBuf[5971] = 256'h11f043f05bf076f09af0a2f0b8f0daf0def0e5f0f0f0dff0ddf0eff0ebf0f4f0;
    inBuf[5972] = 256'h0af1fff0f6f0f7f0e1f0d9f0e5f0ddf0e4f002f10ef128f153f169f18ff1c9f1;
    inBuf[5973] = 256'he9f10bf233f239f23cf246f239f236f243f235f22af22af215f20ef21ef21ef2;
    inBuf[5974] = 256'h29f246f250f266f28ff2acf2d7f214f33bf366f397f3acf3bff3d7f3d4f3d7f3;
    inBuf[5975] = 256'he5f3dbf3d0f3cdf3b7f3adf3b4f3acf3b1f3c3f3c6f3d9f304f42af461f4a5f4;
    inBuf[5976] = 256'hcef4f3f419f526f538f550f555f55ef56cf569f575f58ff59af5aef5c8f5c8f5;
    inBuf[5977] = 256'hc6f5c6f5b4f5abf5aff5adf5c1f5ebf512f645f681f6aef6e4f61df73ef75cf7;
    inBuf[5978] = 256'h76f776f775f77af776f77af784f782f787f791f792f7a2f7c0f7d2f7e7f701f8;
    inBuf[5979] = 256'h11f82bf855f87ef8b0f8e5f809f927f941f94bf95af96ef979f984f993f998f9;
    inBuf[5980] = 256'ha2f9b7f9c7f9d9f9edf9f7f9faf9faf9f5f9fef916fa30fa53fa83fab1fae1fa;
    inBuf[5981] = 256'h15fb40fb66fb87fb9cfbaafbaefba3fb96fb8cfb81fb80fb8dfb9ffbb7fbd2fb;
    inBuf[5982] = 256'he6fbfdfb1bfc3afc5cfc7bfc8dfc98fca1fca8fcbafcd6fcf1fc10fd30fd49fd;
    inBuf[5983] = 256'h65fd83fd99fda8fdadfd9ffd91fd87fd82fd89fd99fdaafdcafdf6fd21fe52fe;
    inBuf[5984] = 256'h84fea6febffeccfecafec8fec8fec4fec5fecffedcfefdfe31ff68ffa1ffd6ff;
    inBuf[5985] = 256'hf9ff0f001d0019000b00faffe4ffd5ffd4ffe2ff090045008600c50003013701;
    inBuf[5986] = 256'h5e01790183017c016d015b014d014c015e018101af01df010902310255026b02;
    inBuf[5987] = 256'h77027d0273026502620268027b029f02c602ef021a033d035b0381039e03b203;
    inBuf[5988] = 256'hc603cd03cf03e203f903120436044e045304590455044a044c044d044f046204;
    inBuf[5989] = 256'h75048904b804ee041f055d059405be05ec050a0616062d063e06480663067b06;
    inBuf[5990] = 256'h87069e06ab06ae06c106d506e40606072307340757077d07a107d70708082b08;
    inBuf[5991] = 256'h5b088808ae08e808210952098e09c009e009090a280a350a460a4a0a3f0a420a;
    inBuf[5992] = 256'h440a440a5f0a830aa70ae60a250b5d0ba80bed0b220c620c970cbb0ceb0c0d0d;
    inBuf[5993] = 256'h210d470d630d700d8c0d9a0d950d9e0d9c0d8b0d8f0d8e0d880d9e0db60dce0d;
    inBuf[5994] = 256'h070e3e0e6d0eb80efc0e2c0f690f900f9a0fb20fbb0fb10fba0fb20f930f8a0f;
    inBuf[5995] = 256'h780f580f5b0f5a0f4a0f550f590f520f730f980fb50ff30f261042107910a710;
    inBuf[5996] = 256'hc310fb10261135115a116c1160116c11681146113a112311f910f710f210e210;
    inBuf[5997] = 256'hff1021113c118811d71117127b12d2120913531386139813bf13d313c713dd13;
    inBuf[5998] = 256'hec13ea1311142f143314551467145d1478148d149214c114ec1409155815aa15;
    inBuf[5999] = 256'hf4156e16de163117a117fc172f1875189f189f18b118a1186f1868185d184018;
    inBuf[6000] = 256'h591874188318ca1812194c19b519101a481a9e1ad71aed1a2d1b5c1b6c1baa1b;
    inBuf[6001] = 256'hdb1bef1b301c611c6e1c9d1cb01c971c9d1c861c4c1c431c311c081c201c401c;
    inBuf[6002] = 256'h561cae1c041d401da71df51d151e4f1e631e461e4a1e321ef41dea1ddb1db51d;
    inBuf[6003] = 256'hc81dd51dc61ddf1de41dc81dd71dcf1da71dae1da81d871d9a1da61d981db41d;
    inBuf[6004] = 256'hc01dad1dbf1dba1d931d891d5f1d0e1dd91c871c161cca1b6e1bfc1ab71a6f1a;
    inBuf[6005] = 256'h201a041ae319be19c619c019a619ad19981965194319f91889182818aa171217;
    inBuf[6006] = 256'h95160a167f151c15b1144114f2138e131913b9123d12af113411a3100a10910f;
    inBuf[6007] = 256'h140fa30e610e230eee0dd20d9e0d580d140da40c170c860bcc0af9092c095008;
    inBuf[6008] = 256'h7f07d2063006a4053a05d00473042a04d60383033503d2026702fc017e010801;
    inBuf[6009] = 256'ha4003b00e5ffa0ff57ff1cffebfeaefe72fe33fedbfd79fd0afd81fcf7fb6bfb;
    inBuf[6010] = 256'hdefa6cfa0dfabff997f981f976f989f99df9a8f9b4f99cf95ff917f9acf82ef8;
    inBuf[6011] = 256'hc2f74cf7ddf696f652f61cf60ef6fbf5e6f5e3f5bff584f54ef5f2f488f430f4;
    inBuf[6012] = 256'hc0f359f31df3d9f2a6f2a1f28df27df285f261f221f2def15bf1bcf024f067ef;
    inBuf[6013] = 256'hb2ee23ee82edffecb8ec65ec2dec2aec0bece4ebc9eb72eb01eb97eaf3e944e9;
    inBuf[6014] = 256'hace8f0e742e7c3e62fe6b6e571e50ce5a7e459e4cee331e3a2e2e1e126e193e0;
    inBuf[6015] = 256'he4df54df07dfaede7cde8dde87de8edeadde8bde57de25dea6dd1bdda1dcecdb;
    inBuf[6016] = 256'h45dbccda2edab3d978d924d9f5d8fdd8ddd8d3d8efd8d0d8c2d8dad8b9d8afd8;
    inBuf[6017] = 256'hd8d8d2d8e8d82ed942d96cd9c0d9d3d9e6d909dad9d9a4d97fd913d9bfd897d8;
    inBuf[6018] = 256'h3bd80ad81ad806d81ed873d89ad8dbd842d96dd9a6d9f7d906da28da67da68da;
    inBuf[6019] = 256'h83dac4dad2da04db5cdb75db9edbdddbd4dbd3dbdfdba1db6ddb4ddbeedaaada;
    inBuf[6020] = 256'h91da5ada57da88da9cdadeda4adb90dbf6db72dcb3dcfcdc43dd45dd4edd60dd;
    inBuf[6021] = 256'h49dd53dd74dd7eddb9dd12de5ededede72dff1df9ae04ae1e0e19fe262e30de4;
    inBuf[6022] = 256'hdee4abe55fe633e7f3e792e84de9f5e988ea45ebfdebb5eca4ed9ceea4efecf0;
    inBuf[6023] = 256'h3ef2abf354f5f8f6a5f875fa29fce2fdb5ff5a01f902a50415067707e408160a;
    inBuf[6024] = 256'h430b7d0c850d960ebf0fc710ec1136136b14c7154417a818321ad11b4e1df01e;
    inBuf[6025] = 256'ha3202d22ce237225e4266928e929372b8e2ccb2dc62ebe2f893004317931bc31;
    inBuf[6026] = 256'hb231a73179311f31e630ac306c30673071308630da302b316d31c831f031dd31;
    inBuf[6027] = 256'hbc31423179309d2f762e232de52b892a30291028e526ce25f8240d241d234a22;
    inBuf[6028] = 256'h3c210720d81e6a1de01b6f1ae1185e170916a71463134d121911e80fc00e4c0d;
    inBuf[6029] = 256'hb30b090a0e0802060f040b023900c1fe73fd7ffcf5fb8cfb5dfb65fb4ffb22fb;
    inBuf[6030] = 256'hd8fa31fa49f935f8d9f664f5f5f385f23af125f03bef96ee2ceee5edc8edbfed;
    inBuf[6031] = 256'hb4edb3edaded9eed9beda1edc2ed0aee62eed9ee7aef1cf0c7f083f11bf28af2;
    inBuf[6032] = 256'hd7f2e0f2b8f277f20cf2a5f15af115f108f141f194f126f2f1f2aef376f441f5;
    inBuf[6033] = 256'hbff512f641f60cf6a2f51df546f463f39ef2b6f1eff06ef0e2ef81ef6def47ef;
    inBuf[6034] = 256'h2cef36ef05efc2ee8dee0fee74ede9ec17ec37eb79ea82e98ae8c8e7dae6ede5;
    inBuf[6035] = 256'h2ce52fe428e342e217e1dedfcede8cdd4ddc48db1fda10d950d880d7d1d66bd6;
    inBuf[6036] = 256'he8d578d53ad5c4d441d4ced30dd337d272d173d07bcfaacebacdf5cc76ccfbcb;
    inBuf[6037] = 256'hc8cbe4cbf7cb3acca2ccdbcc2bcd86cd9bcdbbcddecdbbcdb6cdd1cdc2cdedcd;
    inBuf[6038] = 256'h56ceb1ce59cf47d02ad155d2b9d306d58ed640d8ced983db47ddd2de6fe0fde1;
    inBuf[6039] = 256'h37e37be4a2e55fe618e7b5e7e9e71ee846e819e8ffe7eee7a0e780e782e772e7;
    inBuf[6040] = 256'hace72be8a9e873e988ea89ebc3ec2fee5def98f0e1f1ccf296f34ef498f4b1f4;
    inBuf[6041] = 256'ha5f425f471f39ff26cf12ef008efb9ed8feca9ebcdea3cea02eacde9c7e9e0e9;
    inBuf[6042] = 256'hb4e968e9f9e821e821e712e6c2e478e35ee24fe18ae031e011e036e09ee015e1;
    inBuf[6043] = 256'h92e1fee149e276e272e24ae220e2e0e1a6e194e17ee177e195e196e17ee154e1;
    inBuf[6044] = 256'hd4e01fe053df50de6bddecdcc4dc63dd04df83e132e50eeaa2ef00f6d4fc6403;
    inBuf[6045] = 256'hb0095e0fc71333178d19781aa01a451a38195018e117a7174918d019ac1b3f1e;
    inBuf[6046] = 256'h4f2124241e27122a722cca2e233127338b356e388d3b7a3f0c44d1481f4e7653;
    inBuf[6047] = 256'h3858b85c7160e762ab647d653965c36416643463fe624b63ed63776569674e69;
    inBuf[6048] = 256'h726b1b6dd06df16d026de86a4f680d6562611b5e1b5bb7588c57245794571a59;
    inBuf[6049] = 256'hd85ab05cc45e16609f60bf60b95fc05d7a5b6a58eb54a851204e924a73471244;
    inBuf[6050] = 256'h9440493d5f39f5347a30512bcb259220501b6e169012600f330d690c670c480d;
    inBuf[6051] = 256'h230f0911eb12dd14ff15661676169015fa1361125f10370e960c0d0ba609d708;
    inBuf[6052] = 256'h0d08140743060e0546035e0109ff4cfccdf977f76cf552f409f48af444f6dcf8;
    inBuf[6053] = 256'h10fc160062049408e70cd41011140d177a19371be61c5d1e7c1ff0208f221324;
    inBuf[6054] = 256'h03262028ff29032ce12d2a2f48301631473159314e31063108315e31f5313833;
    inBuf[6055] = 256'h06353037f439f83cff3f3c433f46c848264b004d3c4e4f4f02504c5092509050;
    inBuf[6056] = 256'h2f50c64ffe4eb54d3c4c2b4a764782440f41483dbd394a362c33e730432f642e;
    inBuf[6057] = 256'h962e6b2fd730e332e334bb366b384a396639f53881375435d732c22f7e2c8229;
    inBuf[6058] = 256'h7226a2236d21501f681de41b301a531878162c149a110f0f530caa0952071605;
    inBuf[6059] = 256'h4c0317022001a400a0009400a300ce00a70063002800b6ff4cff18fff9fe01ff;
    inBuf[6060] = 256'h66ffe5ff74002a019a01b2016a0180000aff25fdd3fa57f8f1f5cdf33af25bf1;
    inBuf[6061] = 256'h43f115f2adf3e4f5aaf89ffb7dfe2c015303c804a005b50523053304d7024701;
    inBuf[6062] = 256'hdeff79fe31fd4efc87fbd4fa56faabf9c2f8bef74df68bf4baf29bf06dee90ec;
    inBuf[6063] = 256'hbeea36e94de893e72ae74ee760e75ce787e757e7dce665e67ce54fe446e3fae1;
    inBuf[6064] = 256'hace0b6df8ade52dd52dce1da25d95ed7ead402d2fcce50cb63c7b6c3e6bf78bc;
    inBuf[6065] = 256'he7b9a2b713b690b553b592b579b621b7acb73fb816b885b7dbb677b5e2b38fb2;
    inBuf[6066] = 256'hf1b093afd7ae1aaecead26ae59aecaae96afebaf32b096b060b026b034b0eaaf;
    inBuf[6067] = 256'hedaf83b0ffb0eab168b3bbb44eb623b876b9b0bac1bbffbb1bbc19bc55bbdcba;
    inBuf[6068] = 256'h98baf6b9efb951ba84ba2dbb2dbcb1bc47bde2bdc8bda1bd7ebdc5bc3abc09bc;
    inBuf[6069] = 256'ha6bbcfbb95bc41bd65bed7bfafc06fc1ecc147c128c09abef3bb12b93eb6fdb2;
    inBuf[6070] = 256'h4ab06aaeb8acf1ab24ac70ac49ad93ae5faf19b0adb052b095af95aed6ac15ab;
    inBuf[6071] = 256'h84a9c5a78aa6dca53da52fa57ca586a5b2a5bca526a56aa454a3a3a103a0559e;
    inBuf[6072] = 256'h789c249b209a3399d798a0983698f39767977c96b895e6945f94e89463965199;
    inBuf[6073] = 256'h6b9e55a549ae6fb9bcc5e9d287e018ed53f8e9018808750c150ebb0c65093905;
    inBuf[6074] = 256'h060001fb52f791f481f3aff424f717fb8e0041063f0c93122e187c1df422f527;
    inBuf[6075] = 256'h1c2d053335391b40f04702506d58d8605668216fd6745a78037a237abc783077;
    inBuf[6076] = 256'h9975e4733b737e73537425769d78f27a287dca7e2e7f697e557cf478d3742a70;
    inBuf[6077] = 256'h886bb167c5644563a06353656e68e26c83710776397adc7cdc7d6c7dc47a4e76;
    inBuf[6078] = 256'hc170c1690062445a3052624a56435e3cce35d82f9e2967236f1d0c17b710cd0a;
    inBuf[6079] = 256'heb04c3ffa4fb29f8faf51ff5d8f48ff509f745f88ef9bbfae3fa5efa4ef91af7;
    inBuf[6080] = 256'h41f428f175ed8de9c1e5cbe1dadd0bda0bd6e1d193cdf2c824c45bbfaeba69b6;
    inBuf[6081] = 256'heab26ab01faf47af0ab164b43cb95bbf67c611cee7d56ddd61e46bea40ef05f3;
    inBuf[6082] = 256'ha6f506f7b0f7d7f76cf70bf7f0f6dbf646f750f879f90bfb19fd08ff13016903;
    inBuf[6083] = 256'h8505a207150a7a0c080f1d1277153a19a11d6d22ac27642d3d333d395a3f0245;
    inBuf[6084] = 256'h724a7a4f94531657bd59525b1c5c0d5c0c5b6c5939576d545e51214ec24a8a47;
    inBuf[6085] = 256'h8344b541633f8e3d443ca13b843bfe3b1a3d8c3e5b40784268443346cb479848;
    inBuf[6086] = 256'hb5484448ca468144b541033ec7397535b530e72b7627f822a91ed81a10177c13;
    inBuf[6087] = 256'h53101f0d100a4a076904b3015bff0efd33fbf4f9edf877f8aaf8fff8b8f9e3fa;
    inBuf[6088] = 256'heafbf3fc0ffebffe27ff66ff23ff87febbfd7efcf8fa48f940f7fff49bf2f6ef;
    inBuf[6089] = 256'h2fed69eab0e732e50ee355e12fe0a8dfd5dfcce069e296e442e729ea21ed14f0;
    inBuf[6090] = 256'hc1f209f5ebf644f810f96ff96df926f9bef84df8f4f7b2f783f788f7acf7cef7;
    inBuf[6091] = 256'h04f82cf81bf8faf7b8f72af799f60df65bf5ccf476f430f444f4c6f478f592f6;
    inBuf[6092] = 256'h1ff8cff9c4fbfbfd15002402180491059e062f07ec06010676040a0205ff9cfb;
    inBuf[6093] = 256'hb4f7acf3c4efe8eb79e8ade550e39de1abe018e0fadf4ee09ae0eee054e161e1;
    inBuf[6094] = 256'h2fe1ebe041e05adf85de8bdd9bdc00dc7adb18db07dbfddafada17db03dbb8da;
    inBuf[6095] = 256'h41da5ad91ad897d6a3d47dd249d0decd94cb91c9a1c725c64ac5ccc4f7c4ebc5;
    inBuf[6096] = 256'h4ac747c9e9cbc5cefed181d5d8d82bdc68df25e29ae4bee63ce869e94eea9fea;
    inBuf[6097] = 256'hbeeab4ea32ea94e9d8e8a4e75ee606e545e38fe1f9df36dedadc0cdc6fdb78db;
    inBuf[6098] = 256'h40dc4addecde24e158e3bee545e84eea11ec8fed45ee98eeb1ee28ee70edbbec;
    inBuf[6099] = 256'ha7eba1eac0e981e83fe703e639e445e245e0c1dd3adbefd872d64ed4ccd277d1;
    inBuf[6100] = 256'hb9d0c4d004d1a8d1b9d296d367d441d59dd5a7d593d50dd541d471d373d25ad1;
    inBuf[6101] = 256'h4cd03ccf20cee3cc8dcb20ca68c895c6dac4f4c219c1a3bf43be11bd58bcbdbb;
    inBuf[6102] = 256'h36bbf2ba98ba32baedb99db9a9b97aba13bc17bff4c390ca64d375de15eb3bf9;
    inBuf[6103] = 256'h4a08ef16d22425318b3a0a4177442144ea408c3b0b34e32b3224191dd8171215;
    inBuf[6104] = 256'h4414f115ff193d1fbd25362d22340c3afb3ef242c646aa4a884e1a535258d75d;
    inBuf[6105] = 256'h0f64696a4770eb757a7a4d7dfa7ef67eec7cf5791f7675713b6db069da668865;
    inBuf[6106] = 256'h9065a066e3689e6b516ef070aa7248731473ac716f6f0c6d686a2968f2666e66;
    inBuf[6107] = 256'h0267ce68e26a3c6da76ff57021712770256d7b689e623d5b1053bc4a1f42f739;
    inBuf[6108] = 256'h9a32a92b95254e20291b7516fa11180d4e08a203befe6afacff6a7f3b6f1fbf0;
    inBuf[6109] = 256'he0f0d5f186f302f56df664f7fdf670f5bff270eefee8d5e2f7db00d569ce42c8;
    inBuf[6110] = 256'he9c27cbecebae4b784b55db364b16eaf61ad6aaba8a954a8cea753a827aa88ad;
    inBuf[6111] = 256'h68b2a2b806c030c89dd0c0d82ae060e6f0ead4ed0fef84eeafec1aeadce68be3;
    inBuf[6112] = 256'hc8e087de23ddf5dc92dd02df64e116e40ce77deadced37f1fbf4daf8f7fcc801;
    inBuf[6113] = 256'h01079d0cd5124419b11f0326c62bd830163528383a3a6a3b9a3b453bce3a273a;
    inBuf[6114] = 256'hc239ee396e3a563baf3c143e513f38407540ea3f893e573c8b39623630335730;
    inBuf[6115] = 256'h252ef22ce32cdb2dd72f94328c357b38f53a5d3c9a3c8b3be538fd342630762a;
    inBuf[6116] = 256'h8024b61e3019631477102a0d9f0ab008df063205860378013cffe3fc4ffaf1f7;
    inBuf[6117] = 256'hfaf554f467f343f39cf394f4fbf555f7a1f8a4f9eef997f995f8c2f667f4b0f1;
    inBuf[6118] = 256'hafeebcebf3e857e618e423e262e0e2de6dddeadb6fdadfd853d70bd60ed590d4;
    inBuf[6119] = 256'hd8d4d1d58ed71bda25dd85e00fe450e70bea13ec20ed3ced76ecd6eabae861e6;
    inBuf[6120] = 256'hefe3d0e131e011dfafdeefde84df83e0aee1a5e28ce345e496e4d8e423e560e5;
    inBuf[6121] = 256'h01e62be7aae8bdea59ed11f0e9f2b9f50ff8eff940fbc3fbbdfb49fb56fa59f9;
    inBuf[6122] = 256'h82f8abf732f721f714f734f771f747f7cbf602f68ef4a7f283f0feed86eb6ce9;
    inBuf[6123] = 256'h8fe74ee6e4e500e6bee620e8a7e943ebdbecf7ed99eecdee4fee50ed0bec63ea;
    inBuf[6124] = 256'ha8e818e796e55ee492e3eae274e233e2d9e16de1ede027e04bdf6ede6fdd9cdc;
    inBuf[6125] = 256'h13dca6db9adb00dc7ddc38dd32de00dfcedfade045e1dfe1ade264e350e498e5;
    inBuf[6126] = 256'hdbe652e804ea66eb9bec97edbded44ed4eec68ea00e86fe56ee289df1cdddada;
    inBuf[6127] = 256'h41d989d825d86dd872d97adab8db2bdd1adecbde63df51dff7de8fdea3dd9cdc;
    inBuf[6128] = 256'hc0db8eda60d966d808d7a2d55dd4acd2f2d05fcf7dcdc8cb76ca1ac92ec8dac7;
    inBuf[6129] = 256'h93c7afc738c88ac8e2c84ac92ac9c0c82fc80ec7aac540c493c2f6c093bf3ebe;
    inBuf[6130] = 256'h2fbd58bc88bbedba52ba85b9c8b8dcb798b64eb5d1b30fb26cb0c7ae1cadccab;
    inBuf[6131] = 256'hc3aa25aa55aa46ab4aadbab065b598bb82c39ccc01d781e21feeb3f9d404560e;
    inBuf[6132] = 256'h2f16251c501f3020261fdc1b6f17c012c40dab0936071306ff06240aa40eb314;
    inBuf[6133] = 256'hf41b3e23b12afd314338fc3d2e437647a44bdf4fe7537c587b5d6662a867bb6c;
    inBuf[6134] = 256'he9708d742377257824781177ed743172956ed96a8d6886678e673469df6b1e6f;
    inBuf[6135] = 256'h0d73d676157aec7caa7e517f547f5a7ecd7c467b7879d477bb768a7574749b73;
    inBuf[6136] = 256'h1972f76f486d50695464ab5ef357c550a6496942bd3bf135a430552cfe28f125;
    inBuf[6137] = 256'h7a236321ea1e771c021af716f41323110c0e5b0b37090e075d051f049002f600;
    inBuf[6138] = 256'h39ff98fc5df9a3f5eef0abeb2de63ee05bdaded4a8cf18cb54c71cc4a6c1ebbf;
    inBuf[6139] = 256'h87be93bd0cbd9fbc71bcabbc18bdd7bd23bfd2c0e8c298c5b0c8fbcb89cf0ed3;
    inBuf[6140] = 256'h2fd606d962dbe4dccadd25deb7ddefdc1ddc10db43da21da72da8cdbbbdda1e0;
    inBuf[6141] = 256'h63e41de94dee02f43bfa6900a906fb0cd4127118e91db62221275b2be92e1032;
    inBuf[6142] = 256'hfc343437f0384d3ade3ae93a823a5839d63738365434c332db31883151327734;
    inBuf[6143] = 256'hc737763c5442e148f04fe856235d6a622b6607682e6879660a638c5e2b595153;
    inBuf[6144] = 256'hb94d7c48e14357408b3d5d3be2398038ff3673356f330731912edf2b4f295927;
    inBuf[6145] = 256'hd52521257a255d26dd27f129c22b2f2d252ede2d692c072a5a26c821e41c9e17;
    inBuf[6146] = 256'h7912000e150a0307ef04710391023102c2014401a9009bff57fefefc78fb2dfa;
    inBuf[6147] = 256'h3bf981f84ff897f8fff8a5f956fa9efa93fa1afaf1f84af746f5eaf282f035ee;
    inBuf[6148] = 256'h1cec6dea1be915e858e7a5e6e4e504e5c7e349e2b1e0e8de47dd28dc7cdb89db;
    inBuf[6149] = 256'h93dc59dedbe00be467e7bfeae2ed53f005f2f1f2d5f2f6f18ef094ee7aec7eea;
    inBuf[6150] = 256'h82e8e3e6b9e5a8e4dee351e388e2afe1d2e091df44de24ddf8db2cdbfcda13db;
    inBuf[6151] = 256'hbedb1bdda8de80e09ee269e4f3e53ce7c9e7cde76ce75ae6fbe48be3c0e103e0;
    inBuf[6152] = 256'h89deecdc76db3ddabfd83bd7cad5f9d31ed273d0b0ce49cd83cc11cc61cc9acd;
    inBuf[6153] = 256'h39cf71d135d4d5d65dd9afdb2cddfadd27de54ddecdb33dafad7d2d502d44bd2;
    inBuf[6154] = 256'h25d1abd061d093d031d1a3d12ad2c7d2f9d224d36bd36cd39fd330d4afd484d5;
    inBuf[6155] = 256'hc3d6dfd725d991da84db4edcf0dcd9dc7ddc01dcebdac5d9c5d874d756d68cd5;
    inBuf[6156] = 256'h7dd49bd3fdd2fdd110d151d022cf17ce67cd70ccc8cbaccb71cb8ecb22cc67cc;
    inBuf[6157] = 256'hc0cc3ccd11cda1cc10ccb0ca04c953c717c5e9c217c127bfa5bdc4bce4bb72bb;
    inBuf[6158] = 256'h7dbb4abb2abb2abba4baeeb933b90cb8ddb6d9b5c4b4efb35cb3dab2a5b27fb2;
    inBuf[6159] = 256'h30b203b2adb1feb067b0b3afd1ae40aecfad72ad8badccad22aeceae79af46b0;
    inBuf[6160] = 256'h89b109b340b5afb827bd33c33acbaed4b9df35ecf8f8b505d511e81bc0231729;
    inBuf[6161] = 256'hf72afb29bb2610215c1ad3139f0d1d093907a507030b481150190723c02d0d38;
    inBuf[6162] = 256'he541d34ada51ad57795ca15f11628c641c67756a6a6e6072a8768d7a117d657e;
    inBuf[6163] = 256'he67d0f7be576aa717c6bbb65f060495dae5b135c225e0162f2664f6cef71e876;
    inBuf[6164] = 256'hc97ab67d1a7f1a7f527e887c347a0a78b1757a73c671cd6f926d326bc9676763;
    inBuf[6165] = 256'h595e16581951074aba42e83b26363031882d3e2b8e29a02823280e2792258d23;
    inBuf[6166] = 256'h3e20351cc817a812b60d6b098005a402f500c1ff3fff33ffa3fe93fdd7fbbcf8;
    inBuf[6167] = 256'h92f49eefbbe992e3b5dd39d8b5d377d049ce4acd53cdd0cd97ce60cfa5cf5bcf;
    inBuf[6168] = 256'h99ce4bcdc0cb65ca6cc92ac9f3c9c1cb84ce3bd27bd6d0da0fdfc2e278e555e7;
    inBuf[6169] = 256'h4de835e89de7e5e607e699e5f6e5d8e67de8f4eaaaed9cf0b6f36df6edf863fb;
    inBuf[6170] = 256'h7ffda9ff44022005a008050deb115d17341dcb220828b42c4930ef32b9348135;
    inBuf[6171] = 256'hd7351536443603378b38a43a8b3d1241a1441a481a4b094de74d934dec4b5449;
    inBuf[6172] = 256'h204699424d3f923cb03af339323a593b503d853fab419343a944d9444244aa42;
    inBuf[6173] = 256'h5a40b63db63abd371c359c326e30982e982c722a22282b25ae21db1d86191e15;
    inBuf[6174] = 256'h0a11490d550a78087c078f079508ff09bc0b800da60e2f0f070fcf0dd60b5d09;
    inBuf[6175] = 256'h590649037f00e7fdcffb46faf9f8f4f712f7e5f573f4b2f26bf0d9ed36eb95e8;
    inBuf[6176] = 256'h4ce699e496e373e31ee471e55fe78ee9adeba3ed23ef06f067f02ef078ef93ee;
    inBuf[6177] = 256'h86ed86ecd4eb57eb24eb4aeb78ebaaebe6ebd6eb96eb48ebb3ea1ceacee990e9;
    inBuf[6178] = 256'hace961ea4eeb94ec49eedeef5cf1d0f2b3f325f456f4e5f328f378f288f1b8f0;
    inBuf[6179] = 256'h63f01af018f094f0f3f044f1b5f1b8f161f1f3f01cf01eef3fee50edbbec83ec;
    inBuf[6180] = 256'h8aec02edbbed73ee19efa0ef8eef03ef1aee79ec6fea4be8dae581e38fe1bcdf;
    inBuf[6181] = 256'h43de45dd5bdc92dbebdafbd9e6d8c3d753d6e6d4b1d392d2ebd1e3d141d242d3;
    inBuf[6182] = 256'hd7d48bd66ad848daa2db8fdcf7dc8ddcabdb72dac2d821d7bad560d486d334d3;
    inBuf[6183] = 256'h06d33dd3bad306d465d4bad49fd488d487d45ad4a1d47ad588d649d8b5da2add;
    inBuf[6184] = 256'he6dface2b3e435e60be79be66de5a5e3ece011de68dba3d889d65bd58cd49ad4;
    inBuf[6185] = 256'h7fd568d69ed705d9c8d943da89da08da5cd9dcd81cd8c1d705d853d814d94ada;
    inBuf[6186] = 256'h29dbe6db6adcf3dbcdda1bd96dd65ad34bd00fcd4aca58c800c7a7c64bc760c8;
    inBuf[6187] = 256'hf6c9cbcb43cd6cce18cff8ce64ce70cd18ccdecae0c914c9c1c8b9c8ccc804c9;
    inBuf[6188] = 256'hf4c866c866c795c512c34cc023bd06ba9fb7d0b5f9b47fb5efb652b9a4bc10c0;
    inBuf[6189] = 256'h94c325c702ca89cc2dcf8fd16fd48dd89ddd35e4a8ec1af67300440b1a15831d;
    inBuf[6190] = 256'hea231b274727ae241b1fd21707103e0809028afee9fde6008107ce10751c6d29;
    inBuf[6191] = 256'h3a365342d74cdb54a15a285e7f5fa75f185f3b5efb5d4b5e175faa6046626463;
    inBuf[6192] = 256'h2564d6633762d35fa55c2a59ff55f7521451a3512e5479588c5e4f65426c0f73;
    inBuf[6193] = 256'h7678507cb67ee17e557dc87adf7667722a6eb0697565d361ed5dea59da55dd50;
    inBuf[6194] = 256'h554b97452d3fea387933a22e452bcf29a3291a2bf92d0c312a34c636a537cf36;
    inBuf[6195] = 256'h1d34fe2e2b282220fa16db0d5f0588fd32f779f2d0ee7fec2febfae9f1e8f4e7;
    inBuf[6196] = 256'h4ee65de45fe207e0f7dd6fdc42dbcbdaf5da52dbdedb3ddce4dbd5daedd801d6;
    inBuf[6197] = 256'h6cd283ce87ca02c75cc4cfc294c2b3c3f4c51ac9cfcca6d03cd45dd7e3d9b0db;
    inBuf[6198] = 256'hfcdc0bdeffde2be0d8e1f8e39ee6c8e90eed40f030f369f5dcf695f76bf7b4f6;
    inBuf[6199] = 256'hdbf5eff479f4fcf473f622f933fd3a0207085c0e8914461a541f3723fa25ba27;
    inBuf[6200] = 256'h582849280528a927bd27a728632a2b2dfd306c35403a173f5a43be46e0487249;
    inBuf[6201] = 256'h8f483a469442303e8139fb343f31a62e6e2dd42db22fd432f236663bb33f7043;
    inBuf[6202] = 256'hf8450c4799466644b540f33b4b3643305f2ad0240020241c15190217d3151115;
    inBuf[6203] = 256'hbc14ab1474143214e6135b13cd124b12a9111c119d10ef0f320f450ee90c3d0b;
    inBuf[6204] = 256'h3709b906f4030001d3fdbafabff7d2f430f2c9ef7bed76eba0e9dee779e66de5;
    inBuf[6205] = 256'hbbe4c1e47ce5e0e623e910ec52efd8f22ef6d4f8a9fa45fb60fa22f882f4a7ef;
    inBuf[6206] = 256'h1dea30e445de07d9c2d4aed11dd0f3cf04d145d355d6ded9c6ddaee166e5f8e8;
    inBuf[6207] = 256'h30ec02ef91f1b0f34cf56ff6dbf677f653f546f362f0deecc1e857e4ffdfe7db;
    inBuf[6208] = 256'h77d8ffd57dd41ed4edd49dd622d952dcbbdf4ae3dfe61bea13edd8ef2ef238f4;
    inBuf[6209] = 256'hfff53af7fbf730f87bf7edf583f301f0b4ebd6e673e11fdc49d710d300d062ce;
    inBuf[6210] = 256'h11ce43cfdfd157d58cd924de61e21de628e90cebeaebe9ebe3ea39e93be7e6e4;
    inBuf[6211] = 256'h9ce293e09edeeedc87db1ddad0d89bd73bd6e9d4bad388d2b4d16ed18bd159d2;
    inBuf[6212] = 256'hefd3f1d577d876db70de67e142e495e67ae8f4e9bbea16eb1deb9aeadde900e9;
    inBuf[6213] = 256'hc5e77ae632e5aae335e2eee0a3dfb9de48de1bde9adecddf4ee16ae309e68be8;
    inBuf[6214] = 256'h10eb77ed1aef1df086f0e3ef91eed4ec73eaece79de558e389e167e09fdf68df;
    inBuf[6215] = 256'hb7df0ae087e018e138e122e1dfe013e025df42de2add54dceddba3dbc8db67dc;
    inBuf[6216] = 256'hfedcb0dd75ded6deeedec7de18de17dde5db6ddaf8d8a0d75fd66dd5b3d41dd4;
    inBuf[6217] = 256'hd3d38fd334d3efd27ed2d8d14cd1b4d016d0cacfaecfd0cf5cd018d108d233d3;
    inBuf[6218] = 256'h4bd485d503d788d882da3edd8ee0f5e4a4ea30f1d6f85b01ce0903126e19ef1e;
    inBuf[6219] = 256'h7a22d1235e22c91ea21922139e0c1307f3027601030348079f0e661862234c2f;
    inBuf[6220] = 256'h163b6945454e20555c59bf5b875cbb5b7d5a2859bb57fc56b8568556c756f256;
    inBuf[6221] = 256'h85560f564d551c545b531a5376532555d157635b6c6044663c6c47727f77697b;
    inBuf[6222] = 256'h2c7e3a7f9c7ee17cd379df75b6711d6d74682f64c55f615b4957e1526c4e5a4a;
    inBuf[6223] = 256'h4446a34200400f3e423ddc3d3d3f6e4127446146f0476348c2463943d13d3136;
    inBuf[6224] = 256'h3c2d8e234019770fd70646ff84f9b8f53ef345f27ff200f3caf3a0f4dbf4bbf4;
    inBuf[6225] = 256'h48f433f3e4f173f097eea3ec85ead1e7b2e405e170dc49d7c3d1d9cb1bc601c1;
    inBuf[6226] = 256'hadbc90b906b8fdb774b95bbc4dc0e4c4d3c9abce10d3e6d60fda73dc45dea6df;
    inBuf[6227] = 256'h95e050e1efe13ce257e23ce2a2e1b1e090df1bdebcdcdfdb85db37dc61ded4e1;
    inBuf[6228] = 256'hc4e640edacf4d9fc8a05eb0db415ba1c6622ba26e129a52b532c442c6e2b262a;
    inBuf[6229] = 256'hb028f7264925d02365225921de20d72095215223f2259c294a2ea4337639663f;
    inBuf[6230] = 256'hf544c8497b4dc74f9150bf4f7c4d174abf45f040203c75374f33ef2f292d132b;
    inBuf[6231] = 256'ha229682860277c265c251b24d2224e21d71f9c1e741da11c2c1ccd1baa1b981b;
    inBuf[6232] = 256'h2e1b8f1a9419d4179815df12600f870b81071703b8fe97fa85f6dcf2d0ef3bed;
    inBuf[6233] = 256'h61eb55eae8e942ea51ebc8ecaaeebaf098f22df423f528f548f459f24def7ceb;
    inBuf[6234] = 256'h12e74be2b3dd99d93bd6f9d3eed217d374d4c9d6d0d939dd9ee0c3e367e64ce8;
    inBuf[6235] = 256'h84e912eae0e934e934e8d2e65fe502e49ae25de161e07cdfe1dea5dea7de20df;
    inBuf[6236] = 256'h1ae069e130e357e59be719ea9fecdaeeeef0b1f2d7f3a6f423f516f5def499f4;
    inBuf[6237] = 256'h14f4a6f35ef3f0f294f24df2c5f12ff197f0bbefe2ee2cee6aedf2ececec1ced;
    inBuf[6238] = 256'hbdedd1eef2ef3af192f281f321f46df4fef306f3a8f1a9ef5fed14eb97e836e6;
    inBuf[6239] = 256'h2ee43ce293e05ddf55dea9dd7edd88ddecddcbdecfdf0de18fe2eee326e52de6;
    inBuf[6240] = 256'h9ce67ee6e0e57ee496e266e0d4dd32dbd1d89fd6e0d4bad3ffd2d4d23dd3edd3;
    inBuf[6241] = 256'h03d578d6fbd7b1d99ddb75dd63df63e122e3c6e446e651e70de877e84fe8d0e7;
    inBuf[6242] = 256'h08e7cee58be45be316e228e1aae057e07ee01de1dbe1f3e24ee483e5dbe64ee8;
    inBuf[6243] = 256'h78e9aceaf3ebf5ec0fee4aef2ff00bf1ddf11af2f7f175f11cf03aeef2ebf9e8;
    inBuf[6244] = 256'hc7e5aee28edfeedc18dbd6d996d963dabbdbc8dd67e0e9e25ce5a3e727e910ea;
    inBuf[6245] = 256'h6beadee9b7e82ce70ae5a9e240e0a4dd27dbf8d8eed646d514d42cd3afd295d2;
    inBuf[6246] = 256'hb3d214d382d3c9d3eed3afd3f6d2fad1a5d012cfa1cd60cc86cb6acb07cc79cd;
    inBuf[6247] = 256'hbbcf70d297d502d930dc39df23e2a0e42ee720ea53ed53f158f6ebfb2b02c508;
    inBuf[6248] = 256'hba0ed913a9174219e018ab168d12960daa084704c701d4015804dc09ff119d1b;
    inBuf[6249] = 256'h67265b31033b204330498d4ce64d9e4de34bdd490c488346fc455f463447ac48;
    inBuf[6250] = 256'h3a4a4f4b384cb24cb14cff4cb04dec4e73511d55af59555f5b65256b8370a074;
    inBuf[6251] = 256'h0f77ea77da7629747670d66bf6667f624c5ec65a2f58e255ea533c521350994d;
    inBuf[6252] = 256'hfc4ad047a344fd41bd3f743e5f3ef93e584010421c4356432642a93e3339cf31;
    inBuf[6253] = 256'h5628f31d6113df08b3ff72f8f2f2c4efb7eeefee4ff037f2b7f3c6f409f50df4;
    inBuf[6254] = 256'h44f2bcef5decc3e801e5f4e0f9dcdcd841d46fcf4ecab8c434bf07ba59b5c6b1;
    inBuf[6255] = 256'ha6af0caf2eb000b321b722bc7ec1a5c60acb50ce52d0fbd072d01bcf46cd62cb;
    inBuf[6256] = 256'he7c901c9dac87cc995ca0bccb1cd0ecf3bd062d152d281d36ad5f1d78edb97e0;
    inBuf[6257] = 256'h80e636ed97f4bafb450201082e0cc70e0410b90f800e050d720b8d0ae70a5b0c;
    inBuf[6258] = 256'h510fe5137c191a208927f42e37361c3dfd42ed47e74b874e0d509d500050984e;
    inBuf[6259] = 256'haa4c304a8d47f644794278400f3f513e923eb13f82411c4422473b4a554d0050;
    inBuf[6260] = 256'hf0510f530a53db51aa4f654c65480044243f333a8135e630b82c2b29ec253023;
    inBuf[6261] = 256'h1121331fca1dee1c3b1ce31be71bd81bdf1beb1b831bce1aab19ad1720150b12;
    inBuf[6262] = 256'h260ef309a5051201c4fcf4f876f5b7f2cef061efa1ee7bee89eee4ee68efbcef;
    inBuf[6263] = 256'hf6eff5ef77efa3ee6cedb7ebbfe974e7cfe419e255df96dc32da33d8a6d6c5d5;
    inBuf[6264] = 256'h80d5ced5bbd613d8aed96fdb13dd87debbdf8be01be178e18be18ce187e152e1;
    inBuf[6265] = 256'h1fe1e8e070e0dfdf2ddf27de1cdd20dc1fdb80da60daa3daa6db6add9edf6de2;
    inBuf[6266] = 256'hace5e8e838ec73ef36f2a8f4aef6f5f7b8f8f4f873f88af746f67cf48ef291f0;
    inBuf[6267] = 256'h62ee79ecf9eabde929e941e9b3e9b8ea38ecc5ed84ef56f1bbf2d8f3b6f4e0f4;
    inBuf[6268] = 256'h94f4ebf397f2eaf005efc1ec6eea49e846e6aae4a0e30fe321e3d0e3cee418e6;
    inBuf[6269] = 256'h7de78ae83ee985e90be905e89de6abe486e283e08adee3dcc5dbefda7ada78da;
    inBuf[6270] = 256'h95dad6da47dba5db05dc71dcc2dc2bddbcdd47de00dfdfdf9de06ce147e2dde2;
    inBuf[6271] = 256'h68e3e7e3ffe3e9e3ade3fee225e245e121e000df0ede22dd87dc5ddc75dc04dd;
    inBuf[6272] = 256'hfadd12df78e0f8e139e370e46ae5c6e5dde5a9e5dde4ebe3f1e2a4e175e08ddf;
    inBuf[6273] = 256'ha8de1bde02de11de73de1ddfc0df92e072e11de2e7e2ade322e4c0e47fe5fce5;
    inBuf[6274] = 256'h9ae64be78ee79fe779e7b4e69be54ee49ee2eae061dffadd0edda1dc86dcdddc;
    inBuf[6275] = 256'h64ddcfdd26de1cde92ddbedc72dbc8d930d89ad629d544d4cad3bbd345d417d5;
    inBuf[6276] = 256'h53d6e7d76cd938db25ddc7de90e089e245e45de611e903ecd3efbff446fab500;
    inBuf[6277] = 256'hd007a00eff144b1a781da51e9c1d071afc14300f2909b104a9023c038707550f;
    inBuf[6278] = 256'h6e19a425b732b63e33494351ba55335702563a525e4d4b484e43a03f763d6a3c;
    inBuf[6279] = 256'hff3cbe3edd40b943e046c549214dca506054a4585b5de6619f66046b4d6ea770;
    inBuf[6280] = 256'haf710e71536f826cdf685165f261185f815dd95c015d315ea05fdb60ec611262;
    inBuf[6281] = 256'h2a619b5f1f5d105a23573e54d3515750534fda4ed34e464e044dd64ad6464041;
    inBuf[6282] = 256'h6a3a0c3206292a2081170410590a2906da036803e9033f0509074308ed08df08;
    inBuf[6283] = 256'h75071305ed01aafdd8f8bbf306ee2ee860e252dc77d612d107ccdfc7e6c415c3;
    inBuf[6284] = 256'hc9c21cc4cec6b7ca8ecfa1d478d99ddd79e0c3e15fe139df8fdbe0d69cd155cc;
    inBuf[6285] = 256'hcdc77fc4a4c295c251c469c7b1cbced0fed5f8da8fdf50e35be6efe8f6eadbec;
    inBuf[6286] = 256'hebeee2f0fbf248f541f703f9a9fac9fbbafcebfd47ff5f01b50408098c0e3315;
    inBuf[6287] = 256'h1c1cf7226729792e02320f34583473332532bc301130c230bd323b36133b7540;
    inBuf[6288] = 256'hf745094bd44e1c51b7518e50304e104b8f47704413429c405f403d41ed424245;
    inBuf[6289] = 256'hb847fc49e44bfd4c4b4df34ca74b99490747a943cb3fb23b22377a32082e9529;
    inBuf[6290] = 256'ha2258a221320a11e461e741e3f1f65202d2191213f21951fca1ccd186a13580d;
    inBuf[6291] = 256'hf506620084fabaf5fbf1caef1cef85ef00f1fff2c1f415f67ef694f573f31ff0;
    inBuf[6292] = 256'h93eb71e60ae191dbc9d6e4d2ffcf72ce0ece9fce21d036d295d410d731d9d1da;
    inBuf[6293] = 256'hd9dbf2db2fdbafd945d729d4aad0cfcc08c9c9c531c3a0c15cc147c279c4cfc7;
    inBuf[6294] = 256'hdccb6cd00dd51ed970dcb3de8cdf3edfefdda9db08d974d61bd48fd20bd275d2;
    inBuf[6295] = 256'h0ad495d6aed965dd5de10ee58ce892ebb9ed4fef48f06df035f0a4ef89ee62ed;
    inBuf[6296] = 256'h41ec09eb47ea08ea1aeae0ea4becffed2ff099f2b5f49df604f867f805f8edf6;
    inBuf[6297] = 256'hf1f49ff249f0dfede9ebb3ea11ea4dea76eb18ed20ef52f11df36ff41cf5baf4;
    inBuf[6298] = 256'h79f37af195ee3eebe0e772e469e125df74dd8bdc93dc28dd39deb8df2be179e2;
    inBuf[6299] = 256'h8fe317e436e4fee32ae3fde1ace0f7de2add8ddbded94dd804d7cad5ded46ad4;
    inBuf[6300] = 256'h39d48dd485d5d2d69fd8e4da37dda9df08e2bbe3cce426e569e4e5e2d2e016de;
    inBuf[6301] = 256'h34db8ed828d691d413d47cd406d688d862db81de86e1c5e34de5f9e55ee5eae3;
    inBuf[6302] = 256'hdfe12edf8bdc61da90d88ed774d7d5d7ded876da1bdcf3dde2df7ae107e38fe4;
    inBuf[6303] = 256'hb6e5dde608e8c7e862e9d0e9a2e92ae976e836e7d2e573e4e2e289e18ce0b8df;
    inBuf[6304] = 256'h5fdf77df9fdfffdf80e0d4e020e150e12ee1e6e06be0b1dff0defcddc0dc7adb;
    inBuf[6305] = 256'h0ada6dd800d7d7d504d5c4d423d53cd609d844dae7dca1dfdce1a8e309e5c6e5;
    inBuf[6306] = 256'h7de6c6e7c7e936ed79f242f98601a70a5e13d71af01f7a216e1fe71952116f07;
    inBuf[6307] = 256'hc4fda6f532f17af18df6c700240f8f1fa1305e40a04cb9541858805633514d49;
    inBuf[6308] = 256'he33feb36782f0d2a8f27a6279829662d3b326037323d45434549d94faf56545d;
    inBuf[6309] = 256'h1e64666a546fd172337426733470846bd0654b60415b6b57c055e355c257875b;
    inBuf[6310] = 256'h0c608c64d368e46b746dd26db36c716aac675264f860255e8b5b785901586156;
    inBuf[6311] = 256'hba540a539250954d384ad545d740a63be93541301d2b2d26e8217f1e8c1b8119;
    inBuf[6312] = 256'h4a184b17cc1679168d154e149512cc0f600c3e08ec02fdfca8f6caef29e913e3;
    inBuf[6313] = 256'h5fdd99d8ead425d2b1d084d036d1cbd2cfd4a9d64dd85fd96fd98ed88fd641d3;
    inBuf[6314] = 256'hfbce06cab4c4a5bf4cbbf3b7f8b593b5c3b676b981bd70c299c785ccd0d0f0d3;
    inBuf[6315] = 256'hd0d5a2d64cd618d593d3f4d1b9d062d0e5d063d2d2d4a1d7cbda49de92e1dce4;
    inBuf[6316] = 256'h6ae8d6eb85effbf3e2f879fef404860be611e317a41c07202922aa22fc21b520;
    inBuf[6317] = 256'hf71ea61d871d921e4021b125272b6a312838753e04449748a14b464db64df24c;
    inBuf[6318] = 256'h804bb34991478345ac430442d7402d40fa3f6b405941ae427c446b463d48cd49;
    inBuf[6319] = 256'h904a4d4afe486946de42c73e3e3ade352632142f162d4f2c412cde2cc52d282e;
    inBuf[6320] = 256'hfd2d032da92a57274123411e0619f313f90ebd0a7807e00441036e02de01bc01;
    inBuf[6321] = 256'hc0016201d500d3ffdafd34fbcbf766f38fee68e9eee3bede06daded5dbd214d1;
    inBuf[6322] = 256'h76d038d103d36dd554d81edb4fddc1dee7de82ddcbdab7d696d117cc9ac6a8c1;
    inBuf[6323] = 256'hd8bd58bb6fba35bb48bd83c088c49ec888ccfbcf70d2f8d395d412d4cbd2f1d0;
    inBuf[6324] = 256'h81ceffcbaac988c724c6b1c525c6ebc7edcad1cea5d3e6d8e3dd85e243e685e8;
    inBuf[6325] = 256'h8ce93ee983e719e55de288df69dd42dc08dc27dd74df88e287e60deb8bef13f4;
    inBuf[6326] = 256'h3af879fbfefd89ffc0ff02ff4dfd83fa49f7f0f399f002ee77ecdfeb8cec63ee;
    inBuf[6327] = 256'hdff0f0f335f708fa50fcccfd1cfe80fd1ffce8f94df793f4abf1ffeed5ec15eb;
    inBuf[6328] = 256'h0eeae9e967ea9aeb7ceda4eff1f12af4c3f58cf669f615f5c4f2d2ef5cecd5e8;
    inBuf[6329] = 256'hb8e526e36ce1cae017e13be20ae413e61fe804ea78eb82ec2ded4bedfcec62ec;
    inBuf[6330] = 256'h61eb29eae6e881e71fe6e4e4c1e3e9e286e28ee223e33ce49ee547e703e97cea;
    inBuf[6331] = 256'hb5eb7eec81ece8ebbaead8e8a7e670e434e265e045dfc5de2bdf79e05ce2d0e4;
    inBuf[6332] = 256'h8de70eea4bec0beef0ee32efdbeec4ed64ecf9ea76e94be891e7fbe6b2e69fe6;
    inBuf[6333] = 256'h64e62ee6ffe59ae540e502e5bae4bee427e5bde59fe6a8e76fe8f0e80fe9a5e8;
    inBuf[6334] = 256'he5e7cee662e5f3e37fe20ee100e044dfabde5dde3dde21de30de7dde16dfffdf;
    inBuf[6335] = 256'h0de14ae298e38de446e5d2e5d9e5b2e5ede5ace692e83eec98f198f8cd002609;
    inBuf[6336] = 256'hd010b0168619fb18d714300d880370f950f068ea24e9c8ecc2f552038713dc24;
    inBuf[6337] = 256'h3d354842f44a734e704c3946173d4e320d28951f71199f16f816ac199e1ee924;
    inBuf[6338] = 256'h902ba932b5393940c246f34c3252c456185a775b265bf358e254e54f7a4a6845;
    inBuf[6339] = 256'hfc4180403e41af44fe4961508457215e566304677f68b46743654c61785cb357;
    inBuf[6340] = 256'h2053454f9f4cd84a1f4a934a8a4bf24c994e924fc14f094fbf4c2a498e44ad3e;
    inBuf[6341] = 256'h29389531042b5225f720c31d1d1cd71b2e1c291d531eda1ed61ef01d891b0918;
    inBuf[6342] = 256'h7d13ac0d5707cd0002faaff316ee21e963e5e7e262e10fe19ae16fe290e392e4;
    inBuf[6343] = 256'hebe4b7e4c1e3b4e1d3de2fdbbbd6e2d1f5cc22c8dcc37cc033be45bddbbde0bf;
    inBuf[6344] = 256'h23c350c7dbcb23d0a5d3ecd59ed6c7d58ed32ad048cc8bc84cc544c3e4c203c4;
    inBuf[6345] = 256'hc9c634cbafd01ed761decfe543ed87f4e6fa3e006104a30620070006140324ff;
    inBuf[6346] = 256'h17fb5cf71af538f5c3f72efd6905760fc61a7626fd30a839ec3f104360435c41;
    inBuf[6347] = 256'h4f3d3938f8320e2e722aad28cb28202b782f3835273cae43004bbf514a57f85a;
    inBuf[6348] = 256'hab5c395caf599c556d50af4a19450b40fd3b583909382838a339e03b9f3eac41;
    inBuf[6349] = 256'h6944a9464c48ce480e48ef452742043dcf36b52f8828d521db1b6c17d814e313;
    inBuf[6350] = 256'hba14eb167919f91bb51dd31d5e1c3f196014790efb072e01f4faa3f544f142ee;
    inBuf[6351] = 256'h69ec50eb12eb4aeb87ebf2eb33ece1eb2bebd1e991e7b9e437e10addaad834d4;
    inBuf[6352] = 256'hf5cf7dccd2c910c881c7e3c7ffc8c8cac6cca8ce4dd049d182d108d1b7cfcecd;
    inBuf[6353] = 256'h9ccb2ec9e4c618c5d9c37bc322c49dc5f8c7f2ca0cce2cd1fdd310d67fd734d8;
    inBuf[6354] = 256'h11d88dd7dcd614d6c8d50fd6c3d630d82ada53dce1dea0e13ce4f4e6a3e901ec;
    inBuf[6355] = 256'h52ee67f0f0f11ff3bdf37ff3c7f2a5f120f0eaee4eee5dee9def0ff252f56ef9;
    inBuf[6356] = 256'hf0fd1202a1052c081f09aa08f6060b04920011fdb7f913f76ef5a4f4e3f411f6;
    inBuf[6357] = 256'hb3f7b1f9cffb88fde3fedcff1b00c6fffafe67fd35fba0f880f519f2c8ee81eb;
    inBuf[6358] = 256'h90e858e6cde42ae4a1e4dde5bfe70fea2decdbedf1eef4eeefed17ec46e9dbe5;
    inBuf[6359] = 256'h5fe2ecdef5dbe7d99ed833d8b2d8b2d921dbeadc97de16e04fe1d7e1c6e13ae1;
    inBuf[6360] = 256'hf6df47de67dc2cdafbd724d693d4b5d3c0d363d4b7d59ed790d98adb66ddabde;
    inBuf[6361] = 256'h75dfbbdf32df41de2addd1dbb2dafad966d944d9a8d94ada75db28ddfade0ee1;
    inBuf[6362] = 256'h41e321e5d9e64ce80fe94fe901e9eae77fe607e583e373e2f4e1d5e156e260e3;
    inBuf[6363] = 256'h9de428e6c5e7fee8eae971ea65ea17ea9be9dbe813e843e762e6b9e544e5fde4;
    inBuf[6364] = 256'h19e55ce599e506e67ee6e0e661e7f1e775e809e9ade978ea6feb4fec09ed75ed;
    inBuf[6365] = 256'h23ed36ec05ebabe9c1e805e9c4ea70ee41f4cffb9404840d1c15421adc1b1919;
    inBuf[6366] = 256'h7312c10829fddbf1d0e874e363e327e909f41f03751467250e34913e8f433143;
    inBuf[6367] = 256'hee3da6347329031ea413240c3908af079b0a341045176b1fd827c32f4737ee3d;
    inBuf[6368] = 256'h2a434e47024acf4a224ae347e943043fae39703480306d2e892e58315c36e53c;
    inBuf[6369] = 256'h9b445c4c24539e580a5c015ded5bec5874546f4f3e4a634581419c3eeb3cb03c;
    inBuf[6370] = 256'h913d7b3f4b4243450e485b4a604be94adf48d644233f39385a307a2865216f1b;
    inBuf[6371] = 256'h58175515fd145b16ea18a41b321eed1fec1f401eec1acb159b0fdb08b80105fb;
    inBuf[6372] = 256'h20f50ff05becf8e977e8fae725e85fe8cee83ee92fe9c8e8f1e746e600e439e1;
    inBuf[6373] = 256'hd9dd2bda4fd648d275ce1dcb6dc8d3c682c656c73fc902cc29cf4dd212d5fbd6;
    inBuf[6374] = 256'h9fd7dfd6b7d45fd17bcdacc973c680c42fc468c554c8d4cc3cd231d84fdec9e3;
    inBuf[6375] = 256'h63e825ece0eef3f0aaf2e2f3e4f4c1f516f632f645f605f6f2f58bf6d2f792fa;
    inBuf[6376] = 256'h73ff4e064b0f101a4f2520307239db3fd34218427b3df135b72c0b23ea1ad115;
    inBuf[6377] = 256'h77149417ec1e5a29e7351f43444f3559e75fae62cc61aa5d0857354f0c47483f;
    inBuf[6378] = 256'hcd38f633f73015301b31df332a385a3d23433849bc4e30532256ab567d54b24f;
    inBuf[6379] = 256'h58482f3f2535012b03220d1b8b1639150717111bd3203027972c6530ef318530;
    inBuf[6380] = 256'h7a2c1526941d14146a0a330192f9e2f30cf05fee65ee77ef9df136f46ef630f8;
    inBuf[6381] = 256'he6f8f3f798f5d1f1a5ecaee61be034d9bdd202cd6cc8b5c5c8c472c5b9c7faca;
    inBuf[6382] = 256'h93ce3cd245d51fd78ad727d60dd3acce60c9e9c308bf10bb86b8bcb78db8fdba;
    inBuf[6383] = 256'hc2be2dc3d9c738ccb2cf35d29cd3d0d331d3d6d1dccfdecd0ecc8bcaeec944ca;
    inBuf[6384] = 256'h75cbdfcd58d19fd5d8da84e012e668ebdaefe6f2c3f43cf548f499f26bf008ee;
    inBuf[6385] = 256'h50ec89ebd4eba0ed9cf04ff4b2f834fd550133057708ce0a7b0c5f0d620df70c;
    inBuf[6386] = 256'h240cd30a6509d8071906ab04cf0391035204120680088b0be70e1412e514fb16;
    inBuf[6387] = 256'hd6176e17c215ca12030fe50aa306b70280ff03fd83fb32fbd9fb5cfd90ffe701;
    inBuf[6388] = 256'h0904c1059a0671064b05ff02bbffe6fbaef790f31bf060ed8bebc5eab6ea2beb;
    inBuf[6389] = 256'h0fecf5ecabed24ee13ee8aedb8ec7deb0aea9ae8eee618e54ee368e198df2cde;
    inBuf[6390] = 256'h07dd4bdc1cdc37dca2dc52ddd8dd1bdef8dd12ddaadb0eda37d8a2d6a3d5fbd4;
    inBuf[6391] = 256'hdcd465d535d64ad794d893d93fda9ada7cda48da31da01dafad915daf1d9ddd9;
    inBuf[6392] = 256'hd8d9aed9dcd976da22db15dc55dd82debbdfcce022e1d4e0ebdf4ede96dc29db;
    inBuf[6393] = 256'h0bdaaed926da2ddbecdc39df9fe10ce426e687e75fe89be82de880e786e60ae5;
    inBuf[6394] = 256'h60e393e1a6df14de2bdd19dd1ade17e006e3bde697ea39ee5cf150f30bf412f4;
    inBuf[6395] = 256'hb0f3a6f3dff4b2f750fc70022809a70fbc140d172f16ee11750a5a015bf805f1;
    inBuf[6396] = 256'h6eedc2eefbf4f2ff640e211e632d003af541b9440f42793a083076244619a210;
    inBuf[6397] = 256'h800bfa098d0c9d12ee1ae3243b2fc3385b416c48934d60517b53825314521c4f;
    inBuf[6398] = 256'h904a7e456240ac3b74381c37f937ab3bb2416a496a52385b9f624368446b576b;
    inBuf[6399] = 256'h1d69c464e95eac5897526f4d084a50485d48274ade4c2f50d853ee563359815a;
    inBuf[6400] = 256'h145ae7572f54b44e0248b640f6389131242bcc254322bd20bd205a220f25b627;
    inBuf[6401] = 256'h072a7e2b362b43299725e81fea182511dc081e0171fadbf4f2f0b4eea9edf6ed;
    inBuf[6402] = 256'h30ef87f0d4f185f2f2f156f0b0edd9e959e56ae012dbe6d538d125cd17ca14c8;
    inBuf[6403] = 256'he4c696c609c712c8bdc9cccbe4cdc1cf08d16ed1e1d05dcff3ccc7c91ac64fc2;
    inBuf[6404] = 256'hd5be4bbc4bbb04bc90beddc25bc89ece49d596db0fe169e514e813e9c4e847e7;
    inBuf[6405] = 256'h44e572e3eae126e1a1e12ce30be67beafcef7bf6d6fd41058b0c9213a1199f1e;
    inBuf[6406] = 256'h6e226924be24cd238c21b91e141ccd199918fb18dd1a951e0f24872aa031af38;
    inBuf[6407] = 256'haf3e5e43784698471e47544566421c3f0a3c94394f3848384e394f3bc83d5340;
    inBuf[6408] = 256'hd042c84402468a462e460e459243cb41f63f4d3e923cd23a2a396f37e0359634;
    inBuf[6409] = 256'h43331d32383149308e2f0d2f472e2f2d842bca2844252621741cca1764133d0f;
    inBuf[6410] = 256'heb0b8809d8071207d1066206b1055b04010205ff74fb52f73bf354efa1eba8e8;
    inBuf[6411] = 256'h61e698e46ee37be25be124e096de9cdc94da6dd82dd62ad440d273d00ccfd0cd;
    inBuf[6412] = 256'hc6cc0acc49cb8eca09ca96c95ac97ac9aec9e9c928ca22cae0c967c987c877c7;
    inBuf[6413] = 256'h5ac619c515c494c388c32ac476c524c743c9a9cb06ce6fd0a7d25bd4bed5ced6;
    inBuf[6414] = 256'h72d70bd8a7d830d9f4d9dedac2dbeedc50debadf69e13ae3fbe4f1e608e91ceb;
    inBuf[6415] = 256'h5fed8eef5cf1f4f22bf4ddf45ff59ff585f563f535f5fcf425f5a4f551f667f7;
    inBuf[6416] = 256'hb4f8f4f94cfb95fca0fd9bfe59ffafffd2ffb6ff57ff01ffa2fe1bfea8fd2ffd;
    inBuf[6417] = 256'h94fc23fcd5fb8afb72fb78fb70fb81fb9efb99fb88fb50fbc6fa0bfa18f9e9f7;
    inBuf[6418] = 256'hc3f6aff590f493f3b2f2c6f1fff069f0e1ef89ef56ef09efadee43ee98edb1ec;
    inBuf[6419] = 256'h87ebfce92fe83fe63de48ce259e192e070e0f9e0d1e1f3e24be44fe5c2e5c5e5;
    inBuf[6420] = 256'hd9e42ce341e1eadeaedcf3daa1d9f5d813d9b9d9e5da68dcc3dde9dec1df04e0;
    inBuf[6421] = 256'heddf91dfbfdebfdda1dc44db18da47d9afd89fd805d98cd974daa3dbbddce7dd;
    inBuf[6422] = 256'he7de5ddf83df49df95dedfdd35dd80dc1adcdddba4dbcfdb36dca9dc74dd4fde;
    inBuf[6423] = 256'hf8decbdfa8e079e18ee2a2e380e447e593e55be5f4e40de4b1e258e1dadf6bde;
    inBuf[6424] = 256'habdda3dd7cde75e01fe345e6abe996ecd6ee54f077f06aefaced69eb80e9f1e8;
    inBuf[6425] = 256'h22ea9fed7ff30afbaa033b0c1f136b174018ed141b0ee504b0fac9f10dec9cea;
    inBuf[6426] = 256'h86eeacf7d9049f14b424b832153d37427a41cc3b46328e261d1baf11970b0e0a;
    inBuf[6427] = 256'h040dd913ce1d3929a8342a3f6e470e4d6c5062515a502b4ecd4a98466342763e;
    inBuf[6428] = 256'h1e3b15397938af39283d73427649be51ef594361fb66f0690c6a9667a2623a5c;
    inBuf[6429] = 256'h6b55c74e6949ff45834459453948224cbb505255e758725bb25c245c345afe56;
    inBuf[6430] = 256'h4052964c6346c93f8b39dd33b32ecb2a3c28c126e1266128632ac32cdb2eb22f;
    inBuf[6431] = 256'h3d2f312d2a29b8231f1d9d155b0eea077e02e1fef5fc14fc4afcfbfc44fd34fd;
    inBuf[6432] = 256'h66fc3efa1bf725f364eea3e932e514e1cbdd42db34d9f6d744d7aed65ed603d6;
    inBuf[6433] = 256'h3bd563d491d3b8d234d2f9d1bfd18bd128d16ed079cf17ce37cc2fca34c892c6;
    inBuf[6434] = 256'hdbc56ac654c879cb88cf0dd46ed832dc29dfffe080e1e1e074dfc8dd8bdc31dc;
    inBuf[6435] = 256'h1fdd4ddf1fe23ee54ee8b0ea70ecd7edcceedbefd7f119f53bfa8d015c0ab413;
    inBuf[6436] = 256'h901c6023202783274224271e5916f90df8060503ef0273075010021c2d294136;
    inBuf[6437] = 256'h7741e149d14ed24f664d36481c41b5392433fd2df22a022abc2a122db0303435;
    inBuf[6438] = 256'h7d3a01404945264afa4d5c5041513150e84ca147924082389e30ca290e250b23;
    inBuf[6439] = 256'h9823a626ce2bf9316a38373e044239439641fa3c3636342e95256c1d6716c110;
    inBuf[6440] = 256'h340de30b4b0c340ece100713a6145315b5144f133a11380ea00a7a06bb01f3fc;
    inBuf[6441] = 256'h42f899f35aef6debd2e73fe5eee3cae3ece4bae665e8a6e902ea33e95ee758e4;
    inBuf[6442] = 256'h1fe034dbf4d508d150cd1acb7eca75cb60cdb4cf21d228d480d5fcd565d5f5d3;
    inBuf[6443] = 256'h10d209d07ccec1cdb0cd2dceeace7dcfebcf37d05cd0a9d02bd1d8d1f8d299d4;
    inBuf[6444] = 256'hb5d672d961dcf0de0fe18ce24ee3bde3f1e3f5e328e48ce42fe584e67be8d9ea;
    inBuf[6445] = 256'h9aed42f070f261f419f6a0f760f946fb20fd0effd50036023f039503e1025b01;
    inBuf[6446] = 256'h30ffd0fc24fba7fa88fbf8fd8f01a905f609ef0df010b412f1127811b10e310b;
    inBuf[6447] = 256'h8e0778044802fb009400eb00cb01430329050c07bf08240afe0a770bd90bf70b;
    inBuf[6448] = 256'ha20bb20ac608d2051702c4fd55f962f525f2fcef56ef2cf07bf21df63efa1afe;
    inBuf[6449] = 256'h1e017f020302ebff33fc35f78cf170eb7ee58ee0eddcf1dacedaf1dbfeddbee0;
    inBuf[6450] = 256'h87e314e642e86fe97ee9a2e8c7e669e40fe296df31ddf9da7ed802d6f3d327d2;
    inBuf[6451] = 256'hf0d09ad0d5d0cad1a3d3f1d599d835dbdfdc6dddd0dcc8dafbd7fad4d0d11ccf;
    inBuf[6452] = 256'h3ecd0dccf0cbffccacced6d00ed394d479d5c6d54ed588d49bd352d20ad1e0cf;
    inBuf[6453] = 256'hcdce4ace55cea1ce5ccf50d03cd183d217d4b3d57ad717d914da92da9dda55da;
    inBuf[6454] = 256'h1bdaebd9d0d9f1d9fbd901da56dab6da29db24dca8dd0ce003e4b9e928f1d4f9;
    inBuf[6455] = 256'h8702290a8c0f70119d0f3e0a900100f768ec64e317de26dee7e338efe7feb910;
    inBuf[6456] = 256'hb1228132d73da1434443bf3cbe3145245316a70a25037a003603d50ae6153b23;
    inBuf[6457] = 256'h0c31783d9047494e08518650354d8f47fb40363a9c33492ed42a8329e62ad02e;
    inBuf[6458] = 256'hcd34973c21458d4d8355de5bbd5f1f61915f1e5bcf54644dc5452b3f153aff36;
    inBuf[6459] = 256'h5f36e4375f3b7740f645154b514fb9512e5204510e4ea4494b44023e5137cb30;
    inBuf[6460] = 256'h902a39251c21fd1d371cd71b621cf51d44205522d4234d2407233720171cb416;
    inBuf[6461] = 256'hca10c60ad504c3ffd1fbe4f860f7fef608f76cf7c0f770f79ff638f509f36ff0;
    inBuf[6462] = 256'h84ed5cea7be7f7e4bde201e181dfe3dd41dc81da8fd8bad61ed5c5d3ead29dd2;
    inBuf[6463] = 256'he0d2b5d3e0d424d644d7f3d702d862d71dd655d428d2dacfc5cd22cc54cbabcb;
    inBuf[6464] = 256'h0dcd6fcfbdd280d67cda8bde3fe27ae527e8e7e9d8ea2eebd0ea2beaa3e919e9;
    inBuf[6465] = 256'h05e9e9e9b8ebd7ee86f340f9c9ffae06010d7a12cd165f195a1aed1903186c15;
    inBuf[6466] = 256'hf212e5102010181187139017fc1c13239229ee2f42354e39c13b4b3c6b3b8539;
    inBuf[6467] = 256'hda362f34ef314230b32f6130303233350539273d5d411a45f547eb49aa4a174a;
    inBuf[6468] = 256'h7b48e1459442243fcc3bf138e3368135f2343535dd35ec364a386039123a423a;
    inBuf[6469] = 256'h7539c4374635d831df2d9529ff24bc20181d021ae617a516b6153415d5140514;
    inBuf[6470] = 256'he9124a11ac0e5c0b6607c9023afe01fa26f62bf3f8f04aef6cee0feeb7ed65ed;
    inBuf[6471] = 256'h94ecc9ea48e808e519e11ddd2ed95cd51bd262cf35cde9cb44cb0fcb4ccb9acb;
    inBuf[6472] = 256'hdccb41cc96cce2cc43cd64cd30cdb5ccbccb6fca07c970c7e6c596c470c3c7c2;
    inBuf[6473] = 256'hc2c23bc353c4ddc574c728c9d1ca3bccaecd13cf32d059d175d264d388d4ced5;
    inBuf[6474] = 256'hffd656d8a2d9bbda06dc73ddf7def5e02ae360e5e8e780eaf4ec91ef0bf21ff4;
    inBuf[6475] = 256'h17f6bdf7f0f80afad7fa2cfb55fb33fbdbfaddfa4cfb45fc29febd00c3035107;
    inBuf[6476] = 256'hf10a310e0311fe12da13d61306138a11d00ffa0d190c760a20092708d0071a08;
    inBuf[6477] = 256'hed08590a310c280e2d100a125a13f613bc1371123210480de1095c0622035a00;
    inBuf[6478] = 256'h3bfefefc90fcebfc05fe79fffe0068025303a7038b03df02b001320030fea7fb;
    inBuf[6479] = 256'hdcf8bff57bf27cefc7ec8aea1ce962e864e835e95dea8feba1ec09edacecbceb;
    inBuf[6480] = 256'h11eae1e781e5d1e20de08cdd2fdb35d9e6d702d7a0d6e5d66ed737d84bd93cda;
    inBuf[6481] = 256'h08dbb2dbe4dbc7db76dba7da98d96bd8d1d618d57ad3bdd13dd03bcf86ce68ce;
    inBuf[6482] = 256'hfecef9cf73d142d3ead475d6abd723d81cd890d747d6bed430d394d183d03ed0;
    inBuf[6483] = 256'h9bd0d6d1c6d3f6d55bd89bda5fdccadd9edeb7de87de06de36dda6dc5adc32dc;
    inBuf[6484] = 256'h7bdc23dd13de88df60e186e3f6e525e8d0e901eb5aeb00eb8bea26ea4deab8eb;
    inBuf[6485] = 256'h99ee25f357f97200bd07360e8b122814cc12490e9207efff72f8cef27bf014f2;
    inBuf[6486] = 256'h12f80f02a40e601c56298333ed39d23bfe38af323a2af8201119f9133c126d14;
    inBuf[6487] = 256'h1c1a15225f2b9034603c5d42e445ca46e2457943fa3f8f3c8c3901378f352d35;
    inBuf[6488] = 256'hb0356f37313ac93d50422547d64b4c50a75363559955c553e64fcc4ad744d43e;
    inBuf[6489] = 256'hea398a362f352f36f738223d3342f346bc4a324d8d4de94bd8487c448e3fca3a;
    inBuf[6490] = 256'h3c364c32262f712c592ad72869274f269525cd2448242024d0236123a122fa20;
    inBuf[6491] = 256'h801e2a1bd7161f12490d69083f04070199fe62fd35fd67fdd3fdf7fd23fd5cfb;
    inBuf[6492] = 256'h8ff8b9f479f028ec14e8ece4d0e2a2e17de1e0e122e20ce231e149dfacdca2d9;
    inBuf[6493] = 256'h7fd6e3d331d298d132d2c6d3edd52ed8f8d9f1daebdad4d9e1d76cd5d4d286d0;
    inBuf[6494] = 256'he3ce3eceb7ce2cd084d285d5bcd810dc73df8ce25ee5fce719eac3eb22edfbed;
    inBuf[6495] = 256'h69ee8aee33eeaded43edf5ec45ed6dee25f0acf205f6b1f9e6fdc202e207740d;
    inBuf[6496] = 256'h89139d19911ffd2400294c2b752b1129c024371f221907141311d8102414ff1a;
    inBuf[6497] = 256'h97242b30563c6a4759500756bb57c4557d509e48aa3fd1362d2f072ae627e728;
    inBuf[6498] = 256'hf92c4d33043b5343084b5951dd55da572a571854ad4e7e476f3f16376d2f5329;
    inBuf[6499] = 256'h2a259223a724ce27b22c7932bb37cd3b053e9c3dcf3af3353d2f9d27c51f1e18;
    inBuf[6500] = 256'h94117b0cc108c5063606750694071009340a130b410b380a4a086805780106fd;
    inBuf[6501] = 256'h16f89cf21aed88e706e23edd3ad90fd642d494d3c0d3e1d45ed6a7d791d888d8;
    inBuf[6502] = 256'h54d735d51fd26bceaacaeac684c3edc009bffbbde5bd5cbe3ebf64c054c10dc2;
    inBuf[6503] = 256'h8fc29ec286c278c25dc295c233c3efc3dfc4c1c520c621c6bac5e7c44bc430c4;
    inBuf[6504] = 256'hb6c463c622c9a0cceed089d5dad9d9dd04e1f7e204e41ce458e375e2a2e10fe1;
    inBuf[6505] = 256'h59e179e25be44ce7e8eacceef5f2dcf62ffa2bfda0ff88014603a50480051e06;
    inBuf[6506] = 256'h52060f06be056405190553052706a907150a260d8010ec13de16ed181c1a421a;
    inBuf[6507] = 256'h5819bf17a91549131b11690f4b0eeb0d3e0e040f1a10551173125e1301143814;
    inBuf[6508] = 256'h1014a013dc12e011c210550f980dad0b7e0935073005730320026c0124012501;
    inBuf[6509] = 256'h6a0190015801b90066ff64fd07fb59f8a4f552f347f18def4bee30ed33ec79eb;
    inBuf[6510] = 256'haeeabee9c9e87ee7efe568e4c4e224e1bddf3edeb1dc47dbc6d959d839d714d6;
    inBuf[6511] = 256'hf8d407d4f5d2f8d14dd1abd039d011d0dbcfc8cf0bd053d0b5d021d10fd183d0;
    inBuf[6512] = 256'h85cfe5cd11cc55caa6c887c73ec7a7c717c97acb2fce04d184d305d595d533d5;
    inBuf[6513] = 256'hc2d3bdd16acfefccfacaddc9bbc9fbca60cd73d024d4e9d73edb35de74e09ae1;
    inBuf[6514] = 256'hd3e117e181dfaeddf3dbb4da67dae8da3adc81de3fe136e46fe75aeac9ec0def;
    inBuf[6515] = 256'h33f1a6f3eff6fbfab9ffc6042209430ca90d930c32091304aefd7cf71bf399f1;
    inBuf[6516] = 256'h28f425fbb605db12db20752d3737c63c143d9a383f304a25351a1c115c0b5c0a;
    inBuf[6517] = 256'h340ee0157b20502c7337e2406c47464a034a0f471b42c93ce937e3338631bd30;
    inBuf[6518] = 256'h37313a3360364c3a203f2944e4486b4d0951515387542b541052da4eb04a2146;
    inBuf[6519] = 256'h4042573fbf3de53d3a3f764185447247cb49754bb04b7e4a734891456c42b33f;
    inBuf[6520] = 256'h343d133b6939a937e4352934fe31a72f642df32ada287d277526db258225a324;
    inBuf[6521] = 256'h2e231821171ea71a0e173113a70fa80c000a1808e906e105ff04ff0360025400;
    inBuf[6522] = 256'he3fdf1faf4f708f523f2c5effeed9beccbeb42eb71ea44e983e704e51de20bdf;
    inBuf[6523] = 256'h09dc8fd9d1d7f4d62fd761d841da8adcb3de3fe0ebe083e000df8cdc6bd9fed5;
    inBuf[6524] = 256'ha7d2f3cf6cce4aceabcf82d24bd68adae5ded7e21de6a0e820eabbeaadeaf8e9;
    inBuf[6525] = 256'h0de94fe8a2e748e788e73de8bbe95fecf9ef95f40dfaacff31054e0a540e3a11;
    inBuf[6526] = 256'hf612261330129710920eef0c500cc60cb00e12126d16ae1b6a21cf26992b5e2f;
    inBuf[6527] = 256'h8e316a3236321731be2f9b2ecb2db52d612ea62fa6311c34ac3649398b3b1d3d;
    inBuf[6528] = 256'h173e503ec03db93c423b8839f0379236ac357235a2351e36b736e936a636fd35;
    inBuf[6529] = 256'hb134fe321831da2e8e2c6c2a542889260b2583231622b220131f891d121c5d1a;
    inBuf[6530] = 256'ha418d1169d1459120210540d900a96073304de00b8fdc9fa8bf8eff6acf5edf4;
    inBuf[6531] = 256'h64f4b0f3e1f299f186efdcec8fe9c4e51be2beded3dbb4d933d82bd7bad693d6;
    inBuf[6532] = 256'h86d697d670d6f4d53fd531d4f3d2bcd177d04acf51ce65cdadcc3ccce3cbb8cb;
    inBuf[6533] = 256'hb3cb99cb89cb88cb84cbbccb2fccbbcc8fcd87ce7bcfaad0f6d131d393d4e7d5;
    inBuf[6534] = 256'hfdd61ad827d914da32db5fdc84ddecde73e009e2f7e3fae5dde7c9e974ebc1ec;
    inBuf[6535] = 256'h05ee1fef0af016f118f201f321f453f585f6f1f762f9b7fa26fc8ffdeafe7600;
    inBuf[6536] = 256'h1902c103990576073609ed0a630c650d0d0e480e100eaf0d4d0df70cf00c4f0d;
    inBuf[6537] = 256'hf80df10e201040113112dc120c13ce123d12521139102a0f1e0e330d960c1a0c;
    inBuf[6538] = 256'hb90b850b340baf0a120a2609f007b6065e05fa03cd02a30170005bff1ffeaefc;
    inBuf[6539] = 256'h36fb6ff95df743f5eff28af07bee9aec00ebfae934e99de85ae8f8e74fe76de6;
    inBuf[6540] = 256'he5e4bfe24ee07adda7da58d86dd625d5bbd4bdd41cd5cfd532d622d6a6d550d4;
    inBuf[6541] = 256'h56d217d077cde7cad5c820c72cc637c6ebc666c88ecab3ccbece78d03fd132d1;
    inBuf[6542] = 256'h69d0a0ce57ccf0c96fc773c553c4eac391c443c67dc851cb77ce4ed1dbd3dad5;
    inBuf[6543] = 256'hdad625d7c7d6b1d58bd497d3d3d2ced28cd3bfd499d6e2d833dba7dd01e002e2;
    inBuf[6544] = 256'he3e36de579e653e7c0e78fe71be750e62ce531e483e34ae3ece35de5a2e7d7ea;
    inBuf[6545] = 256'h8bee78f27cf6e7f964fc02fe86fe2efe94fdfffcfcfc00feedffc30232065309;
    inBuf[6546] = 256'hab0bc70c130ce409e506b00384016301a903bf084e1030197822c52a8a302f33;
    inBuf[6547] = 256'h4d32e02d1e27441f8417ab11c40e210f2a13421a2023d72ce935ef3c82412043;
    inBuf[6548] = 256'hc1416c3ec1396c34b42f0e2ca129fd28e929092c792fab333038173db5419445;
    inBuf[6549] = 256'hc948b14aed4ad14931474043dd3e623a6d36da33b2321e335435a0388f3ce340;
    inBuf[6550] = 256'ha4445147d948b84809475244a7409b3cd1384e3572327f30032f012e6c2da62c;
    inBuf[6551] = 256'hbe2bd42a932942282527f225d124c9236d22cd20d31e251c0d19ae15ea11510e;
    inBuf[6552] = 256'h300b660857061c055804180431042b04fb0367032102610033fe92fbf5f889f6;
    inBuf[6553] = 256'h39f441f28ef0cfee01ed02ebade83de6e6e3d9e182e023e0bfe055e2a7e438e7;
    inBuf[6554] = 256'h87e917eb7deb88ea41e8e7e4e4e0cddc35d996d66fd5fad50fd87cdbd0df4ee4;
    inBuf[6555] = 256'h7de8f3eb3eee69ef9befe6eed5ede3ec2dec1dece1ec27eee9ef12f249f4a7f6;
    inBuf[6556] = 256'h3af9d6fbc6fe16027e053609240db210dc137616fd179c188b18d117fc167016;
    inBuf[6557] = 256'h4b161017d7185f1bc81eb8228326082aee2cce2eeb2f68305630343026302230;
    inBuf[6558] = 256'h6030b630e330f830bc301a30542f722eab2d6c2da82d642eb52f2e319332cd33;
    inBuf[6559] = 256'h7c3490341a34ed324431592f1f2df42a0729212777250f249e225b215420441f;
    inBuf[6560] = 256'h631ea71dc61cfc1b3a1b2e1a07199917861515134510f90cb40985064b037200;
    inBuf[6561] = 256'hf5fdaafbf3f9bdf8c0f730f7caf638f6a0f5c0f44df374f1fceecdeb58e8b7e4;
    inBuf[6562] = 256'h1ce110de9bdbb7d998d802d8c7d7f6d741d87cd8b4d8b1d874d831d8ced75bd7;
    inBuf[6563] = 256'hf0d657d693d5b3d49fd38ad29dd1d3d065d06ad0d3d0ced154d332d560d796d9;
    inBuf[6564] = 256'h7ddb13dd29dea7ded6deb3de42dee0dd93dd66ddb8dd7fdea9df64e17de3cce5;
    inBuf[6565] = 256'h7ae84ceb14eee5f067f361f5fcf612f8a4f811f953f96ef9b8f92afac9fadffb;
    inBuf[6566] = 256'h58fd14ff2f017403b4050c084f0a580c3f0edb0f0311e5117e12b912c812aa12;
    inBuf[6567] = 256'h38129311d010e50f0c0f6b0ef30dc30de50d2b0e9e0e3d0fba0f08101e10aa0f;
    inBuf[6568] = 256'hb30e610d890b4b09f2066204c80184ff85fde7fbe2fa27fa9bf94df9dcf83ef8;
    inBuf[6569] = 256'ha0f7abf662f504f43cf219f0ebed6aeba4e8efe515e349e0fddd10dcb3da2dda;
    inBuf[6570] = 256'h1bda72da46db0bdca4dc13ddbedc92dbbad9e3d65fd3b6cfe5cb65c8b9c5bac3;
    inBuf[6571] = 256'habc2bac26cc3b9c47cc60bc85dc967cab6ca85ca01cadcc86fc7efc52ec49cc2;
    inBuf[6572] = 256'h7ac19fc072c006c103c2a3c3c0c5ddc711ca1ecc8acd8bce11cfecce9bce3ace;
    inBuf[6573] = 256'hb3cd85cdb7cd1fce20cf95d02dd218d404d69ed732d99edad0db3addbfde42e0;
    inBuf[6574] = 256'h11e2ebe3a6e57ae70ce932ea2debc0ebf4eb47eca0ec10edeaedf5ee2ff0d8f1;
    inBuf[6575] = 256'hb9f3eaf598f856fb17fee300330302057e065c07d8075c08f208120a1c0ce00e;
    inBuf[6576] = 256'h70127d16301a3b1d301f6c1f391eee1bc518d015f613a913b9153f1a91203128;
    inBuf[6577] = 256'hf02f5f36d43a823cf53af0361d315a2a622440207d1ed11fdc23a92997306737;
    inBuf[6578] = 256'hfd3c1c41324319439441da3e523b0b383535e532a231223132313132d2330036;
    inBuf[6579] = 256'h0b39673cb63f03439045f6465d474b46bf4356402b3cd5375134cf31b1305b31;
    inBuf[6580] = 256'h3833f1354739423c763ec43f963f113eb63b85380f35f1310f2fa52cd42a1f29;
    inBuf[6581] = 256'h8a27162655248722e720371fd61d021d581cf21bbb1b201b151a7418de159c12;
    inBuf[6582] = 256'hd90e950a7306d202b0ff89fd74fc14fc69fc21fda1fdc0fd2dfd9cfb4ef96bf6;
    inBuf[6583] = 256'h18f3e8ef19edb1eae9e8a1e786e686e566e4f1e246e178dfa6dd25dc28dbccda;
    inBuf[6584] = 256'h2bdb28dc8cdd0fdf51e004e1f4e007e053de12dca1d970d7d3d528d5a9d52ed7;
    inBuf[6585] = 256'h91d996dcb2df8fe209e5dce622e816e9c0e96dea54eb48ec61eda1ee9fef63f0;
    inBuf[6586] = 256'h0bf168f1d2f1baf231f4a6f655fae9fe4904160a6f0ff0133217951843188d16;
    inBuf[6587] = 256'ha5137210cd0d230c2c0c2f0ec811c8169b1c58229727db2b9c2e01302730222f;
    inBuf[6588] = 256'h992df42b632a5b29ee28f1287d29642a792bdb2c5a2ed72f7031e53214341735;
    inBuf[6589] = 256'hb135ca357a3599343f33af31f02f532e212d382cbb2baf2bad2bab2b942bfe2a;
    inBuf[6590] = 256'hf929912895265f242922e21fec1d5b1ce91ac319c91891173d16ad148a121d10;
    inBuf[6591] = 256'h760d720a8907df0459025700d1fe83fd9afcd8fbd9fabbf940f820f6aaf3dbf0;
    inBuf[6592] = 256'ha5ed75ea61e765e4d7e1b4dfe9ddabdccfdb2cdbe0daadda6bda39daead965d9;
    inBuf[6593] = 256'hccd8fed7f3d6c6d55fd4d6d257d1e4cfbfce23ce10ceb2ce12d0ecd122d46ed6;
    inBuf[6594] = 256'h64d8e4d9c1dad6da65da92d97bd899d717d7fbd69bd7e6d8a5daeedc82df0de2;
    inBuf[6595] = 256'ha3e408e7ffe8baea17ecf9ecbeed67eeedeeb6efb7f0caf133f3d2f474f64ff8;
    inBuf[6596] = 256'h39faf0fb9afd06fffbffbb0042017b01c5013302ac028203b004f8057207f108;
    inBuf[6597] = 256'h100adb0a3c0bfe0a650a99098a088d07ca0614069e0571053c051305fe04af04;
    inBuf[6598] = 256'h4104d60331037102b401b5008bff4cfeb3fcdefa01f9e4f6c3f4f3f24ff102f0;
    inBuf[6599] = 256'h4eefddee9bee87ee28ee61ed40ec77ea34e8d6e551e308e16fdf5adedbddffdd;
    inBuf[6600] = 256'h3dde62de67dee7ddfadcd9db60dad7d887d73dd629d568d498d3c8d20dd223d1;
    inBuf[6601] = 256'h50d0d1cf7ecf8ccf05d084d016d1a3d1c6d1a3d13cd156d051cf67ce8fcd3fcd;
    inBuf[6602] = 256'h91cd3cce5ccfb9d0dbd1dcd294d3c0d3bdd39bd355d379d31bd415d5aad691d8;
    inBuf[6603] = 256'h54da0cdc7bdd66de28dfbbdf10e091e02ae1c1e1ade2bbe3bce4f6e538e761e8;
    inBuf[6604] = 256'hcfe95febefecb8ee72f0e2f134f333f4def494f542f607f73ff8baf964fb64fd;
    inBuf[6605] = 256'h53fff0004302050336031e03cc029202c60255036b041406e907d309be0b480d;
    inBuf[6606] = 256'h770e780f51106111ec12eb147417341a861c201e881e481db11a22171613ae0f;
    inBuf[6607] = 256'hc70def0dc9102516471d73254b2d69331d37a237c234532f1b28302047195614;
    inBuf[6608] = 256'hfb11dd1293164b1c6b23a92aea30bd356438b13843374c344e30522c8e283b25;
    inBuf[6609] = 256'hf32297212021eb21aa233726b0296d2d123193342a377038883809370a344430;
    inBuf[6610] = 256'h002cde27b724ad22092206231025e0273f2b432e8330ea31f231b430a72ed82b;
    inBuf[6611] = 256'hc128e62543232621bb1fa61ef41d901df51c321c531b0f1ab7188c1765167e15;
    inBuf[6612] = 256'he7144414a013d9129711fd0f020e7b0bca0815065103f7002effcafdfefcadfc;
    inBuf[6613] = 256'h74fc53fc11fc67fb78fa34f98df7dff53cf499f23cf110f0d9eea6ed55ecc2ea;
    inBuf[6614] = 256'h20e983e706e6fce484e4a7e47ee5dbe672e805ea3debcdeb99eb91eac6e86ee6;
    inBuf[6615] = 256'hd7e35ce161df46de49de70dfa3e1abe419e894ebceee69f143f353f48ff439f4;
    inBuf[6616] = 256'h94f3b8f2f5f17cf12cf130f1aef186f2ecf308f6b4f804fce3ffeb03ff07d20b;
    inBuf[6617] = 256'hd70efa101b12f111d110160fee0cfe0ad2099509b10a360dc7103d15211ac41e;
    inBuf[6618] = 256'he62228262128fe28d528b42722266c24b2225e218e203c209a209221fd22e124;
    inBuf[6619] = 256'hf226f228e12a712c7c2d212e372eb92de22cb02b422ad4285727ec25b0247b23;
    inBuf[6620] = 256'h7422c2213421ed2004212f216b21aa21952127215a20f41e2d1d221bbb185216;
    inBuf[6621] = 256'h0e14ce11dd0f4f0edf0cb40bbd0aae09aa08a807730643051604c00280014e00;
    inBuf[6622] = 256'hf3fe97fd1bfc3bfa1ff8ccf537f3b9f078ee7bec09eb21eaa4e9a8e9fde95cea;
    inBuf[6623] = 256'hbceae7eaaaea15ea1fe9c7e738e687e4d5e25ce131e06bdf21df3adfacdf69e0;
    inBuf[6624] = 256'h47e138e222e3e2e37ce4ede42ee562e587e590e59ce5a3e5a1e5cae51ce683e6;
    inBuf[6625] = 256'h21e7dbe791e869e95aea54eb7eecbeedf5ee40f078f17bf271f339f4b5f427f5;
    inBuf[6626] = 256'h90f5eff590f676f781f8d4f94afba7fc04fe41ff2900e4006601850172013401;
    inBuf[6627] = 256'hb3002900abff25ffd4fecafee0fe48ff0600cf00ac01890203031503c502dc01;
    inBuf[6628] = 256'h8300e9fef7fcf2fa17f94bf7d1f5d9f41ff4b5f3a9f39af389f385f338f3adf2;
    inBuf[6629] = 256'h03f2f1f095ef20ee53ec59ea70e86ee692e422e3ece115e1b3e068e041e058e0;
    inBuf[6630] = 256'h55e050e065e03ee0ebdf8bdfd8def5ddf4dc8adbe3d926d834d683d473d3f0d2;
    inBuf[6631] = 256'h47d383d433d63dd85cdafadb09dd5adda6dc50dba0d9abd711d61cd5b4d424d5;
    inBuf[6632] = 256'h55d6e9d7ead90edce2dd7adfa1e019e142e12fe1d4e0a9e0b5e0d4e056e125e2;
    inBuf[6633] = 256'h11e366e403e6abe78de965ebdbec15eed5eeeeeebeee43ee92ed3ced5eedfced;
    inBuf[6634] = 256'h70ef83f1d4f350f684f80efafcfa1efb82fa9ef997f8adf76cf7d5f7d3f87bfa;
    inBuf[6635] = 256'h78fc6efe4200ab018602ef02db0277021d02cf01a601c101e101dc01b6015e01;
    inBuf[6636] = 256'hfb00cf00fe00c7013f0338059207ff09f30b1e0d440d440c7a0a66089306b405;
    inBuf[6637] = 256'h1e06c907990af00dfa102513cc139512e00f340c5d0895059a04c1053c09680e;
    inBuf[6638] = 256'h3c14d619021ecd1f0a1fb21b4b162a10620af8050904c404ce07c70ca3124218;
    inBuf[6639] = 256'h0d1d452098216d21f71fa91d681b7319e4171c17da16d4163a17e317c918461a;
    inBuf[6640] = 256'h381c851e52212a24b226ea285a2ab92a422ae528d726c424f422c621b1218a22;
    inBuf[6641] = 256'h2a247c26e9280d2bcb2caf2d9a2dcf2c4a2b5d298a27df259924f023a323ad23;
    inBuf[6642] = 256'h0e2463249924ac244f249f23cb22b12189207a1f4b1e1e1d0f1ce71acb19c518;
    inBuf[6643] = 256'h8d173f16e2144613b0114410d60e980d990c9d0bc80a1a0a4d096a085607c805;
    inBuf[6644] = 256'hf203f001b0ff87fd98fbbff926f8def6bdf5def43af496f3f6f253f28cf1d0f0;
    inBuf[6645] = 256'h45f0d7ef9cef94ef80ef48efdcee0deed5ec4aeb79e9a6e741e692e5e4e56ce7;
    inBuf[6646] = 256'hf6e918ed6ef06cf396f5cbf6f8f62ef6d3f444f3daf126f16bf19af2b8f46bf7;
    inBuf[6647] = 256'h1cfa92fc97fef1ffdf0094012102eb021e04ab05bd07310a900cb90e6f105e11;
    inBuf[6648] = 256'hbe11c21185117811d8119d120314f41519185f1a801c1b1e401fef1f28203820;
    inBuf[6649] = 256'h3a202f2051209620ea206921f3215d22b422e022de22dc22d822e12217235323;
    inBuf[6650] = 256'h9023da23fb23e5239b23f022f521ce20751f261e081dfc1b2a1b991a131ab019;
    inBuf[6651] = 256'h6c1904198e180318311748164615f5137912bd108b0e2c0cbf09470728057e03;
    inBuf[6652] = 256'h22024401c5005e002900fcff8cfff5fe15febffc33fb72f96af758f530f3d8f0;
    inBuf[6653] = 256'h9cee90eccaeaa4e921e924e9b0e983ea5aeb25ec9cec89ece2eb84ea85e842e6;
    inBuf[6654] = 256'h03e427e203e196e0d1e08ee17ee279e35be4efe43be549e520e50de541e5c1e5;
    inBuf[6655] = 256'ha9e6cce7d5e8abe920ea0eeaaae903e92ae87be712e705e7a5e7e1e885ea9bec;
    inBuf[6656] = 256'he1ee05f110f3def445f676f75bf8e0f842f977f971f974f970f943f92ff932f9;
    inBuf[6657] = 256'h41f9b1f996fad3fb8bfd8bff6d0116033a0482041104f7023f0166ffc5fd7cfc;
    inBuf[6658] = 256'heefb34fc05fd4ffec7ffe200760163016900c6fec8fc8bfa7ff8fff6faf595f5;
    inBuf[6659] = 256'hcaf529f693f6eaf6c3f622f627f5acf3ebf134f078eeefeccbebd4ea1feac1e9;
    inBuf[6660] = 256'h70e938e92fe9fae89ce829e857e73de60be594e307e29ce031dffedd34dd95dc;
    inBuf[6661] = 256'h3adc26dcfddbd1dbbbdb83db5edb72db81dba7dbe5dbe6dbc1db79dbd6da16da;
    inBuf[6662] = 256'h61d9a1d831d839d889d84fd973da89db97dc7cddf3dd41de81dea3def5de72df;
    inBuf[6663] = 256'hd4df47e0b3e0e4e028e182e1cbe153e222e31fe49be587e78ee9a9eb77ed91ee;
    inBuf[6664] = 256'h27ef43eff5eeb2ee8bee68ee90eefaee8aef79f09af19bf288f349f4e3f4c9f5;
    inBuf[6665] = 256'h25f7e5f802fb06fd74fe3fff4aff99fe8efd4ffcf8faedf96cf9a4f9c6fa9efc;
    inBuf[6666] = 256'hc5fedd0072025803bb03b1035703d8022c025c01a1002e003800d100ce011003;
    inBuf[6667] = 256'h6e04b905fa062208eb082c09c0089e072206b904bb0384030d04190596063b08;
    inBuf[6668] = 256'ha909c30a2f0b940a2609320732050204160477052f08c00b890f3d133b16d717;
    inBuf[6669] = 256'he9172c16b912860e720a3d07cf0545064308a60be40f5b14c9187d1cd01ecb1f;
    inBuf[6670] = 256'h681f041ea61cc41b701bea1bd21cc41df21e42208421d022c7233924a4244025;
    inBuf[6671] = 256'h522645289a2a942ced2d3c2e882d762c422b0d2a26296f281b28b528312a582c;
    inBuf[6672] = 256'hd92ebb3066310331ba2f162ec02ca32ba52ad329fe286c287528c62817291729;
    inBuf[6673] = 256'h33289926e52450232d228c21d420d01f9d1e391d051c2f1b451a181993178d15;
    inBuf[6674] = 256'h8a130312c810c20fb30e210d400b87091e084207ca061506fd049603eb017a00;
    inBuf[6675] = 256'h7dff88fe65fdeefbf6f9dcf710f697f47af3a6f2eaf189f1e8f11bf316f571f7;
    inBuf[6676] = 256'h57f93bfaf2f968f8e1f5c3f232ef79eb35e807e693e55ae729eb40f0b4f584fa;
    inBuf[6677] = 256'h00fe02008400a1ffb3fd03fbf7f763f5e7f3c0f30af55ef705faa7fc1fff6501;
    inBuf[6678] = 256'hb8031e065808540ae70bf30cbe0d5c0e910e5f0eb80d970c7f0b010b710b100d;
    inBuf[6679] = 256'hb60ff7128d16201a531d0120c92141226e217f1fe31c621a8d18ab17d917e718;
    inBuf[6680] = 256'ha31af31c951f4522b0245226f226a226892509247622c820001f1f1d2e1b8c19;
    inBuf[6681] = 256'h88182c188a185e193b1a1a1bdf1b421c451cb21b371a0b187a15d2129e10ec0e;
    inBuf[6682] = 256'h750d290cbb0a00095807d5054f04eb028301f3ff9bfea3fd02fdbdfc5efc6ffb;
    inBuf[6683] = 256'hfdf9fef79df55df33af112ef11ed2ceb78e952e8aee74ce701e75fe64ce516e4;
    inBuf[6684] = 256'he4e2f5e182e146e113e1ece09ee02de0a9dfc7de71ddb4db99d992d712d635d5;
    inBuf[6685] = 256'h22d5bfd5acd6e8d766d9ecda7ddcdcdd93de98dee8dd96dc2edb00da1cd9d0d8;
    inBuf[6686] = 256'h09d98ed999da17dcc8ddcbdfe7e1c2e37ce5fae60be8ece87be985e94de9d2e8;
    inBuf[6687] = 256'h0fe87de736e731e7cee709e9b3eafceca5ef36f29ef484f693f70df80bf891f7;
    inBuf[6688] = 256'h0bf786f6e1f563f510f5d3f4fff48ff540f62af729f8f3f8c2f9aafa8ffba6fc;
    inBuf[6689] = 256'hd8fdcffe80ffbfff43ff33fea3fc8afa4df846f69ef4c8f3f7f3edf47ff64df8;
    inBuf[6690] = 256'hc6f9c6fa46fb2afba6facef976f8c7f6f6f421f3b2f1e8f098f0aef0fbf02cf1;
    inBuf[6691] = 256'h48f15ff13ff1dcf012f0aaeed6ece9ea1ee9d2e71be7bde6bde620e7d3e7fee8;
    inBuf[6692] = 256'h8eea0dec26ed8eed0eede8eb64eaa2e8e0e62ae57ee340e2bbe100e22ee3fde4;
    inBuf[6693] = 256'he0e6a1e81cea3ceb38ec0eed89edaeed70edd3ec38ecc4eb5deb0eebb3ea31ea;
    inBuf[6694] = 256'he4e911ead1ea44ec23eef9efaaf119f33ff45df568f626f798f7a6f752f7fff6;
    inBuf[6695] = 256'hdcf6e6f638f7aaf70bf876f8ecf852f9aaf9c1f977f905f9a6f8a2f851f99dfa;
    inBuf[6696] = 256'h32fcdafd4eff6000250197019101ff00cdff24fe68fcf0fa01fab2f9c3f903fa;
    inBuf[6697] = 256'h6bfa04fbf6fb5bfd0fffe0009002f3031605f3055c062c0623051a036d00a3fd;
    inBuf[6698] = 256'h4cfb0cfa22fa71fbdbfdf70043046e07e5091f0b190be809ea070806e204be04;
    inBuf[6699] = 256'he2050808ac0a990d58106f12cc131f144313c011f20f430e730da30d9c0e7310;
    inBuf[6700] = 256'hd21262155118681b561e25216c23d024842568256e24072337210f1f321dda1b;
    inBuf[6701] = 256'h451b011cfa1deb20d3241e29412d0e31de333135153561335530d52c60297e26;
    inBuf[6702] = 256'hd8245524cc2437260728db299b2bce2c542d792d1e2d6f2cbc2bc12a73290e28;
    inBuf[6703] = 256'h7a26ff2405245f230123dd228222002299212021a62025201a1f7f1d941b6219;
    inBuf[6704] = 256'h5d17d7158b147c13a912cd111f11c3105110a40f920ec50c8a0a510833067804;
    inBuf[6705] = 256'h1b03b801630046ff59fee5fde9fde1fd92fddafc8cfbfbf979f803f7b1f583f4;
    inBuf[6706] = 256'h55f362f2e4f1d3f136f2d6f23af32cf3a5f297f13af0d4ee82ed7dec07ec3fec;
    inBuf[6707] = 256'h37edddeecff099f2ddf34af4d5f3c2f255f1d1ef91eed0edb2ed70ee23f0a3f2;
    inBuf[6708] = 256'hb4f5f1f8d8fb20feaaff7300c000c900a10078006b006d00a4002801d701aa02;
    inBuf[6709] = 256'h990382048105c4065808510a930cc70eab100812b412d712b41281128b120313;
    inBuf[6710] = 256'he7132a15a016ff17081986195d19a41894177a16aa155815991561168c17fb18;
    inBuf[6711] = 256'h801ae71bfc1c731dfc1c8f1b441963167813e410c80e300de90bc50ae7097209;
    inBuf[6712] = 256'h9109760ae40b660db10e550f080fe70dec0b14099f05aa0170fd7af912f66df3;
    inBuf[6713] = 256'hd4f123f127f1d4f1d4f2c6f37df495f4e4f3a2f2fbf045efe7edd0ecd8ebedea;
    inBuf[6714] = 256'hc5e959e8f2e6a4e590e4d4e335e393e2e5e106e11be061dfdedec4de37df0fe0;
    inBuf[6715] = 256'h49e1d5e262e4dae517e7c9e7e5e75be70ce642e443e242e0b5ded5dd92dd0fde;
    inBuf[6716] = 256'h30dfb3e0a6e2e6e423e75fe960ebdeecfbeda6eebfee82eee3edc7ec8feb76ea;
    inBuf[6717] = 256'hace9bee9d7eacbec98efd1f2eaf5b2f8ccfae9fb35fcb2fb6dfaeaf869f702f6;
    inBuf[6718] = 256'h1bf5bef4c4f457f567f6bdf768f937fbd4fc3bfe48ffcfff09000200a1ff1aff;
    inBuf[6719] = 256'h73fe91fdb7fc10fc99fb87fbe3fb6cfc17fdc1fd2ffe79feb8fee4fe28ff84ff;
    inBuf[6720] = 256'ha7ff6fffb5fe3cfd31fbecf8a4f6b8f46cf3b0f283f2dbf283f37df4c1f509f7;
    inBuf[6721] = 256'h38f829f984f942f981f83ff7b5f529f49df220f1bbef3aee95ecd5ea02e96de7;
    inBuf[6722] = 256'h7de662e659e75fe902ecdfee8bf17ff383f487f464f335f12fee89eac3e665e3;
    inBuf[6723] = 256'hc8e04bdf04dfb3df3de175e30fe6fae80eece4ee3bf1cff25df303f3e7f132f0;
    inBuf[6724] = 256'h3bee2eec14ea41e8f4e650e6b2e632e894ea9deddcf0c5f30ef672f7cdf749f7;
    inBuf[6725] = 256'h00f61cf411f22bf0a9eef9ed48ee8fefd9f1f0f470f807fc3aff8b01ba029102;
    inBuf[6726] = 256'h1d01c2fedefbe0f84ff66ff46bf37ef3a9f4d6f6e8f981fd2a017204df063208;
    inBuf[6727] = 256'h69089407fe05fd03bd0178ff65fd9cfb5dfaf5f992fa67fc5fff0f030007880a;
    inBuf[6728] = 256'h040d4a0e620e800d2f0cd00a84097b08b0070d07c606e9066f076c089a099a0a;
    inBuf[6729] = 256'h630bd40bec0b230cb00ca20d3c0f4e1171137f15041791173917fa1516144f12;
    inBuf[6730] = 256'h0a1184100e114f12cd137e1514176818cb19291b591c861d7d1e241fcc1f5620;
    inBuf[6731] = 256'hab20fc200621a4202b20931fea1e961e7e1e911e141fdb1fd120232277238824;
    inBuf[6732] = 256'h6225a8254225862464230422dc20e81f481f521fdc1fd6205c220d24b7255227;
    inBuf[6733] = 256'h6628c6287b2838271b2586227b1f491c6919de16ee14fe130014041503176c19;
    inBuf[6734] = 256'hde1b071e591fc11f571fe61d961ba91817154411b80da10a550805076c067a06;
    inBuf[6735] = 256'h250722087209090b790c940d3c0e310e900d8a0c000bf0084f06ed0208ff22fb;
    inBuf[6736] = 256'habf741f54cf4aff438f692f82afba9fddeff7c016e02c1025902370171fffdfc;
    inBuf[6737] = 256'h00fadff60cf41ef2a1f1aef208f529f846fbbbfd49ffdcff97ffd6fed0fda9fc;
    inBuf[6738] = 256'hb0fb1ffb1bfbcffb24fdc7fe7000cc019e02f102d7026a02f601b701dd01a602;
    inBuf[6739] = 256'h1004d00596070109cd091e0a3e0a740a000bd80bb90c7d0d0b0e660eba0e130f;
    inBuf[6740] = 256'h4e0f470fdb0e050efe0c130c870b820bfe0be30c0e0e560f9710a81155127712;
    inBuf[6741] = 256'hfd11f310860fee0d5f0c110b170a790947096309ac09130a690a880a730a0a0a;
    inBuf[6742] = 256'h370905086406650451025700affe91fddcfc61fc02fc80fbd8fa48fad9f997f9;
    inBuf[6743] = 256'h88f952f9b1f89df702f616f43ef293f033ef32ee57ed98ec11ecadeb81ebabeb;
    inBuf[6744] = 256'hfdeb67ecdbec0aedd7ec34ecfcea6de9e9e7a8e6f7e5dde5ede5d9e574e5ade4;
    inBuf[6745] = 256'hf4e3c4e33ee461e5c9e6d5e755e850e8f4e7bde7d8e707e82ee81ae8ade756e7;
    inBuf[6746] = 256'h74e723e880e936ebb5ecc3ed2eeee9ed56edb1ec20ec07ec82ec7eed15effff0;
    inBuf[6747] = 256'hccf263f49cf568f622f7dff771f8cbf89bf8aaf758f60ef539f462f489f54bf7;
    inBuf[6748] = 256'h69f97efb30fd91fe8ffffaffe9ff61ff79feacfd47fd4bfdbffd4cfe72fe26fe;
    inBuf[6749] = 256'h76fd77fc96fb10fbd4faf8fa77fb1dfcf0fcd6fd7dfed2febffe1dfe2bfd21fc;
    inBuf[6750] = 256'hf9fae6f905f92af871f7eff66ff6f1f572f5b6f4ddf316f358f2d1f194f15bf1;
    inBuf[6751] = 256'h1ff1e9f099f066f08bf0ebf086f137f27df221f210f125efb9ec49ea1ae89fe6;
    inBuf[6752] = 256'h1ee66de67fe72ce9fdeab6ec1eeec9eea6eecfed50ec93ea01e9bae7fee6d0e6;
    inBuf[6753] = 256'heae640e7b3e7fde73ce896e80ee9eae942ebc8ec3bee37ef58efc1eec0eda9ec;
    inBuf[6754] = 256'hf5ebb0eb86eb48ebcaea0cea8fe9bde9c0eab2ec3cefd2f122f4c8f571f626f6;
    inBuf[6755] = 256'hedf4f2f2c6f0e5eeb4ed91ed5ceebcef76f131f3b8f426f665f763f838f9d4f9;
    inBuf[6756] = 256'h4afadbfa7ffb16fc83fc67fc90fb27fa58f879f6fcf40cf4daf398f441f6d3f8;
    inBuf[6757] = 256'h26fca3ffb702e504bb054b05110487024601b900e300b201eb0222042105ba05;
    inBuf[6758] = 256'hbb054d05ad04fe039803a4031204ff046d063f08860a050d3b0fda108b112a11;
    inBuf[6759] = 256'h2b10ff0ef60d6a0d3e0d1f0d110d100d2d0dc70dd90e2a10b41130136f14aa15;
    inBuf[6760] = 256'hca169f174a189f1886185c1833180a18151831184e18c21883196f1a7d1b101c;
    inBuf[6761] = 256'hb41ba71a2d19e317b817d218de1a771dc41f3f2114224e222b221222c8211e21;
    inBuf[6762] = 256'h4020121fbb1db11cec1b661b481b501b741bf01b961c641d871eb31fcd20ee21;
    inBuf[6763] = 256'hb222dd2270221e21fd1e901c1c1a1e181117cf162f170118ab18f418e5184718;
    inBuf[6764] = 256'h42172c16f814d41301135212c2116011e91068100610a90f730f800f810f5b0f;
    inBuf[6765] = 256'h030f270ed60c500b9c090408d706fd0578053205c90429046a038802d701b401;
    inBuf[6766] = 256'h0d02d102d2039404de04b20403040703f701ca009dff99febbfd36fd33fd7dfd;
    inBuf[6767] = 256'hddfd28fe16feb4fd60fd5afddefd03ff7500d801f1028703a303760308036a02;
    inBuf[6768] = 256'hbd01040163001c003700ab006b013a02fa02be038904620551062307a507d407;
    inBuf[6769] = 256'hb50773075a0789070708ce08b0098c0a520be00b1e0cfe0b680b6e0a47093008;
    inBuf[6770] = 256'h7a076307ef070309670ac80be70c970dbd0d6e0dcf0c130c870b490b4e0b750b;
    inBuf[6771] = 256'h630bbe0a7509a1079b05f903220340034a04ce0543075408b6086308a307a206;
    inBuf[6772] = 256'h89058d049b03a102b401b40097ff7dfe44fde4fb92fa57f95df8f4f712f894f8;
    inBuf[6773] = 256'h50f9cdf9b7f904f99ef7bff5d3f300f279f075efd5ee93eebdee1bef93ef18f0;
    inBuf[6774] = 256'h56f02cf0a2ef98ee3deddbeb85ea67e99be8f7e777e720e7dce6d5e62be7bde7;
    inBuf[6775] = 256'h8ae870e915ea68ea5beacde9ece8dde7a3e680e598e4e5e393e3a5e3f6e3a7e4;
    inBuf[6776] = 256'hb7e50ae7bee8a9ea74ecfeedfaee27efbbeedfedbcecbeeb0eeba9eac5ea61eb;
    inBuf[6777] = 256'h65eceaedb2ef4ff196f238f312f38ff205f2b8f1fff1b9f28bf366f424f5c0f5;
    inBuf[6778] = 256'h97f6b2f7d8f8f2f9b0facdfa90fa48fa33faacfaa8fbcdfcf1fdc6fe13ff01ff;
    inBuf[6779] = 256'h9cfedbfdf6fc02fc02fb4afa11fa63fa6ffb24fd2cff58014e039004f7047004;
    inBuf[6780] = 256'hf602f100d9fefbfcaafbfbfaacfa9dfab2facafa12fbadfb77fc60fd3dfebafe;
    inBuf[6781] = 256'hd8feb6fe51fecdfd31fd3ffcf0fa63f9b4f750f6a4f5bdf594f6e5f721f9eef9;
    inBuf[6782] = 256'h17fa72f93bf8b9f60af575f330f23bf1c7f002f1d3f12ef3d1f42ff6edf6ccf6;
    inBuf[6783] = 256'habf5e4f3f0f124f0e8ee61ee5deebbee41ef9aefb5ef86ef09ef8fee59ee7dee;
    inBuf[6784] = 256'h1def0cf0e1f065f177f114f191f02ff0faeffeef05f0d0ef68efd5ee27ee9aed;
    inBuf[6785] = 256'h40ed25ed88ed84ee2af085f23ff5d9f7f9f943fb9efb45fb6bfa3bf9e4f768f6;
    inBuf[6786] = 256'heaf4b1f3e6f2c1f25af379f4f1f5abf781f97bfba0fdbaff9f011e03fe035304;
    inBuf[6787] = 256'h4304d5033b038c02c4012001d600fa00ba01000382043406f4079709440bdf0c;
    inBuf[6788] = 256'h200efa0e460fe80e340e600d8a0c080ce40b100cd30c290ef20f36128c146f16;
    inBuf[6789] = 256'hc1173e18db171b1740167b1542158d152e1641178018a219b81a851bec1b3c1c;
    inBuf[6790] = 256'h701c971c111dbc1d6e1e4d1f12208b20e8200121ca2091204120ea1fec1f3020;
    inBuf[6791] = 256'hae2097219622642307242c24bf2313233222612117214721ef211a2342241025;
    inBuf[6792] = 256'h75251725fc238a22d820371f161e601d0e1d211d301d1f1d0d1ddd1cc41c091d;
    inBuf[6793] = 256'h721ded1d641e5f1ec11da51ce81abc187d1635143012c010d00f6d0f8c0fc00f;
    inBuf[6794] = 256'he70f0310da0f900f4b0fd10e160e1c0db30b160aa1087607de06eb0634077507;
    inBuf[6795] = 256'h6e07b9066505b903d8011700c7fee9fd8ffdbbfd35fee9febcff6800da000c01;
    inBuf[6796] = 256'hcf002a003afff7fd89fc35fb1efa6cf93ef973f9e2f96efaf2fa71fb04fca4fc;
    inBuf[6797] = 256'h43fdc3fdf0fdb4fd29fd74fcc9fb58fb2bfb2ffb58fb97fbe6fb4efccdfc51fd;
    inBuf[6798] = 256'hc8fd1ffe45fe45fe38fe2bfe3afe7dfeeefe7cff15008f00c300ac005700e3ff;
    inBuf[6799] = 256'h83ff57ff62ff9bffe8ff34008700e00037018701ae0183010e016c00b7ff2aff;
    inBuf[6800] = 256'he7feddfe00ff40ff74ff95ff9dff6cff06ff7efedbfd51fd15fd18fd47fd7ffd;
    inBuf[6801] = 256'h72fd0dfd6afc91fbb1faf3f93df995f80df889f71df7e7f6bcf692f678f64df6;
    inBuf[6802] = 256'h21f612f6f2f5a4f517f512f4b4f252f113f03feffceef8eef5eec8ee24ee2bed;
    inBuf[6803] = 256'h27ec26eb5aeadde96fe90fe9d8e8b8e8dbe85fe900ea9cea0aebf3ea67ea8de9;
    inBuf[6804] = 256'h57e803e7c2e583e491e32be340e3ece30be516e6e1e645e70ae772e6aee5a8e4;
    inBuf[6805] = 256'h98e3a2e2c5e16ae1c8e1b2e21ce49ee59fe619e71de7aee642e6fce5a1e54fe5;
    inBuf[6806] = 256'h0be5c9e4f4e4ace5a6e6cae7b1e8e5e8a2e826e89ae77fe7ebe79fe8ace9e0ea;
    inBuf[6807] = 256'he9ebd9ec7aed79ed11ed67ec9feb4beb95eb3eec35ed1bee8aeeaeee9dee5dee;
    inBuf[6808] = 256'h42ee51ee6beed9eeb5eff6f0ccf2f4f4ecf679f83df9f3f8e3f747f652f48df2;
    inBuf[6809] = 256'h44f18af09bf05df17ef2e0f341f56bf685f795f892f9a0faa5fb6afcf4fc28fd;
    inBuf[6810] = 256'hdbfc26fc0efba3f946f846f7d5f633f740f898f9f1faf5fb67fc6cfc39fc01fc;
    inBuf[6811] = 256'h0dfc73fc18fde7fda7fe0fff0eff95fea1fd68fc17fbc5f9a5f8d9f771f79cf7;
    inBuf[6812] = 256'h6ef8ccf992fb7afd20ff4f00ee00f2006f0077ff08fe41fc4afa5af8c9f6d1f5;
    inBuf[6813] = 256'h75f5b0f565f663f7a1f81ffabefb50fd94fe39ff15ff23fe7efc6cfa3df835f6;
    inBuf[6814] = 256'hadf4edf314f415f5adf66af8e0f9ccfa2ffb44fb44fb51fb60fb42fbd9fa38fa;
    inBuf[6815] = 256'h9df95bf99ff952fa2efbcbfbddfb6efbbafa13fae0f943fa22fb66fcdcfd4cff;
    inBuf[6816] = 256'hb100f501e902800395030b031402d40081ff8afe24fe62fe7dff550194031406;
    inBuf[6817] = 256'h78085d0ad20bdd0c870d240eab0ee70ef20eab0e120ea80da20dfc0ddb0ee40f;
    inBuf[6818] = 256'ha61038119c11f711d6123e14f5150218fd19971b151d6b1e791f752017210e21;
    inBuf[6819] = 256'h9020961f411e291d7a1c551c271dc71ef320a3233426152845298129e6282228;
    inBuf[6820] = 256'h6827d826cb26fb263827b8273d28ad282f2965293129ec288d284e28a5284c29;
    inBuf[6821] = 256'h072ad22a372b1b2bd12a302a4e2972285b271b26142521245c230623c1227b22;
    inBuf[6822] = 256'h62222d22ed21d92197211b218420801f2d1ee11c761b241a42199c1849186f18;
    inBuf[6823] = 256'h9e18aa188c18d8179c1625156a13b31157102c0f4f0ee80daa0d980dc00db90d;
    inBuf[6824] = 256'h6d0de70cdc0b5f0ab208c306d1043803000266019b015a027403bb04b6054806;
    inBuf[6825] = 256'h8d066906f9055e056d042b03d00171005affd3febefef5fe45ff56ff19ffbdfe;
    inBuf[6826] = 256'h57fe16fe20fe57fea4fe06ff6dffe2ff74001401b1013b029002ab0293024202;
    inBuf[6827] = 256'hcf016001100104015b010402ce027903cc03ae0332039702280210025a02fb02;
    inBuf[6828] = 256'hc9039c04640509066c066906d505a70408034501d4ff27ff66ff890054025404;
    inBuf[6829] = 256'h23068a0759088e0847088c0779062c05a303fd016600ebfebbfd0dfdd7fc15fd;
    inBuf[6830] = 256'hc4fda7fe94ff750009012001990042ff37fdd1fa67f87ff685f564f5f3f5f2f6;
    inBuf[6831] = 256'he1f785f8e0f8d2f86ef8d2f7edf6def5cff4b2f3a1f2a4f186f05bef57ee80ed;
    inBuf[6832] = 256'h1aed4cedcfed73ee04ef20efc8ee14eeeeec84eb04ea6be81be771e66ce61ee7;
    inBuf[6833] = 256'h4ce847e9b8e97ee987e85be77ce60ae634e6d4e66ce7f0e759e879e88ae89ce8;
    inBuf[6834] = 256'h5de8dce728e729e642e5bfe491e4dce47ce5fbe556e67ee649e614e616e62ee6;
    inBuf[6835] = 256'h8fe62de7a5e708e852e84ce83ce843e83ee86ae8cce824e995e914ea5feaa5ea;
    inBuf[6836] = 256'heeea0beb2deb4ceb1debbeea34ea66e9bfe87de899e852e98eeaf2eb82ed10ef;
    inBuf[6837] = 256'h43f01ff174f1f2f0d0ef49ee9fec75eb20eb90ebc2ec50eebbeff7f0ecf18bf2;
    inBuf[6838] = 256'h25f3c6f341f4aff4eff4c8f465f4d3f316f37cf218f2dcf1e9f11df24ff2a8f2;
    inBuf[6839] = 256'h2cf3d5f3d5f411f649f77bf883f944faeefa7cfbc1fbb9fb35fb18faaff846f7;
    inBuf[6840] = 256'h2af6c8f530f637f7c7f89bfa63fc0efe68ff30005e00dfffaefe13fd45fb75f9;
    inBuf[6841] = 256'hfbf702f79ef602f72cf8e5f9fefb22fee7ff2701d501ed019901ed00e1ff8efe;
    inBuf[6842] = 256'h08fd70fb16fa31f9c1f8c0f8fff834f951f96ff9a6f927fa06fb15fc1afdd6fd;
    inBuf[6843] = 256'h0cfeb4fdedfcd5fba0fa75f962f87ef7e3f69cf6bbf647f724f82df937fa14fb;
    inBuf[6844] = 256'ha8fbedfbecfbb4fb53fbcefa1efa3df929f8eaf696f55cf460f3cff2dbf299f3;
    inBuf[6845] = 256'h02f50ff785f90efc69fe4c007c01f601b801c9005dff9afdb1fb0ffa00f9b2f8;
    inBuf[6846] = 256'h5cf9d6fabcfccefeb00018022603f00382041d05bd0538069b06ce06b3068606;
    inBuf[6847] = 256'h5b0634065806d2069707e408b10acb0c340f99118e13111508167716c7161917;
    inBuf[6848] = 256'h5e17b717ec17c51779171217a2168016aa160d17e3171f19b31ac91c191f4521;
    inBuf[6849] = 256'h30237624e524c0240924de22ab218120881f311f7e1f6220e2218523e6240426;
    inBuf[6850] = 256'had26fb264c277c2771272c275326e42445238721e11f9f1e801d6d1c991bf61a;
    inBuf[6851] = 256'hbd1a491b631cdb1d871fd3208521a821f620741f571d7c1a2217d213c5106c0e;
    inBuf[6852] = 256'h3a0d080dc20d510f2611eb126c142115dd14bf13ba11210f6e0caf091107c004;
    inBuf[6853] = 256'h8e029a0032ff5ffe56fe3cffb8007f024e049f0545065106b40598044003a901;
    inBuf[6854] = 256'he9ff2cfe76fcfbfa00fa93f9c3f987fa8dfb98fc8efd3bfe96feb2fe75fecefd;
    inBuf[6855] = 256'hd0fc84fb20faf9f848f835f8cdf8e9f959fbf5fc80fec3ff9700d5007f00d0ff;
    inBuf[6856] = 256'h1effc4fe01ffcbffde00e0018402ac0274020b02a2015b0144016601cf018702;
    inBuf[6857] = 256'h7f038b047005f7050606b3052e059a041404a503490312032903a5038904ac05;
    inBuf[6858] = 256'hc706a0071b083e0830080d08bc0725073906fb04ad03ac022b023502a5021b03;
    inBuf[6859] = 256'h4d031f038402a401b300c1fff0fe62fe18fe24fe88fe09ff74ff9cff45ff6ffe;
    inBuf[6860] = 256'h3efdb9fb0efa72f8f4f6d5f55af582f54ef692f7caf8a1f9e6f967f94ef8e2f6;
    inBuf[6861] = 256'h34f57bf3e4f162f01fef3bee8ded22edf8ecd4ecdcec3deddaedcbee03f019f1;
    inBuf[6862] = 256'heef170f261f2e1f10bf1b2ef08ee3fec5dead7e80ce8eee79de8fde988eb12ed;
    inBuf[6863] = 256'h6cee2fef6def38ef72ee6eed73ec7aebd2ea93ea7aeaa1ea08eb6bebeeeb91ec;
    inBuf[6864] = 256'hffec48ed6eed4bed39ed74ede3eda5ee8bef0cf01ef0bcefd4eedaed1ded88ec;
    inBuf[6865] = 256'h41ec32ec04ecd6ebbbeba6ebe4eb84ec4ced4cee5aef18f097f0ccf089f013f0;
    inBuf[6866] = 256'h8befe4ee5beefdeda9ed97edd2ed44ee12ef0cf0caf02bf1f6f008f0c9ee97ed;
    inBuf[6867] = 256'hb1ec84ec13ed20ee94ef25f181f2a2f358f469f4eff3e6f25af1baef52ee5fed;
    inBuf[6868] = 256'h41ed09ee8cefadf107f428f6d9f7d9f80df9b4f8f4f7f0f6f5f50ff536f491f3;
    inBuf[6869] = 256'h25f3ecf208f371f30ef4e4f4e4f504f75ef8e1f962fbbffca9fde1fd6cfd69fc;
    inBuf[6870] = 256'h13fbd2f9ecf87ef899f827f9fbf9fcfa07fcf9fcc7fd67fed0fe14ff3eff4bff;
    inBuf[6871] = 256'h3dff0dffb0fe30fea3fd20fdc1fc94fc96fcc1fc0cfd6afdd2fd3afe94fed8fe;
    inBuf[6872] = 256'h13ff59ffbeff54000e01b9011b0206025d013b00e6feaafdcdfc81fcbcfc54fd;
    inBuf[6873] = 256'h16feb9fe11ff1affdffe89fe57fe62feb5fe54ff1000bb00440182015d01e700;
    inBuf[6874] = 256'h1d0011ff0bfe3dfdd7fc19fdf3fd37ffc0003f02760376043405b10515064306;
    inBuf[6875] = 256'h0e067e057e041603b10195000c008100ef011c04e006bf09420c600eed0fd710;
    inBuf[6876] = 256'h5c116311c710af0f190e2b0c850a820965098d0abe0c940fe81241163b19dd1b;
    inBuf[6877] = 256'hd81deb1e3d1fb21e551daf1bfd198418d517f317cf18841aa41cc41edd209022;
    inBuf[6878] = 256'hbf23c52496252d26c9261a27ee268526cc25ee246f2439243c24a22413257625;
    inBuf[6879] = 256'h1f26ef26df271a292c2ac72a012b9a2ab629da28fa2726279726ea2503252c24;
    inBuf[6880] = 256'h4723802244225b22b2225f23ec2330244b24eb2314230c22a9200c1f931d161c;
    inBuf[6881] = 256'hb21aaf19d1181f18cc1786173417eb1653167915b014f3137d139013d1130914;
    inBuf[6882] = 256'h1314741322125d10210eb50b77095e079f058b041b047504ae0552070109620a;
    inBuf[6883] = 256'he60a710a3c09670751055a038401f3ffd0fe12fee6fd6afe66ffa900f801ef02;
    inBuf[6884] = 256'h7b03b803ae0385035103e6022f022a01ceff50fef4fce2fb4efb53fbe2fbeffc;
    inBuf[6885] = 256'h57fed6ff3b015c0214036c037b034803e102430266015d0055ff84fe20fe3cfe;
    inBuf[6886] = 256'hbbfe6fff2500c3005301e90192023e03bd03e3039f03fd0230026f01cb004000;
    inBuf[6887] = 256'hb1fff6fe13fe1ffd43fcb8fba1fbfcfbc3fcd2fde6fed0ff5d006200eaff0fff;
    inBuf[6888] = 256'he7fda6fc66fb28fa0df932f89ff777f7b0f70df86af89df87ff830f8c8f73df7;
    inBuf[6889] = 256'h9df6dbf5d5f4b1f39df2a9f109f1c4f0a5f0a7f0b9f0aff0a0f08cf04af0f2ef;
    inBuf[6890] = 256'h96ef22efc8ee98ee67ee3fee1feee0edaeed9bed79ed50ed12ed8becf4eb85eb;
    inBuf[6891] = 256'h33eb27eb4feb49eb12ebb9ea33ead7e9cfe9dbe9f4e9f7e9a0e92fe9e6e8c1e8;
    inBuf[6892] = 256'hfae888e90aea82eaf1ea25eb5debb0ebe3eb12ec3fec29ecfaebbfeb3beb99ea;
    inBuf[6893] = 256'hf2e926e984e835e80ae826e882e8d7e851e9ffe9a4ea5aeb09ec52ec57ec33ec;
    inBuf[6894] = 256'hd1eb85eb6deb45eb1eebe8ea63ead6e970e920e92de99ee927eadaeaa3eb38ec;
    inBuf[6895] = 256'hc2ec44ed84eda7eda3ed35ed8cecc0ebccea18eadbe9f8e98dea6beb22ecaaec;
    inBuf[6896] = 256'hefecccec90ec6aec49ec6decdaec5ded1bee0cefebefc2f06bf194f15af1d2f0;
    inBuf[6897] = 256'hffef42efc8ee71ee50ee44ee0ceed1edb7edc5ed46ee4bef9af02ff2dbf346f5;
    inBuf[6898] = 256'h68f620f730f7b4f6c9f575f411f3d7f1c6f012f0ceefedefa5f009f2e6f31ff6;
    inBuf[6899] = 256'h62f835fa73fb0dfcf1fb52fb49fac4f8f0f603f531f3f3f199f11cf265f327f5;
    inBuf[6900] = 256'hebf68cf801fa3cfb61fc6efd2cfe83fe5cfe9ffd7efc2efbcdf997f8b1f714f7;
    inBuf[6901] = 256'hdcf60bf781f73ef82ef926fa1ffb03fca9fc0bfd1cfdd1fc4dfcb2fb16fba7fa;
    inBuf[6902] = 256'h72fa70faa9fa12fb98fb38fcd9fc65fdd7fd20fe3bfe35fe09fec1fd7cfd49fd;
    inBuf[6903] = 256'h3bfd5bfd7dfd76fd29fd8afcd3fb65fb7cfb41fc97fd17ff780091015102e702;
    inBuf[6904] = 256'h7303d9030a04e7035e03b3023002f6013202ca0279033d041205eb05f6062608;
    inBuf[6905] = 256'h3e093f0a110b990b0d0c6a0c8d0c910c680c0a0cca0bc40bea0b600cfb0c890d;
    inBuf[6906] = 256'h430e370f65100d12fb13d5159117ea18b2192a1a491a031aa5192a199d186b18;
    inBuf[6907] = 256'h99181a191e1a561b751c971d801e111f951fe81ffe1f222032201a201a20fa1f;
    inBuf[6908] = 256'h9e1f591f161fee1e481ffb1fe5202b227923b62423267e2795286b298229a828;
    inBuf[6909] = 256'h31272d25fd224421fb1f281ff81e111f601f1a20f320ce21c5227623cd230024;
    inBuf[6910] = 256'hcf2338236b2222216e1fb21de91b591a5d19c2188d18e8189819a31a1e1c8a1d;
    inBuf[6911] = 256'h921e021f651ed61ccd1a79183f166f14cc1254112610240f8b0e930ef70e920f;
    inBuf[6912] = 256'h33106a103310b30fd50ec90db80c870b650a8c09f108b108ca08e108db08a708;
    inBuf[6913] = 256'h1e086707a806cf0502056304ee03d40321049204f60408057a046003ef015000;
    inBuf[6914] = 256'hd3fe9cfd9ffcf6fbabfbb7fb2afce5fca3fd40fe9bfea9fe9bfe8cfe76fe59fe;
    inBuf[6915] = 256'h0bfe6ffd9ffcb4fbdafa48fa05fa0cfa61fae7fa84fb2bfca6fcd0fca2fc0ffc;
    inBuf[6916] = 256'h3bfb5afa82f9c6f82df89af70cf795f635f602f60df63bf689f6f8f675f70ef8;
    inBuf[6917] = 256'hc4f86ef9f6f942fa26fab5f913f94ef898f708f781f607f691f5fff46bf4e9f3;
    inBuf[6918] = 256'h72f32df32bf356f3bef358f4eff478f5d4f5ccf56df5c5f4d4f3dbf206f25af1;
    inBuf[6919] = 256'h03f10af14af1ccf176f204f369f386f32cf380f2aaf1bcf004f0a6ef8eefd4ef;
    inBuf[6920] = 256'h6bf024f107f2f3f29af3edf3ccf313f302f2caf07aef50ee58ed7decf4ebe0eb;
    inBuf[6921] = 256'h3dec2fed8aeee4ef17f1f4f15cf291f2b4f2b1f29df264f2e7f166f10af1d5f0;
    inBuf[6922] = 256'he8f020f12cf113f1d7f078f03ff043f062f0b2f025f19af13bf201f3bbf36df4;
    inBuf[6923] = 256'hf6f429f52ef513f5ccf482f437f4daf3a7f3c1f32cf40bf53bf665f769f817f9;
    inBuf[6924] = 256'h4bf935f9eef87af808f8a2f742f721f757f7dff7cdf8faf91cfb18fcc3fcfefc;
    inBuf[6925] = 256'heafc9cfc18fc8cfb06fb81fa29fa15fa50fa02fb26fc8dfd0bff52000d012501;
    inBuf[6926] = 256'h9f0096ff5afe2cfd28fc74fb1dfb1efb91fb7bfcc0fd3effb100c60153024902;
    inBuf[6927] = 256'haf01b60091ff60fe4ffd7ffcfafbcefbf7fb52fcc6fc42fdb6fd2afea6fe13ff;
    inBuf[6928] = 256'h57ff56fff4fe44fe78fdc0fc48fc21fc33fc62fca2fce6fc35fd91fdd8fddcfd;
    inBuf[6929] = 256'h7efdaefc97fb94faf6f9f4f996fa9dfbb2fc96fd1cfe44fe2ffeeffd8cfd0afd;
    inBuf[6930] = 256'h5efc8ffbbafaf9f964f916f911f953f9def9a0fa7ffb5ffc1ffdaafd05fe38fe;
    inBuf[6931] = 256'h47fe2afecbfd14fd15fc01fb24fac5f906facffae0fbf5fcddfd8cfe14ff81ff;
    inBuf[6932] = 256'hceffeaffb9ff2bff57fe5dfd62fc93fb04fbbbfacdfa39fbf4fbfbfc2ffe69ff;
    inBuf[6933] = 256'h9900a4016602d902e3026e02a001a600b9ff31ff30ffa0ff6f005e012d02e202;
    inBuf[6934] = 256'h7703dd032e0452042804d2036203ef02c202e2022b03a3031d047404d7044e05;
    inBuf[6935] = 256'hd705a20699079408a609b00a890b4f0ce70c2f0d560d4a0df80c950c150c720b;
    inBuf[6936] = 256'h010bd60a000bc20bf00c440ebd0f1911351252135c143515ee153b16e9153b15;
    inBuf[6937] = 256'h4d145b13ec1208139513a014ce15dc16eb17d7189b197b1a501bfd1ba71c131d;
    inBuf[6938] = 256'h2c1d331d141dda1ccf1cca1cad1c981c501cd21b771b421b561bf71bdf1cce1d;
    inBuf[6939] = 256'hb61e351f331fee1e5b1e981deb1c301c6b1bd81a611a251a651aed1a9e1b6e1c;
    inBuf[6940] = 256'hfc1c2c1d241dce1c4c1cd61b3a1b641a5e19ee172e167114c8127611b9106210;
    inBuf[6941] = 256'h6010a510e3100f113a1136110d11cb104110780f870e5a0d130cda0aa3098c08;
    inBuf[6942] = 256'hb607080798066d065b065e0667064106e5054a0553041b03c4015d001eff21fe;
    inBuf[6943] = 256'h53fdb7fc37fcadfb2bfbbcfa5cfa22fafef9caf981f916f986f8faf77cf70bf7;
    inBuf[6944] = 256'hb0f64ef6d4f555f5d6f46bf433f41ef413f409f4dcf38cf337f3e1f298f263f2;
    inBuf[6945] = 256'h18f2a2f103f130f04fef96ee0feed2ede6ed19ee59ee93ee9bee7aee48ee05ee;
    inBuf[6946] = 256'hdeedf3ed2fee96ee1cef8cefecef3ff065f06af049f0d4ef23ef50ee60ed94ec;
    inBuf[6947] = 256'h11ecbeebb2ebe6eb36ecbeec80ed4aee16efbbeff4efd3ef6befbfee18ee95ed;
    inBuf[6948] = 256'h22ede8ece9ec06ed60edeeed79ee09ef86efc3efe8ef03f0fceffeef08f0f7ef;
    inBuf[6949] = 256'hf5ef09f010f028f036f0fdef96ef05ef47eeaeed5ced3eed7ced04eea3ee73ef;
    inBuf[6950] = 256'h5bf01df1bef11df20ef2ccf17af121f104f11af12bf148f15ef156f165f18cf1;
    inBuf[6951] = 256'ha0f1b4f1aef16df12bf100f1eaf024f1a7f14af224f317f4f0f4bef567f6bdf6;
    inBuf[6952] = 256'he0f6bff631f656f525f4a0f22bf112f090efffef53f13ff395f5fbf71bfaf8fb;
    inBuf[6953] = 256'h72fd55fea3fe32feddfce3fa81f807f605f4cdf27ef239f3cbf4d7f628f96afb;
    inBuf[6954] = 256'h50fdd5fedaff3d00150057ff08fe76fce3fa8bf9c7f8a5f8fef8bef9aafa93fb;
    inBuf[6955] = 256'h8afc8ffd94fea1ff8d001c014401f200240010ffd7fd92fc7dfbb4fa44fa52fa;
    inBuf[6956] = 256'hd6fab1fbd1fc09fe28ff1f00d30023011701ad00ebff02ff13fe26fd4ffc80fb;
    inBuf[6957] = 256'ha8fae4f95af933f99ff999faebfb5dfdaffeb3ff6d00dc00f0009f00ceff73fe;
    inBuf[6958] = 256'hb9fce3fa3cf90ef879f770f7e0f7a6f89af9abfabefbb1fc76fdfdfd3afe35fe;
    inBuf[6959] = 256'he8fd4cfd6cfc5afb3bfa48f9aaf86af87cf8b9f8faf839f97ff9e1f973fa2afb;
    inBuf[6960] = 256'he9fb92fc0cfd4cfd5cfd3efdeefc68fca8fbbdfacef904f985f86cf8b1f845f9;
    inBuf[6961] = 256'h12faf7fadffbb5fc5ffdd2fd10fe1ffe12fefbfdd6fda1fd54fde9fc71fc09fc;
    inBuf[6962] = 256'hbffbaafbc9fb08fc69fceefc99fd7cfe8dffa4009b0142026f022b028b01ab00;
    inBuf[6963] = 256'hbcffdbfe14fe8afd51fd76fd1afe34ff990027029b03b9047905d905dd05b005;
    inBuf[6964] = 256'h5805ce0429046a039e02f80191017201bb0163025703a1041c069307e508d509;
    inBuf[6965] = 256'h380a320ae20975092d090209cf088d081f088b071707de06ea064e07df078208;
    inBuf[6966] = 256'h5609580a8c0bfd0c670e7f0f2e104f10f00f5b0fa70ee00d2c0d760cc70b600b;
    inBuf[6967] = 256'h4c0b9b0b640c6d0d860ea90fa7106d111112691267122d12b5112511bd107310;
    inBuf[6968] = 256'h3f102a100810e20ff10f3510bd108f115f12fb125f1365132313cc125012ba11;
    inBuf[6969] = 256'h26117b10d30f5d0f0b0fee0e1d0f710feb0f97104111d31144125d122712ca11;
    inBuf[6970] = 256'h4011ac102010740fa90ed80dfd0c4b0cf00bd00bea0b310c720cb80c160d6c0d;
    inBuf[6971] = 256'hbd0dfa0dee0d9f0d250d7f0cd40b310b6f0a91099e089207ab061706d305eb05;
    inBuf[6972] = 256'h4d06c3064e07e7077008ef0852096c094609e8084d089907cf06d405b6047b03;
    inBuf[6973] = 256'h2f0214015200eaffebff3900aa0048010c02e102cb039e0420054305f7043c04;
    inBuf[6974] = 256'h43032002db0097ff5efe40fd72fc08fcfefb5bfcfbfcb3fd80fe49fff7ff8c00;
    inBuf[6975] = 256'he100cf00590077ff40fefafccffbe5fa6afa51fa81faebfa5ffbbbfbfdfb15fc;
    inBuf[6976] = 256'h05fcebfbc2fb8efb62fb30fbf7facafa9efa72fa55fa31fa02fad6f9a6f97bf9;
    inBuf[6977] = 256'h70f97cf99ff9dff921fa56fa80fa84fa5cfa12fa9bf907f974f8e9f77cf748f7;
    inBuf[6978] = 256'h49f782f7fcf79ef855f90efa98fad9facffa73fae4f952f9d2f87cf860f868f8;
    inBuf[6979] = 256'h8ef8d1f81ff977f9dbf934fa75fa9afa8bfa4bfae9f96ef9f8f8adf899f8c8f8;
    inBuf[6980] = 256'h39f9c9f95efae5fa48fb89fbb9fbdafbf6fb16fc29fc2bfc1dfcf7fbc2fb94fb;
    inBuf[6981] = 256'h75fb76fba6fbf5fb56fcbbfc0cfd48fd7efdb1fdeafd2ffe67fe80fe70fe2dfe;
    inBuf[6982] = 256'hc9fd63fd0ffddefcdafcf0fc17fd54fdabfd2ffef9fef9ff11011102bb02e902;
    inBuf[6983] = 256'h9d02e801f400f6ff09ff42febcfd7efd99fd19feeffefdff20012502e8025d03;
    inBuf[6984] = 256'h7b034a03df0245028b01ca00040047ffa8fe34fe06fe41feebfefaff4a019702;
    inBuf[6985] = 256'ha5035504980483043804be03170343023b011a0017ff5dfe13fe46fed9feabff;
    inBuf[6986] = 256'h9f0094017a024203ca03fb03cd03400374029101ab00d5ff16ff68fedffd97fd;
    inBuf[6987] = 256'h9ffd02feb1fe80ff4f00070196010402520270025a020e028c01ea00380073ff;
    inBuf[6988] = 256'ha3fec9fdeffc41fce5fbeffb61fc15fdd3fd7bfef5fe3fff68ff6fff42ffdefe;
    inBuf[6989] = 256'h3bfe62fd7ffcb4fb19fbcafabffae9fa45fbb7fb2afc98fcebfc22fd51fd75fd;
    inBuf[6990] = 256'h8dfd96fd6cfdf6fc3bfc3ffb26fa2af966f8f9f7faf75ff81ef92efa5cfb7cfc;
    inBuf[6991] = 256'h66fde2fddcfd65fd8bfc7dfb71fa7bf9baf84af826f859f8eef8c4f9ccfaeefb;
    inBuf[6992] = 256'hfbfce3fda1fe1eff5dff62ff14ff7efeb6fdc4fcd7fb17fb8dfa52fa75fae3fa;
    inBuf[6993] = 256'ha1fba5fcbdfdd0fec1ff6900d800230146014f013201ca00250064ffaafe3bfe;
    inBuf[6994] = 256'h3afe91fe30fffdffd500d2010003450482057306c206600668050f04b902ab01;
    inBuf[6995] = 256'hf2009a009300bb002101c9019e029c039f04720509065e066c0659063106f005;
    inBuf[6996] = 256'ha6054d05dc046d041104d003ca0305046d04fc049205010641064a061d06e605;
    inBuf[6997] = 256'hbd05ab05be05e305f405e705a9052d058b04ca03f4022b0286011b0117018a01;
    inBuf[6998] = 256'h6f02ba0337059e06b80750084908be07d806ca05d5040f047303f70282020b02;
    inBuf[6999] = 256'hb0018901a8011202a0021e0374039a03a303bd03f80344048504890435049d03;
    inBuf[7000] = 256'he2022f02ac016201470153017e01c20123029502040363039f03b303a6037d03;
    inBuf[7001] = 256'h3f03fc02c402a902b902eb02210337030b039602f0014401b60059002300fbff;
    inBuf[7002] = 256'hd3ffb1ffabffddff4e00e9008501f70122020b02cc01860153013c0139013a01;
    inBuf[7003] = 256'h2f010d01d30085002b00cfff7bff38ff0eff06ff21ff5effb6ff160062008100;
    inBuf[7004] = 256'h5700daff14ff1ffe24fd51fcc8fb98fbc6fb42fcf4fcc7fda2fe6cff11007a00;
    inBuf[7005] = 256'h96006300edff4dffabfe27fed3fdb6fdbffdd3fde0fdd6fdaefd71fd25fdd3fc;
    inBuf[7006] = 256'h8dfc5dfc4ffc71fcbdfc23fd91fde4fd06fef5fdb9fd69fd26fdfefcf1fcfbfc;
    inBuf[7007] = 256'h0dfd21fd43fd7dfdd4fd49fec1fe1eff50ff4aff14ffc3fe5ffeecfd72fdf3fc;
    inBuf[7008] = 256'h7dfc2ffc18fc3cfc95fc00fd5ffda4fdbffdb4fd8efd51fd0cfdd7fcc7fceefc;
    inBuf[7009] = 256'h53fddcfd5efeaffeaafe49fea7fde4fc26fc92fb35fb20fb5ffbf3fbcffcd8fd;
    inBuf[7010] = 256'hd6fe8effd9ffa2fffcfe19fe26fd49fc94fb01fb86fa23fadff9cdf9f9f95efa;
    inBuf[7011] = 256'he7fa76fbeafb2efc40fc26fcebfba2fb5efb36fb43fb94fb24fcdbfc88fdf5fd;
    inBuf[7012] = 256'hfafd88fdaffc9afb7efa8ef9edf8a9f8b6f8fff86cf9e4f960fadcfa4efba8fb;
    inBuf[7013] = 256'hd4fbb8fb50fbb2fa02fa71f926f926f966f9cff945fabcfa32fb9bfbf0fb2bfc;
    inBuf[7014] = 256'h3cfc25fcf2fba7fb50fbfbfaaefa7ffa86fabefa1afb75fb9afb77fb21fbc0fa;
    inBuf[7015] = 256'h94fac1fa2ffbaffb07fc08fcc0fb64fb1efb19fb5afbb6fb12fc63fc9ffcdffc;
    inBuf[7016] = 256'h30fd7afdadfdb4fd7bfd1ffdd0fca6fcbffc16fd7ffde8fd46fe8efedafe32ff;
    inBuf[7017] = 256'h78ff97ff70ffe3fe09fe0ffd1afc67fb18fb2bfbacfb8dfca2fdc7fec6ff5700;
    inBuf[7018] = 256'h6f001f008cff0dffdcfe01ff7cff2900d0006301cb01e2019d01e600b0ff36fe;
    inBuf[7019] = 256'hc7fcacfb38fb7ffb51fc86fddffe28005b016a022b038c0365039b025401c7ff;
    inBuf[7020] = 256'h30fee5fc0cfca4fbb0fb12fca3fc5dfd2bfefafed6ffbc009c0177022e039703;
    inBuf[7021] = 256'ha4034a039302b401d000f5ff2cff5efe6ffd77fc9bfb10fb19fbc4fbf0fc69fe;
    inBuf[7022] = 256'he0ff180101029902e402f502c50248029001af00c2fff9fe6afe17fe04fe1dfe;
    inBuf[7023] = 256'h50fe9efe00ff75ff0a00c10090016d022f03a803ba035b03a502d30117018d00;
    inBuf[7024] = 256'h3200e7ff90ff33fff1fefafe71ff46003f0115029002a3027602430239026902;
    inBuf[7025] = 256'hbd0212034703550346032d0317030803f702dd02b4027f0245021102ed01e801;
    inBuf[7026] = 256'h13027102ff02a4033a049904a6045704bc03fa022f027b01f4009e008100a700;
    inBuf[7027] = 256'h0e01b701950283035804f0042805020599040c0486032803f102df02e802fb02;
    inBuf[7028] = 256'h1b0351039003d003fa03e8038e03f3022b025f01b800440009000a0034008f00;
    inBuf[7029] = 256'h2501ec01db02d803ac043205550503055404720377029001e40078005a008e00;
    inBuf[7030] = 256'hf9008f0148020a03d1039b044505b805de059005d104bf0372021f01f3fff2fe;
    inBuf[7031] = 256'h29fea5fd66fd8efd4bfea0ff8701d2031a060b086809fc09ce09f90883078705;
    inBuf[7032] = 256'h2e03a10041fe86fcbbfb12fc77fd80ffbf01dd039305de06d6077108ac087d08;
    inBuf[7033] = 256'hc6079b063305b70368027301d20084008500b30003017201e1015502e2028803;
    inBuf[7034] = 256'h560453054b061a07a407c70799074707dc066706e5052a0530041f0321028401;
    inBuf[7035] = 256'h8601160204030b04ce0433055c0564057a05ad05bf057a05c704a40360026b01;
    inBuf[7036] = 256'hff003701f801ea02d1039c043f05d2056b06e70628071f07b506020634055204;
    inBuf[7037] = 256'h6d039302b901f5006e002b00370092001601b8017b0246030904a904e5049f04;
    inBuf[7038] = 256'he903e302dc012101c100ad00c500d400d200e0000c016b01f6017502c202d102;
    inBuf[7039] = 256'ha00250020702bf0170010f018900f2ff77ff2dff27ff61ffaaffe4ff0200fbff;
    inBuf[7040] = 256'he4ffdbffdaffe0ffe7ffd4ffa1ff5cff0dffd0fec3fee6fe38ffaaff12005400;
    inBuf[7041] = 256'h60002b00c9ff5fff07ffddfef3fe3bffa4ff19007700a800a4005e00dbff33ff;
    inBuf[7042] = 256'h7afed6fd6ffd59fd9dfd2cfed4fe5cff98ff6cffe7fe44fec0fd9afdf1fdb3fe;
    inBuf[7043] = 256'hacffa3006101d3010b0225023a0250024c02080270018b0084ff9ffe16fe00fe;
    inBuf[7044] = 256'h52fee0fe77fffcff6c00d4004601ba01180240022002c1014a01e900bb00cb00;
    inBuf[7045] = 256'h01013e016c018a01a201ce011a028302fe027a03e6033a046e0477044a04e603;
    inBuf[7046] = 256'h5703c102530230026102cd02400384037e033603d9029d02a7020303a5037004;
    inBuf[7047] = 256'h4a051a06c0061607f70649061a05ab03570275013a019d0168025e0351043305;
    inBuf[7048] = 256'h1206f306c10758088d084b08a507c506d705fb043d049403040397025d026002;
    inBuf[7049] = 256'h9802ec0247039703e2033b04b0043905c30525063c0600067d05c9040f046903;
    inBuf[7050] = 256'he0027a023202fe01e301ed01210289022503d9038204ef04f20471046b03f501;
    inBuf[7051] = 256'h4900a4fe40fd5efc29fcaefce4fd9dff800132036104d50488048f0301020100;
    inBuf[7052] = 256'haafd24fbc8f809f74ef6dbf69af811fba8fdd3ff4101f6012202e80158016800;
    inBuf[7053] = 256'h0bff63fdb6fb47fa3ff98ef8f5f742f776f6c2f576f5cdf5c0f61ef89bf9f5fa;
    inBuf[7054] = 256'h20fc20fddcfd36fe03fe1bfda3fb02fa9ef8c4f77ef782f76df707f756f6a1f5;
    inBuf[7055] = 256'h37f53df5aef55ef61ff701f834f9cbfaacfc70fe6eff2aff91fdf6fa0ef89ff5;
    inBuf[7056] = 256'h19f48ef3c1f33ff4b5f403f524f534f563f5d0f5a6f604f8dcf9f4fbe6fd31ff;
    inBuf[7057] = 256'h87ffecfe9ffd18fcc7fac8f904f950f875f776f68df5f1f4cbf426f5dcf5c9f6;
    inBuf[7058] = 256'hd7f7eff812fa35fb2dfcd6fc1efdfdfc98fc32fceafbd1fbddfbcefb6ffbaefa;
    inBuf[7059] = 256'h90f94ef83ef79bf68ef620f725f872f9e6fa4ffc8afd76fedcfea7feebfdd9fc;
    inBuf[7060] = 256'hd3fb38fb25fb7cfbf0fb12fca9fbd3fad8f92bf931f9fdf95ffb01fd6cfe4dff;
    inBuf[7061] = 256'h82ff03fffffdbdfc75fb65fac4f99af9e8f99afa77fb50fc0afd86fdd0fd0efe;
    inBuf[7062] = 256'h56fec4fe67ff2600df006d018f011401e9ff18fef1fbfdf9c2f8a9f8c1f99dfb;
    inBuf[7063] = 256'h9efd26ffc8ff90ffdffe12fe74fd1bfdd5fc81fc31fc13fc67fc55fdb5fe2800;
    inBuf[7064] = 256'h4001a9016201b200f2ff7eff7cffccff4000aa00dc00cd007400b2ff75fec1fc;
    inBuf[7065] = 256'haefa98f8f5f619f637f648f7fef8fcfaf9fcb8fe22002d01d00118021602da01;
    inBuf[7066] = 256'h87012f01c300360079ff76fe3bfdeafb95fa54f942f874f70ff73bf709f862f9;
    inBuf[7067] = 256'hf3fa42fcedfcc6fcf2fbf4fa60fa91fa97fb1dfd85fe51ff44ff6ffe35fd04fc;
    inBuf[7068] = 256'h21fb9efa5efa30fa03fadef9d5f9fbf93bfa62fa42fabbf9dbf8e8f72cf7e6f6;
    inBuf[7069] = 256'h46f745f8acf940fbb4fcbffd46fe57fe21fee8fdcbfdc1fd97fd09fdfafb9efa;
    inBuf[7070] = 256'h50f973f847f8aef850f9d7f90afaf2f9cdf9cef905fa64fac2fa0efb62fbe9fb;
    inBuf[7071] = 256'hc2fcedfd2aff1f007d00180011ffc4fd9cfc06fc47fc47fdb9fe35003e018901;
    inBuf[7072] = 256'h1b012300f0fed1fde1fc14fc52fb87facaf956f96af938fab9fb9dfd7dfff200;
    inBuf[7073] = 256'hb501cc0190016d01cd01dd026f0426068b0741084008bd07e506e005b4042f03;
    inBuf[7074] = 256'h3701ecfe8ffc81fa1af980f8b3f8a0f92cfb4efde3ff9d0229052e076d08f908;
    inBuf[7075] = 256'h1a0915092009430958094109e60837083807e4052c043a02660014ffb3fe6fff;
    inBuf[7076] = 256'hfa00cc0252041d052505bb0443040d042d048804fe047505e1054e06ac06d006;
    inBuf[7077] = 256'ha1061c065d05a604350428047f040905940512067806be06fb0635074f074007;
    inBuf[7078] = 256'h01077b06ad05a804830368028a0112011901930169027d039f049d054f067d06;
    inBuf[7079] = 256'h0006e704770323027f01e101410341052a074908470832076a058303ea01c400;
    inBuf[7080] = 256'h1100baffa7ffe6ff840076019502aa038f0436059c05c1059a050005e1036302;
    inBuf[7081] = 256'hcb006fff9bfe54fe70fec8fe43fff2ffff006302d603f1044805ad046703fe01;
    inBuf[7082] = 256'hf6009400bb001001420132010a010e015001a801ca017901ca002500faff7f00;
    inBuf[7083] = 256'h8b01a00249036f034d035703d9039d041505bd045b0339010eff84fde8fc18fd;
    inBuf[7084] = 256'ha2fd28fe94fe0dffcaffe000260259034804ec046f05fc059006120763076707;
    inBuf[7085] = 256'h2507ac06e205a004d6029a005afed2fc91fcbafdf7ff78025504fb045c04d802;
    inBuf[7086] = 256'h1201afff20ff84ffae005002f4031205650501052a045b031303710342043705;
    inBuf[7087] = 256'hfe058006e8066a071708cb082809d808b807d2056903e20086fe92fc39fb92fa;
    inBuf[7088] = 256'ha0fa50fb6cfcc2fd3bffcc008a028804a0068b08ef097b0a320a6e099f082a08;
    inBuf[7089] = 256'h380881089608230800076205bf0362026401bd003400a3ff24ffddfee6fe4cff;
    inBuf[7090] = 256'hfaffd200c901eb024704c70526072f08ba08a70816083b071006980408039e01;
    inBuf[7091] = 256'hce002101b2022505d607f709070b220bc30a7b0a9b0aea0add0af90909085a05;
    inBuf[7092] = 256'h95024900c7fe0ffed3fdd4fd0efe90fe82ff040100035005c707230a330cd00d;
    inBuf[7093] = 256'hbb0ee80e880ed10d140d950c390cbf0beb0a810987075605410386015400a0ff;
    inBuf[7094] = 256'h4dff5cffd1ffc0003c022f046a06aa08900adc0b6b0c220c1e0ba009da071906;
    inBuf[7095] = 256'hac04a7031e032703a9039004de055a07b508ae09ff099709b608bc070c07e006;
    inBuf[7096] = 256'h0f073e0711074b060605a10367027f01e6006000c3ff2affd5fe1eff39000002;
    inBuf[7097] = 256'h19040a064b07a407380749065305e7044e05950681086b0a8f0b6a0bd6092c07;
    inBuf[7098] = 256'h3404b2011c0073ff3ffff9fe58fe5afd4bfc98fb74fbdefbc8fc1cfed9ff0902;
    inBuf[7099] = 256'h8d0420076309fe0ae00b340c210cb60bc60ae208c5059c01f8fcc6f8fdf51af5;
    inBuf[7100] = 256'h0ef657f825fbc1fdd4ff56018302be03440516070309a30a710b010b31093c06;
    inBuf[7101] = 256'haf023cff95fc16fbaafafafa97fb1efc76fcc5fc2ffdc3fd7afe29ffa9ff0400;
    inBuf[7102] = 256'h700020011c023003f103e403c302bd0071fea0fcf3fbb8fcb0fe37019c035705;
    inBuf[7103] = 256'h220614066d055704e1020b01cefe2cfc5df9baf698f439f3b7f2edf288f343f4;
    inBuf[7104] = 256'h06f506f6c1f7bbfa20ff8b04090a540e5510a80fbe0c9e0885046d0192ff8afe;
    inBuf[7105] = 256'ha4fd2dfcc3f995f632f33cf045eea7ed5dee29f0aff28df56ff81ffb94fddfff;
    inBuf[7106] = 256'hfa01c3030c058805f8047b038401a3ff6afe21fe90fe2bff53ff91fed1fc5bfa;
    inBuf[7107] = 256'hbcf78cf53af4f9f3cdf458f603f850f9dff997f9e2f859f866f82df954fa2bfb;
    inBuf[7108] = 256'h39fb73fa47f997f834f95cfbb1fe4402d4046a05a803dafffcfa4af6d7f240f1;
    inBuf[7109] = 256'h67f195f2f6f3d7f4f4f4b4f4b1f458f5daf6faf820fbe6fc1dfec6fe1dff41ff;
    inBuf[7110] = 256'h1effa0fe9afdd4fb5cf952f6d3f24fef59ec6eea06ea43ebb5edb7f09af3d3f5;
    inBuf[7111] = 256'h60f79ff801faeafb56fed600ed020f04c3030d022aff67fb53f772f31bf0b3ed;
    inBuf[7112] = 256'h71ec41ec04ed51ee70efeaef79ef28eeb5ec14ecedecb0ef30f484f9adfeba02;
    inBuf[7113] = 256'hcf048d04ff0184fd11f8eaf242ef04ee44ef1ff248f560f795f733f62af482f2;
    inBuf[7114] = 256'h21f216f397f4daf529f615f5f8f274f0feed22ec35eb2eeb22ec14eec5f00df4;
    inBuf[7115] = 256'ha8f713fbeefde1ff8a00defff5fdfffa9af75ef4a5f1cbefcdee35eeb7ed12ed;
    inBuf[7116] = 256'h26ec5ceb33ebf5ebeaede5f042f477f7edf918fb05fbe6f9e9f7a2f58cf3c9f1;
    inBuf[7117] = 256'ha2f02ff033f0a5f079f165f238f3a9f339f3aaf119ef12ecade9e0e82cea94ed;
    inBuf[7118] = 256'h2ff2a0f608fae6fb24fc6bfb51fa06f9d6f7def6fcf542f59cf4a2f312f2beef;
    inBuf[7119] = 256'h9aec26e903e6b3e3c9e298e324e66dea11f03bf600fc450021028301f4fe6afb;
    inBuf[7120] = 256'h3df855f6e6f5bff611f8cef860f89cf6c8f3ccf08cee76ed92ed2cee39ee37ed;
    inBuf[7121] = 256'h3beb12e940e8f5e959eea9f432fbfafff001470145ffbffd01fe28001803d604;
    inBuf[7122] = 256'hb6035fffb3f88ef12eecd9e974ea0ded22f059f25af386f389f31df48af58ef7;
    inBuf[7123] = 256'hbdf99bfbdbfc9afd27feeefe6900c002ac0589084b0a020a6507ca0228fdcaf7;
    inBuf[7124] = 256'h83f37cf06beeccec6aebb6ea48eb6fed0bf161f57bf9d9fc96ff470288056e09;
    inBuf[7125] = 256'h700db61070125812ca10540e6b0b2908440479ffeaf92df43cef05ecefeacdeb;
    inBuf[7126] = 256'hffeda7f035f3a0f521f803fb6cfe2202b505bc08fe0a820c680dbf0d760d7b0c;
    inBuf[7127] = 256'hdb0af008400747063506a506c106ab05b802ddfdf6f754f24ceee9ec72ee42f2;
    inBuf[7128] = 256'h38f72bfc47006303dd054108ed0ac40d391095114611360fd10bc107c3037400;
    inBuf[7129] = 256'h10fe9ffc1cfc72fca1fdabff3d02da0400070a08a80736065404ba0219029a02;
    inBuf[7130] = 256'hd4033b055606f4063e077b07d7072708ef07e6061505b20243005efe2dfda4fc;
    inBuf[7131] = 256'hc8fc93fd2affbb011a05e908b50ced0f53120c141115411584149412600f560b;
    inBuf[7132] = 256'h0607f60291ffeafc02fbfdf902fa4cfbe4fd4c01dd04fc07140a0a0b340bdd0a;
    inBuf[7133] = 256'h5e0a260a620a2c0b840c030e380fd10f850f8b0e790d8c0ccb0b160bed090b08;
    inBuf[7134] = 256'hd705eb03e8024103bf04b50663082e090d096808a007220730078507d6072108;
    inBuf[7135] = 256'h6008d408f209d90b630e1d112613e4135413b111b00f1e0e110d280cf90a0909;
    inBuf[7136] = 256'h740606047f024f027e036d05780767093d0b440dac0ff51167136f139f11520e;
    inBuf[7137] = 256'h9c0a7607b405cc0558079509ca0b200d420d870c6d0bb50a230bd20c690f5212;
    inBuf[7138] = 256'h94147615c0146d12ec0e070b5e07a8048403f403bc058608810b140e3b10f711;
    inBuf[7139] = 256'h7f133315ef164518c318df1780151912270e560a440703059103fc021503d703;
    inBuf[7140] = 256'h5a0549075d098f0bb50dfa0fd5123d16d519191d131f0e1f041d3b195d14440f;
    inBuf[7141] = 256'h5e0afd057d02160049ff9d00e903a608f60d76122815ec15f114ea12d710390f;
    inBuf[7142] = 256'h480e2c0ebe0ef00fd4112d14a916d618ed19721950176f133f0e9b081f0382fe;
    inBuf[7143] = 256'ha0fbd5fa3bfcb8ff8b04d209e40e231376163d19951b5f1d351e491d241a0715;
    inBuf[7144] = 256'hb30e8908f3039801a501d1032e07f90aa70e5b117512cf11540f7a0b4e07be03;
    inBuf[7145] = 256'h9a018901a703c007430dfb1283179b198018c41425108b0c760b270d21104812;
    inBuf[7146] = 256'h0312bb0e78094504d1000000b901dd043808fe0a910cb90c8f0b32093a06ba03;
    inBuf[7147] = 256'hb602e1032607580bf40ebf1032100e0ece0b830a8d0a770b0b0c660b9a097107;
    inBuf[7148] = 256'h2e06c6060d09fa0b250e530e4d0ce2084505b102d8017d02f3037e057706ae06;
    inBuf[7149] = 256'h51069f0511051405c1051b07eb088e0a6d0b470b140a32082d064b048e02de00;
    inBuf[7150] = 256'h3fff26fe4afe3300f403b908ec0c2d0fce0ef10ba3074f03ebffdefd2cfd98fd;
    inBuf[7151] = 256'hf3fe2301e703af06a9081409c207240530022700e4ff6701ff037f06af07e906;
    inBuf[7152] = 256'h5004b80072fdbcfb28fc8efe2602c6057308c909fb098409dc082b082c076205;
    inBuf[7153] = 256'hb5028dff90fc88fa00faa6fa84fbc4fb03fb78f913f8ecf76ef92bfc31ff8401;
    inBuf[7154] = 256'h9b02be02dc02ae0346053007a208cf08950776050d03c300abfe7ffc0ffa91f7;
    inBuf[7155] = 256'h96f5dff401f607f971fd5702b106b9090b0ba50aed08690684037d0046fdaaf9;
    inBuf[7156] = 256'hc1f5ebf1b3eedaecdbec7dee10f1b1f39bf592f6ddf6fef68bf7cef8b7fa30fd;
    inBuf[7157] = 256'hfdffbb022405d00632072d062504b501aeffb2fea7feccfe0cfe83fb0ef761f1;
    inBuf[7158] = 256'hd1ebfbe7e2e6a9e8c7ecf4f1a6f6e3f92dfb76fa70f807f6edf3c4f2cdf2b7f3;
    inBuf[7159] = 256'h30f5f5f6b6f881fa90fce6fe5a0176037904ca0314017cfce5f686f189edd0eb;
    inBuf[7160] = 256'h48ecebed7befbcef0dee1deb48e8bde643e789e943ec5dee59ef67efaeef61f1;
    inBuf[7161] = 256'hcaf48df9bdfe21030f06700768076606c6049302e9ffd2fc3cf946f5f2f054ec;
    inBuf[7162] = 256'h11e8d6e411e325e3c2e4d7e68ae83ce9b0e8a7e722e7c2e71aea38ee66f3e8f8;
    inBuf[7163] = 256'hcafdc100fb003dfee0f85df2b8ec9ce901ea80ed6cf2e0f642f9dbf87bf698f3;
    inBuf[7164] = 256'h7af11af161f234f48af583f59cf34df052ec2de887e4a7e17cdf6ddedadebae0;
    inBuf[7165] = 256'h22e4b5e862ed69f167f431f64af744f81ef9b9f9b0f98bf87bf606f4b6f129f0;
    inBuf[7166] = 256'h57efaaeee7ede4ec97eba3ea6deaafea14ebe6ea49e94de67ce287deb7db00db;
    inBuf[7167] = 256'h67dc9fdfcce3a1e780ea6eecdaedddef4ef31cf8a6fd8d023805ec049101a8fb;
    inBuf[7168] = 256'h97f4b3edcde7aae367e16de037e00de042df21de60ddc4dd3fe0eae4c0ea93f0;
    inBuf[7169] = 256'h14f54cf786f7a2f672f5d3f4f6f454f57ef5e0f4e8f2acef72ebb1e688e202e0;
    inBuf[7170] = 256'hb2dfdee1bee5b6e985ec5ced23ec01ea5ae80ce878e902ec75ee19f0a2f04bf0;
    inBuf[7171] = 256'h1df0f1f0f2f2e8f5d4f868fa15faddf75df4f8f0b0eea3ed70ed08ed5aeb6ee8;
    inBuf[7172] = 256'h09e556e2bde1d9e323e88fedb4f260f637f854f83af7e7f506f5cff454f513f6;
    inBuf[7173] = 256'h41f697f51ff442f2daf043f009f069ef73edc0e922e5fde0b2de25df06e23ae6;
    inBuf[7174] = 256'hdcea59efb4f36ff87dfd0e0233051c06b2040b02a9ffa3fe35ff5d006f0018fe;
    inBuf[7175] = 256'hd6f860f186e948e348e05ae109e608edc1f475fbe2ffc601620167ffdefc66fa;
    inBuf[7176] = 256'h1ef807f6ecf39bf148ef64ed53ec58ec65ed38ef7ef1d5f313f64cf888fadbfc;
    inBuf[7177] = 256'h5fffef01510449066607550725060f048001fcfeadfc68fae3f7f2f4f1f1d3ef;
    inBuf[7178] = 256'h9deffcf1c8f6d5fc7c024d067c073a067f036a00dbfd39fc6cfb27fb21fb32fb;
    inBuf[7179] = 256'h79fb3afca9fdd2ff6202ad040206d305f803e8005dfdfaf941f77af5c1f454f5;
    inBuf[7180] = 256'h77f71ffbd0ff94045308580aa40af0094e096609300a280b8c0bdb0a35091f07;
    inBuf[7181] = 256'h2705b403be0207026a01e2009400ca009a01e5025e047b05ce054d0531040f03;
    inBuf[7182] = 256'hc002b903e0059508c10a730b840a81088206b7059506b808340bed0c390d3d0c;
    inBuf[7183] = 256'h800a9808d9061105e002230017fd98fad2f97afbbbff1f06630d12141a19c41b;
    inBuf[7184] = 256'hf91b4d1a73172f143911cf0eeb0c690bd409e407c505b9033a02da019902f003;
    inBuf[7185] = 256'h3405b1053a057b0478041b06ac094e0e7a12ad14f913c810a90c4e092908cb09;
    inBuf[7186] = 256'h550d4e116e14ba1520158813e111ec101111d61165121a127910990d4a0a5307;
    inBuf[7187] = 256'h49057b049304f3043405380571059a061c09210d5d12bf174b1c5c1f3d20b51e;
    inBuf[7188] = 256'h2c1b1f167e10be0bee089208870aa90d9a108c124d137c130f14281535165516;
    inBuf[7189] = 256'h8c14d410660cad08d606630796094d0cdf0e1411491314166b19d41c951fbf20;
    inBuf[7190] = 256'hfe1fa91d131ae315f311ad0e740ca00bce0b630ce40cb60ce40b470b920b460d;
    inBuf[7191] = 256'h86107b1406187c1a831b541ba91af51974192819aa18ce17a516161566132012;
    inBuf[7192] = 256'h7311ad1117131e15ed16de173417db14b411b30eaf0c2e0cdf0c330ecb0f4d11;
    inBuf[7193] = 256'hd312a31477160118fc18db189a17bf157913fd10b70eb60c350be20a2f0c570f;
    inBuf[7194] = 256'h2f14aa19871ebe217722ad20071d1c189d12390d3308110496010e019702f305;
    inBuf[7195] = 256'h240a450ef9110515b917901a3a1d111f811ff01d941a8a16ec128f10ae0f650f;
    inBuf[7196] = 256'h870e480c6808c8031b00d8fe0a01c906b30eba16cc1c1a1f111d8e1738104d09;
    inBuf[7197] = 256'hcb0479032f05f108170d8410e1121a14c0149d15bc16e117cd18e218b3175f15;
    inBuf[7198] = 256'h3b12e90e390c910afa090d0aed090c096007340552035c0224022802f7015601;
    inBuf[7199] = 256'hf5001f02b205d00b8813ec1a66204f23b82374224020de1ca8174e102907d9fd;
    inBuf[7200] = 256'hcef6cff345f51bfa0c00ec04c007e008ab09890bf30e5d137417a519fb185615;
    inBuf[7201] = 256'h3f0f0508330120fc0bfa7ffbd4ffaf054e0bd80e8e0f170ebd0bed0990093b0a;
    inBuf[7202] = 256'ha00a9509b406b50228ff8efd8ffe98013c051d08700937093c085207b7065406;
    inBuf[7203] = 256'he80532056c043304fb04e5068909ea0b050d4b0ccc0959063a037a018a01fb02;
    inBuf[7204] = 256'ha3046205a1047702aeff40fda7fbc5fa2dfa80f9dcf8f3f894fa22fe49030609;
    inBuf[7205] = 256'hff0d0d11ba115910980d370ace067d03080043fc41f855f43bf1c9ef75f043f3;
    inBuf[7206] = 256'hbff7f2fcd101a7053b08cc09f20a4c0c1d0e1d10941191114a0f8d0add034cfc;
    inBuf[7207] = 256'h2ff5b4ef75ec7eeb6deca6ee94f1cbf4f8f7d4fa32fd12ffa3002e02ed03e805;
    inBuf[7208] = 256'hbe07c0086908ac0601045c01cbffe4ff7901b80371058905600315ff6ef98ff3;
    inBuf[7209] = 256'hc0ee2dec57ecf3ee32f3e7f7ecfbbdfe7b00800122025602a501caff08fd2efa;
    inBuf[7210] = 256'h64f887f890faa6fd89002b0248025a01190017ff70fecffdc6fc0ffbb8f824f6;
    inBuf[7211] = 256'hb1f3b2f190f07ff06ff133f34af5eff6b3f78bf7c2f618f649f699f7f6f9f0fc;
    inBuf[7212] = 256'hcdfffd010e03a102b900a6fddbf909f6d4f26ff0bbee70ed52ec97ebcaeb77ed;
    inBuf[7213] = 256'he7f0a4f5a0fae0fea301a6026e02a101830035ff93fd45fb56f80af59bf169ee;
    inBuf[7214] = 256'hb6eb82e9fbe755e79fe7f4e828eba3ede0ef7bf13af28ef249f31af565f8c8fc;
    inBuf[7215] = 256'h0b01c403bd037d00e4fa94f440ef50ec1beccaed2bf002f26cf290f129f0f6ee;
    inBuf[7216] = 256'hb4ee88efc2f08ff123f114ef06ec3ee9fde74ae935ed92f2def7b0fb2ffdb6fc;
    inBuf[7217] = 256'h50fbf2f94cf942f901f9e2f793f539f2b8eef4eb48ead7e945eae9ea80ebf5eb;
    inBuf[7218] = 256'h38ec8decfeec46ed68ed6ced4bed62edeeedbfeebfefb6f041f178f1a7f1f2f1;
    inBuf[7219] = 256'h95f283f357f4eff443f56bf5f5f52df7cff872fa5bfbb4fa68f8daf495f07fec;
    inBuf[7220] = 256'h31e9b4e621e584e4e0e487e683e958ed60f1a9f460f69cf6d8f5a9f4c8f341f3;
    inBuf[7221] = 256'h71f201f1e1ee47ec16eafbe8d8e848e9b7e9aae985e915ead9ebe1ee82f2a9f5;
    inBuf[7222] = 256'hccf702f9f9f9adfb3afea900c001390098fb09f56aee61e918e765e7e6e84eea;
    inBuf[7223] = 256'hc9ea34ea6ce969e98feac2ec2eefc8f041f1eaf07ff01ef146f384f608fab6fc;
    inBuf[7224] = 256'h9cfdc7fccdfa4cf8e1f5acf346f16bee18ebbde749e56fe467e508e875eba0ee;
    inBuf[7225] = 256'h0cf189f24ff341f404f6b9f85ffc54006203ae04a703020050faa7f323edfce7;
    inBuf[7226] = 256'h2ee535e51de84aed91f383f990fdb8fe28fde0f973f698f4f4f4def617f910fa;
    inBuf[7227] = 256'hc3f88bf590f11aee39ec16ec03ed4fee82ef7ef0abf155f360f588f753f95bfa;
    inBuf[7228] = 256'hc1fab8fa4dfaa7f9b9f859f7c3f578f4f3f38ef433f66cf8b1fa80fca6fd5efe;
    inBuf[7229] = 256'hd1fe07ff02ff89fe79fd20fccefabbf916f98bf86af75af55cf2dbeecdeb10ea;
    inBuf[7230] = 256'heee934eb3ded55ef3ff131f391f5a3f818fc3aff61013302ef01620135018e01;
    inBuf[7231] = 256'h240247025c0162ffbffcfaf98af779f588f39ef1e3efcfeefaee9bf074f3e4f6;
    inBuf[7232] = 256'h0cfa57fce3fd0dff4a0004020d049a05e80582046f016afd97f9e9f6c4f5c9f5;
    inBuf[7233] = 256'h17f6c7f56af46ef2e7f0fef079f347f866fe7a045a094e0c3f0d820c4d0aba06;
    inBuf[7234] = 256'hef0130fc31f61af101ee78ed6cef07f302f73dfa14fc7ffc03fc65fb58fb3ffc;
    inBuf[7235] = 256'h0ffe7000df02e2044c063b07ff07ec082e0aaf0b310d4a0e8a0eaf0d7d0bcf07;
    inBuf[7236] = 256'hf2027cfd1ef8b8f3f9f0f3ef5df0ccf1c2f3eef547f8b4fae8fc8efe75ffb8ff;
    inBuf[7237] = 256'hbeff1a001e0195020d0440053c06a607610aac0ed8138b18ff1aed196a15940e;
    inBuf[7238] = 256'h09077e00f6fb76f985f878f897f873f8f4f748f7dff645f7eff8f3fbc2ff8303;
    inBuf[7239] = 256'h7a063508f1088909bc0ad90cb50f9212a114791504158a138911300f770c5109;
    inBuf[7240] = 256'h890508012afc77f7aef3baf126f2f4f4acf93aff7004a708b10be50de60feb11;
    inBuf[7241] = 256'h91132214d4126d0fa20ac40551025201ac026a053408af096509ef073a064505;
    inBuf[7242] = 256'hc30560074a09dd0aa80bcc0b050cd60c4a0e0c105e11b1111811f40fd60e1e0e;
    inBuf[7243] = 256'h5f0dd20bea08860468ff19fbf9f8c9f963fd7b026907d70aef0be90ae3080d07;
    inBuf[7244] = 256'h7f06e807f70ad40e8e1220151516b7157f1420134d121f126512df12e012d311;
    inBuf[7245] = 256'h8c0ffa0b8b0745032300dffeb5fff2018904a306cd0776089c09cd0b040f9d12;
    inBuf[7246] = 256'h55155d16e3159a149b13bb13a9146f150e15c712de0e830ad206a4043504c104;
    inBuf[7247] = 256'h6e05d905d205b2052c067b077509c70bdf0d780fcc102912f3134a168318b119;
    inBuf[7248] = 256'h0019e215d210350b84061d049a043807b20ae00dd30f8b10cd101f11ad113f12;
    inBuf[7249] = 256'h1212ae106a0e140ccd0a770bee0d591183141f16b715a5137410f20cd9094307;
    inBuf[7250] = 256'h3405cf03ee028a02c3027c03bd04d106ce09b70d4d12b916051a6a1b701a8217;
    inBuf[7251] = 256'ha913e60f310d050cdd0b000ce60b230b050a73090f0a170c3e0f591231142814;
    inBuf[7252] = 256'h3c124d0fc60cac0b5e0c670e8b109911cf10e20d6109530499ff2dfcf4fa43fc;
    inBuf[7253] = 256'h28005a06cc0d2915441b201f7320a61f441de919fd158111a40cef07f4037701;
    inBuf[7254] = 256'h070154029504e3064f08a3087e08a908e509840ce20fdc126f1407140112970f;
    inBuf[7255] = 256'h140e4c0e14101f12e51255113c0dbf07af0269ff8efee5ff71026905ae08640c;
    inBuf[7256] = 256'hc710a615dd19fb1b171b2e178a115f0c8c09d909970cc60f4011c90f730bc305;
    inBuf[7257] = 256'hd8002cfe32fe4700fb0218053e069e06c6063507dd077508d5081009ab09340b;
    inBuf[7258] = 256'ha80d881008133d14cf1317129d0ff80c990a7d089106f904d6034a036303e303;
    inBuf[7259] = 256'h8a044e054706a7077209350b530c4f0cfb0acf08b2065105f0046c053706cd06;
    inBuf[7260] = 256'hff06cc065a06ca0514055004be039003f303d3049b05a2058a044a0260ffa4fc;
    inBuf[7261] = 256'hb7faeff957fab6fbe5fdea00a404b708a10cb50f611184116e10970e420c7009;
    inBuf[7262] = 256'h0606fa0198fdc7f995f7a6f709fa14fe6a02ba054907f40646054d030002e301;
    inBuf[7263] = 256'hf802cd04a306b80792071d067f0301001afc49f805f5cff209f2a8f22cf4e3f5;
    inBuf[7264] = 256'h2ff7ddf76bf8d2f9e2fcc001c507ae0d1d124b144f14ba122d100c0d4e09b904;
    inBuf[7265] = 256'h6cff08fa7ef5bef242f2ccf397f6c6f9a9fce6fe8f00e801f5027d0351033602;
    inBuf[7266] = 256'h0c003ffd97fac4f83ef807f96bfa55fbf4fa09f925f67ef358f261f35cf654fa;
    inBuf[7267] = 256'h2efe0b01a70279031604c1046f05b805f304b70206ff37fa07f56ef05bed83ec;
    inBuf[7268] = 256'h0eee95f156f64dfba7ff2f03fc052508cd09ba0a490a1408180494fe44f813f2;
    inBuf[7269] = 256'ha0ec5be890e553e4a7e47fe6a2e9b2ed24f274f658fa80fdb9ff11015e016200;
    inBuf[7270] = 256'h54fe88fb50f864f56bf382f2a4f293f3c5f4d7f594f6d1f6a7f650f613f671f6;
    inBuf[7271] = 256'hc7f717fa2afd4b007a021d0309027eff43fcfbf8c5f57ff2d7ee8bea06e618e2;
    inBuf[7272] = 256'h98df3cdf0ce165e495e8c2ec2ff0c5f287f455f56ff51ff58bf441f4e9f4caf6;
    inBuf[7273] = 256'h11fa77fe0603a00639081107400396fd62f729f2efeef5edf1eedcf074f208f3;
    inBuf[7274] = 256'h27f2b9ef66eccfe836e512e2b4df21ded1dd5adfefe28ae887ef8bf645fcb8ff;
    inBuf[7275] = 256'h8a006fff89fdc3fbd0faa8fa9cfa1efac2f855f637f3d9ef94ecffe961e89ce7;
    inBuf[7276] = 256'h9ce7fde729e821e830e8cbe8c7ea71ee2af30ef8ecfb99fdfefccbfaeaf770f5;
    inBuf[7277] = 256'he3f3f9f23df237f1b5ef48ee94eddbed0fef65f09cf00bef9eebe8e65ae251df;
    inBuf[7278] = 256'h77def3df0ee38be6b0e921ecebedd8ef90f213f628fa17fed700f60174019dff;
    inBuf[7279] = 256'h2ffda2fadbf7b5f4d0f0e3eb7fe6a6e149de64dd48df55e39fe805ee85f2ddf5;
    inBuf[7280] = 256'h0ef825f96df9d7f818f764f416f19aedc6ea1ce979e8aee854e9e2e94deaabea;
    inBuf[7281] = 256'hf2ea37eb56eb10eb9aea3aea41ea4beb81ed86f01df4caf7ecfa64fd21ffcdff;
    inBuf[7282] = 256'h44ff5dfdf3f969f580f023ec68e9c6e8f2e94deccdee75f01bf105f19ef081f0;
    inBuf[7283] = 256'hc2f0f7f0dbf029f0d2ee5fed3cec75eb30eb60ebd9ebd7ec99eefbf0b0f31af6;
    inBuf[7284] = 256'h87f7cef733f752f608f6aaf6e1f728f9b9f9fbf829f7e8f4ecf2eaf113f2f9f2;
    inBuf[7285] = 256'hf7f353f4b3f379f258f124f1a7f2d0f5bff973fdcafffaff34fe25fb7bf7f9f3;
    inBuf[7286] = 256'h11f1beee02ede7eb6deb84ebe4eb46ecb6ec73ed17ef67f283f7b7fdcf034e08;
    inBuf[7287] = 256'h2f0a7f0910070804700165ff41fd59fa51f677f1f0ec06ea75e93feb9fee71f2;
    inBuf[7288] = 256'hcdf53bf8d6f909fb08fcd9fc6dfd8afd25fda4fc6ffcc7fcddfd90ff6301c402;
    inBuf[7289] = 256'h28032c02a9ffcafb32f7c5f245ef52ed3fedd4ee9af121f5eef89afce9ffac02;
    inBuf[7290] = 256'hcc046606ab07b0084709f3083007b603c6fe6af90df5daf263f36af6f5fac0ff;
    inBuf[7291] = 256'ha403d60518069004b70171fecbfb8bfafdfac1fcdffe320007008cfeb4fca2fb;
    inBuf[7292] = 256'h36fcabfe4702de058a08c0096a0905082306250462022801b2002e019702aa04;
    inBuf[7293] = 256'hde066f08d208ef070c06cd030e025401c1012d032c056e07e309700cef0e1411;
    inBuf[7294] = 256'h25126111830ebe09e60351fe1bfae1f7b3f7faf8f8fa42fdbaff8a02f305c809;
    inBuf[7295] = 256'h800d5d108711a9103c0e260b9808b907fd08140c2110e1134e16f416d915a313;
    inBuf[7296] = 256'h2611b60e680c200a8307b2048402bd01dc02d905a509bd0c0a0e310de70aa408;
    inBuf[7297] = 256'h94072308e0097e0bcd0b6f0acb07f5042303f0025f04e8069c09f40bdc0d520f;
    inBuf[7298] = 256'hc410ba122215a517cd19ac1a96199a163912920d210ac0088b09ec0b8f0e3810;
    inBuf[7299] = 256'h5b10f00e980c3e0a5208ee0606065c0500055a05a406f7080e0c140f6311c412;
    inBuf[7300] = 256'h3513331357139c13c31384137112b810150fef0d760d8a0d7a0dd40ce50b3d0b;
    inBuf[7301] = 256'ha30b860d2b1038127a123710f60b6d0768042304cf066c0b9b102a154c18001a;
    inBuf[7302] = 256'h9c1a241ac018b81622147611580fdd0de90c560cab0be10a810aee0a750c2a0f;
    inBuf[7303] = 256'h5a121a15bc16b5160b155212110fce0bf6089306c204b8038f03990410078e0a;
    inBuf[7304] = 256'h970e9e12cd15b2176c182d186917b21635160b163f167f169b168116e415b014;
    inBuf[7305] = 256'h0213c0100b0e2b0b1d081b05a002f5007e00a80159042508740c61103c13c514;
    inBuf[7306] = 256'hfb1457149213221356132c140b15531580142a129a0e9a0adb062204f5020c03;
    inBuf[7307] = 256'h0004930571079409310c100fc211ce13ad14581459135912fc117d125813db13;
    inBuf[7308] = 256'h7313b111c50e510bca07970411024b0076ffd1ff5001bc039f062109b00a310b;
    inBuf[7309] = 256'hd20a440a5e0a790b930d4d10ca125f14dc1447141a13091270116d11e6115612;
    inBuf[7310] = 256'h2c12f3102e0eaa09a703bffc16f615f1e7ee40f007f53bfc8e04b20c76134d18;
    inBuf[7311] = 256'h241bfe1b3b1b7e19471711152c135d11400f8f0c300987054502e0ff88fe23fe;
    inBuf[7312] = 256'h42fe9cfe2dffe7ffb4007201f4015d022903e604f5070b0c21102f13a6149a14;
    inBuf[7313] = 256'heb139a13e11331148313d910180c360696007efc88fa55fa0ffbfefbccfcb2fd;
    inBuf[7314] = 256'h29ff6c0158046c07e8093e0b3f0b1e0a86084507ec06bf076a09fc0a6d0b060a;
    inBuf[7315] = 256'hb00643023ffe21fcd7fc4f005c054a0a850d2c0e740c60092906c10363029a01;
    inBuf[7316] = 256'hcc00abff57fe74fdb7fd59ff0002eb044907a108f408a008110865075d06a804;
    inBuf[7317] = 256'h1302b0fefafaa9f769f5b7f4b0f51bf887fb53ffd902ae0596078308a3083908;
    inBuf[7318] = 256'h8407cd0658063d065d0656069f05cc03db0066fd75faf2f830f9b5fa50fcc4fc;
    inBuf[7319] = 256'h8dfb20f9bef6c8f5e3f6acf9eefc46fffdff69ff92fea0fe3500ff02fc051408;
    inBuf[7320] = 256'h8e0861071a0558028cffe2fc3bfa77f7b6f443f286f0d4ef53f001f2a9f4e9f7;
    inBuf[7321] = 256'h5ffba3fe4601180315044d0406048603d002e501c70045ff52fd19fbcbf8b7f6;
    inBuf[7322] = 256'h52f5eef4a7f559f796f9cdfb67fdf5fd68fde4fbbaf982f7d1f5faf42ef53cf6;
    inBuf[7323] = 256'h72f72df810f81ff7faf586f541f61df876fa52fc20fdf8fc72fc6cfc59fde3fe;
    inBuf[7324] = 256'h4400a50080ff1afd2ffa72f770f54ff4c8f39cf3aaf3c7f3e1f3d7f37bf3ecf2;
    inBuf[7325] = 256'h7df291f2aff3fdf507f931fcb7fed3ff5fffaefd2efb8df85ff6c1f4a4f3def2;
    inBuf[7326] = 256'h20f252f17ef0b4ef23efe7ee0befcfef5bf197f36df65ff990fb86fc21fc81fa;
    inBuf[7327] = 256'h5df86bf6daf4abf3bbf2c8f1f7f0b3f037f18df26cf448f6cff7cef832f934f9;
    inBuf[7328] = 256'hdff819f81df72ff661f5d6f43ef4d6f236f06eec04e83ae441e28be2f5e4c2e8;
    inBuf[7329] = 256'he6ecd9f07ef4dff738fb70feed002702b5015fffa4fb5af758f385f04def61ef;
    inBuf[7330] = 256'h2df0d1f086f04bef9aed22ecb8eb98ec49ee47f0f5f1d8f231f360f379f3a9f3;
    inBuf[7331] = 256'hdcf3b2f327f368f295f123f169f166f212f424f6fef732f977f9b8f86cf70af6;
    inBuf[7332] = 256'hc5f4baf38af29af0e1edb7eac2e709e619e6b9e761ea29ed40efaff0dcf12ef3;
    inBuf[7333] = 256'h2af5b0f7f2f954fb64fbedf987f710f521f332f252f20bf3d8f32ef4a7f359f2;
    inBuf[7334] = 256'h94f0dbeeefed28ee6aef7ef1b5f347f503f6d7f5c6f442f385f178ef52ed43eb;
    inBuf[7335] = 256'h60e91ae8cde788e863ea39eda0f040f48cf7dbf9effaacfa43f976f7eef5ebf4;
    inBuf[7336] = 256'h8af462f4baf355f252f011ee4aec78eb9beb7eecadedd9ee28f0b9f1a1f3eef5;
    inBuf[7337] = 256'h18f876f9e7f969f934f805f73cf697f5e8f4eaf355f271f0baee6eeda7ec3eec;
    inBuf[7338] = 256'he9ebb1ebdbebd5ec10ef6ff26bf665fa97fd86ff50001300e8fe1afdbefaedf7;
    inBuf[7339] = 256'h2ef5eef258f183f00df058ef2deea0ec1deb71ea21eb40ed9ff0a7f4a7f84bfc;
    inBuf[7340] = 256'h4eff7401c5022d038802fd00cffe50fcfef93cf84ef757f722f84ff973faf5fa;
    inBuf[7341] = 256'h69fad7f877f6dcf3e8f12ff1e0f1d8f358f661f850f9e6f876f7f2f547f501f6;
    inBuf[7342] = 256'h36f847fb4bfea300020275025302ce01d8005bff59fd1efb3ef93cf84ef83ef9;
    inBuf[7343] = 256'h77fa7dfb26fc8ffc26fd50fef9ffe001c4035405810676070608b307f1053402;
    inBuf[7344] = 256'h71fc7cf5c5eee0e911e8b6e929ee0bf4cdf948feff003202c0029d035c052808;
    inBuf[7345] = 256'ha40bf90e551131126911560f850c5909f5052f02d8fd3bf91ef591f293f253f5;
    inBuf[7346] = 256'hdbf994fee001af023a01d8fe21fd3cfd66ffdb024e06a1086509e508d6070407;
    inBuf[7347] = 256'hf2068e077e085b09ab0938094d083c075d061d067d0601073907c8068c05f303;
    inBuf[7348] = 256'hb90269022d03a6041b06e206a8069f0557044303a5028f02d3025b0362040606;
    inBuf[7349] = 256'h3f08e50a760d6b0f8510ad100210d20e3e0d600b76099f07f905aa048c037502;
    inBuf[7350] = 256'h8901fa0023017a02f404ff07e80af30cc80dbd0d640d490db00d480e870e1e0e;
    inBuf[7351] = 256'hf60c670b0f0a3a09ec08f708e9089308370815087908a209410be10c3e0e130f;
    inBuf[7352] = 256'h590f4d0ff50e460e5a0d3d0c390bdb0a4d0b600ca50d420ea20de60b84093607;
    inBuf[7353] = 256'hb3050405c704ab047a04810467056e075b0a820dc90f7a10c30f5c0e650dea0d;
    inBuf[7354] = 256'h15106e1321170e1a901bab1b861a99188f169d14d6124c11a70f8a0def0ac207;
    inBuf[7355] = 256'h3c0405019ffe62fd83fdc1feb7001b0396050308560a3e0c860d2c0e320e060e;
    inBuf[7356] = 256'h610e950fb71192144f173419091ac019c118cb172417be165c16581539131210;
    inBuf[7357] = 256'h210c0c08b8049402be011502fe02f303d1048b056606e907260af00c0110c512;
    inBuf[7358] = 256'hc914fa155e163716c915ed1480136011400e540a5006c80282003d00f2013d05;
    inBuf[7359] = 256'h9d09100eb011271449153f15a214db1326139b12fa110711ab0fcc0d970b6109;
    inBuf[7360] = 256'h4f07a005a3044e04a804b305130795084e0a260c2e0e991023135d15f3168817;
    inBuf[7361] = 256'h1417f2156a14c4122e11700f6f0d4f0b1409f2062d05a3033c0221015300f5ff;
    inBuf[7362] = 256'h55006d01090314057307360a830d3d110d155918391a201a03182d14800f180b;
    inBuf[7363] = 256'hac07c20584057406fa07a309d50a500b520b0a0baf0a860a6e0a200a79095a08;
    inBuf[7364] = 256'he00670055004aa0380039703c203f4032404820437051206e1067b0792072907;
    inBuf[7365] = 256'ha0064a068a06a0074e091f0b9e0c420de30cc20b250a5d08ab0609057c034102;
    inBuf[7366] = 256'h9001a801a10214045905dd054805cc030d02aa0017006f005b016d025f030104;
    inBuf[7367] = 256'h510464044004ff03b5035b030003a4021d027a01f700b500da007b0158022b03;
    inBuf[7368] = 256'he40389043305f3059206a506e9057404c6028f014301d3019702a7027f0134ff;
    inBuf[7369] = 256'h66fc0dfaedf831f99cfab2fce5fee4008f02b6033004f1030d03ce01ac000800;
    inBuf[7370] = 256'h09008e004c01f7015b02650219027201680025fff3fd32fd3cfd19fe57ff3400;
    inBuf[7371] = 256'hf8ff58feb6fb12f9a2f73ef8e5fac3fe8802ed045105fa03bc018bff01fe15fd;
    inBuf[7372] = 256'h53fc41fbb6f90cf8ecf6d9f6eaf7c6f9c0fb39fdfcfd38fe5cfecefeafffd600;
    inBuf[7373] = 256'hdd014e02ec01b800e3fee0fc28fbfcf975f973f992f983f926f978f8a5f7e7f6;
    inBuf[7374] = 256'h4af6cef57df570f5ebf532f749f9edfb95fe99009a019b01e000e3ffeffe00fe;
    inBuf[7375] = 256'h01fddefb9dfa8ef908f908f949f950f99bf81cf743f5c9f37af3b7f433f73bfa;
    inBuf[7376] = 256'heafc76feabfec5fd31fc93fa70f9f6f83ef939fa87fbb4fc4cfddffc53fbe7f8;
    inBuf[7377] = 256'h24f6d6f3b0f20af3fef427f8a7fb98fe2100b1ff7efd60fa6cf7cdf51df6f7f7;
    inBuf[7378] = 256'h72fa70fc05fd1ffc6bfad9f859f855f97afb16fe45003001840058fe19fb90f7;
    inBuf[7379] = 256'h79f43ef220f1fdf069f13df286f350f5c2f7bcfa9afda1ff32000effc4fc56fa;
    inBuf[7380] = 256'hb4f892f8ebf9ecfb96fd0dfeddfc67fa8df72df507f44ef48af519f75bf8e5f8;
    inBuf[7381] = 256'hdaf898f86ff8a7f82af98bf993f934f987f809f827f8edf837fa92fb58fc4efc;
    inBuf[7382] = 256'h88fb4ffa3ef9cbf8e9f858f9a2f93df915f86df6acf469f3f7f238f3ecf3b4f4;
    inBuf[7383] = 256'h28f549f53ef539f59bf592f6fcf7c0f99afb20fd2cfebbfed1feacfe6ffeedfd;
    inBuf[7384] = 256'h01fd71fb0ef934f694f3daf1a5f111f37cf50bf8def95ffabaf992f894f75bf7;
    inBuf[7385] = 256'hfaf7f9f8d7f920fa9af99bf8a2f70cf731f70ff83ff95bfaf1fa9bfa60f983f7;
    inBuf[7386] = 256'h66f5acf3c2f2a8f241f33df435f529f658f7f1f81afb9efde2ff6101c201ff00;
    inBuf[7387] = 256'h87ffd4fd21fc9bfa3df9fcf720f7f2f674f78af8c0f977fa7afae0f9e0f8ccf7;
    inBuf[7388] = 256'ha7f615f5e9f256f0f1edc5ecadedc2f06df574fa74fea300e100a2ffd1fd40fc;
    inBuf[7389] = 256'h5cfb58fbfffbcefc55fd30fd21fc6bfa99f830f7a4f6f6f6a9f73bf855f8f9f7;
    inBuf[7390] = 256'ha9f7e3f7bbf8eef9e4fafefa3bfa1cf94af85bf854f996fa63fb2ffbf5f951f8;
    inBuf[7391] = 256'h02f782f6f5f6f7f7e4f86ef989f950f91bf916f91df908f9b8f818f856f7acf6;
    inBuf[7392] = 256'h38f61df65ff6f0f6dbf71df996fa29fcacfdf7fe26006401c302380458056905;
    inBuf[7393] = 256'he2039400dbfbb0f62df20def98ed85ed3aee5defe1f0f2f2c8f535f995fc28ff;
    inBuf[7394] = 256'h5300e5ff6afec4fcaefb90fb4cfc45fdd2fd8dfd70fce3fa6ff98bf86cf8e3f8;
    inBuf[7395] = 256'h97f942fab5faf5fa42fbbbfb3dfca7fcccfc84fcfafb75fb14fbcbfa6dfabef9;
    inBuf[7396] = 256'hbef8b6f718f749f75ef813fafffbc2fd33ff6d0089017502fd02c7027d0119ff;
    inBuf[7397] = 256'hd3fb02f81af48ef0c7ed36ec35eceaed3df1c0f5c7faa8ffc803b1061a08d707;
    inBuf[7398] = 256'hee05db0270ffa5fc5dfbe6fba5fd66fff1ff95fe94fb18f8a2f53ff50ef745fa;
    inBuf[7399] = 256'h99fddaff8400e0ffa2fe8bfd1cfd4cfdadfdc9fd53fd33fca2fa05f9b7f7e3f6;
    inBuf[7400] = 256'h7ff65ff666f6a9f688f78bf9fffc99016a06110a4c0ba109af05fc0055fdfafb;
    inBuf[7401] = 256'h03fd5aff5a019a0193ffecfb27f8daf5edf559f834fc1800da02fc03b103a502;
    inBuf[7402] = 256'h9701e9007d00f3ffe9fe46fd6ffb23fa0cfa6cfb01fe1101a5030c0528055804;
    inBuf[7403] = 256'h45038d026a0295028e02e8019b0022ff40fe91fe2a0076026e041905f9035701;
    inBuf[7404] = 256'h23fe72fb04fa12fa4ffb29fd28ff27012f0344053d07ce08a909a409ec08e807;
    inBuf[7405] = 256'hed062206750592043503600149ff62fd4cfc77fc02fec20028045c0792093f0a;
    inBuf[7406] = 256'h4109f006f8031801ebfec5fdb5fd95fe1b00fc01ed039a05d706a4070b082608;
    inBuf[7407] = 256'h1d08f0079a073607e606de064207df074108f907b906a4046b02d80079006d01;
    inBuf[7408] = 256'h35030a055306d906ce06ac06ca062c078f0792070707140603053f042104a604;
    inBuf[7409] = 256'hb1052907da08960a410c9e0d760ec40e890ee50d110d0a0cb10af708d4067004;
    inBuf[7410] = 256'h350280008dff79ff1e004201bc025704e605480757080b098c09000a960a690b;
    inBuf[7411] = 256'h510c190da50dcc0d900d150d5e0c810bc20a4d0a520afd0a0e0c020d6a0dea0c;
    inBuf[7412] = 256'h760b7b097307be058a04b4030f03910245025a0206033904d705d007f209270c;
    inBuf[7413] = 256'h660e6310b91128128411fb0f1c0e6a0c430bb50a4b0a7909f1079905d4026100;
    inBuf[7414] = 256'hccfe60fe2effd300d202e304cd068008240ad10b960d7b0f5411db12bf139f13;
    inBuf[7415] = 256'h601238107b0da90a35081f064f04d502be016a016902be04de07eb0ad00ce50c;
    inBuf[7416] = 256'h750b6409c6075a07fe07ed0844096e08a606c5048b0361032304110583056505;
    inBuf[7417] = 256'h0205fa04f5050c08dc0ac90d15104c115c116810d80e2a0d9c0b510a4a092408;
    inBuf[7418] = 256'h9706b504b9023501f0003102b604e007b90a7e0c0e0db60c0a0c900b540b0f0b;
    inBuf[7419] = 256'h5d0ae408c60685049802780161010e022f039704fd055107bf083b0aa80bf50c;
    inBuf[7420] = 256'hd80d070e6b0d090c270a4808de063a066706f6066b077207db06e10500056d04;
    inBuf[7421] = 256'h2d041d04ea0375030703f3028503d2047a0605082509b509f1093f0abe0a650b;
    inBuf[7422] = 256'h0b0c5b0c300cad0be90a010a1209fb07a8062e05a3033a023801ad009400d500;
    inBuf[7423] = 256'h2f017401a301ca012c0215037e0427069b073c08c5077e06fd0409043e048905;
    inBuf[7424] = 256'h5407de086d09d0086c07dd05bc046404b0044f05f60564069706b706d306f006;
    inBuf[7425] = 256'h0307d8064a064d05e30351020a017300e9008202cd0411078e089608ff064404;
    inBuf[7426] = 256'h2b018cfe11fdd7fc8cfdb4fedcffe9001202a303d1056f08e00a6b0c830cf40a;
    inBuf[7427] = 256'h2608f104290276001f00e10036029003630464049b033c02a70053ff8cfe6ffe;
    inBuf[7428] = 256'he2fe9fff74004d01340246038c04ce05c406380710077506b40506057904f403;
    inBuf[7429] = 256'h4a035a022a01daffa3feb8fd47fd7ffd6afecfff4b014b023802d90082fee1fb;
    inBuf[7430] = 256'hcdf9fef8acf995fb36feff00750340052406ec058a044802c9ffd4fd1cfdebfd;
    inBuf[7431] = 256'hdbff1102ae03150435038b01bfff46fe4afda7fc15fc74fbeffad5fa62fba5fc;
    inBuf[7432] = 256'h69fe320083011f0208027101b9002900c0ff49ff6ffed5fc63fa5ff756f4fdf1;
    inBuf[7433] = 256'hf0f06bf13ff3e3f5abf81afbfdfc63fe92ffcd00160255035e04fc041805b304;
    inBuf[7434] = 256'hcd036702830032feabfb46f965f75bf63ef6e4f60ef85cf982fa76fb29fc75fc;
    inBuf[7435] = 256'h52fca3fb41fa56f84af67df459f328f3cbf3fff484f61af89ff910fb62fc80fd;
    inBuf[7436] = 256'h41fe9dfec3fee8fe3dffe7ffa300e20035005efe77fb2df85df5a3f353f335f4;
    inBuf[7437] = 256'h8ff5b1f623f7c4f6eef52cf5dff445f540f66df789f86bf9fbf965fad4fa3dfb;
    inBuf[7438] = 256'h94fbc0fb93fb16fb6efabff942f917f938f999f90ffa64fa7dfa28fa3ef9e9f7;
    inBuf[7439] = 256'h56f6b7f482f3f4f2e6f233f397f3b2f387f34ef32ef35ef3edf3a7f46af52af6;
    inBuf[7440] = 256'heff6eaf733f9b0fa45fcb2fdaefe3eff67ff21ff8ffeb8fd8afc22fb8ef9c6f7;
    inBuf[7441] = 256'hecf510f42bf271f009eff5ed5bed41ed8ded5eeec6efaef116f4c6f640f930fb;
    inBuf[7442] = 256'h5bfc97fc1afc37fb2dfa4ef9c8f89af8c9f83af9acf9f9f9e3f936f918f8baf6;
    inBuf[7443] = 256'h5af572f437f47bf40ef588f565f594f451f300f252f1d0f192f371f6daf9f1fc;
    inBuf[7444] = 256'h12ffc7ffe6fed0fc1bfa53f718f5b2f3fdf2caf2cef2bdf2a6f2b6f20cf3d9f3;
    inBuf[7445] = 256'h0ff562f6aaf7b6f85ff9d1f926fa5cfa93fac8fadafae3faebfaccfa8dfa14fa;
    inBuf[7446] = 256'h29f9d7f744f692f41cf326f2b8f1d9f164f21af3f0f3dff4e3f524f79bf816fa;
    inBuf[7447] = 256'h7bfb93fc21fd39fdfbfc76fce4fb5efbc7fa1bfa41f91bf8c4f662f50ef40cf3;
    inBuf[7448] = 256'h7af248f27af2fbf2a3f38bf4c3f542f714f918fbf7fc77fe5eff7bffe5fec1fd;
    inBuf[7449] = 256'h39fc9ffa25f9d4f7c1f6d6f5e8f40ef477f367f341f424f6bff88ffbd1fdd5fe;
    inBuf[7450] = 256'h72fee8fcbbfaa2f816f733f6f6f532f6b2f680f79ff8eff959fb9efc6bfda6fd;
    inBuf[7451] = 256'h4bfd74fc7bfbb2fa44fa52fabbfa22fb38fbc1faaff94af8f0f6eaf574f57ef5;
    inBuf[7452] = 256'hcaf53df6d4f6a0f7daf88afa79fc54feaeff3a000b006cffbefe69fe82feccfe;
    inBuf[7453] = 256'hf0fe7cfe27fd1afbbcf893f638f5fcf4b9f509f75df83bf980f964f950f9b0f9;
    inBuf[7454] = 256'ha8fa0ffc9bfdfdfe17000a01f001c8026c037e03ac02f80098feeefb74f978f7;
    inBuf[7455] = 256'h1cf672f574f50af61cf76af89df97cfafafa38fb88fb32fc50fdcafe53009901;
    inBuf[7456] = 256'h61028b0210020c01b8ff73fea9fdb0fda3fe3100a6014c02bf011b0013fe94fc;
    inBuf[7457] = 256'h2efcd0fccbfd1efe23fd02fba0f826f76bf76af93cfc99fe97ff23fff9fd33fd;
    inBuf[7458] = 256'habfd7afffd014104810579057104e8025201ffff07ff75fe63feddfec6ffe700;
    inBuf[7459] = 256'hea0182029e025402c9012d019f001d00aeff59ff1cffdbfe71fecafdf9fc41fc;
    inBuf[7460] = 256'h07fca1fc16fe250065025504b1058206d906d0068806fb0528054b04af038c03;
    inBuf[7461] = 256'hf603af042f05f504b0038001fffef0fc03fc8efc4efe9900a002a6035e031102;
    inBuf[7462] = 256'h5b0005ffcafef1ff42022905dc07c309b10acc0a890a5b0a460a040a4009ac07;
    inBuf[7463] = 256'h68051c037701f100a201fe022f04a1041d04e2029f01f50037015e020404b005;
    inBuf[7464] = 256'h0507c507ed07a407f506fe05ee04df031203e5027303b50486066208c8097e0a;
    inBuf[7465] = 256'h6f0ad10916098a084b08550866084a08ff078307e8065606ca054805f604e904;
    inBuf[7466] = 256'h430527067007e108400a350b8b0b380b320a9508b206d0045903b002d902a103;
    inBuf[7467] = 256'hbb04ac052f0663067906ba066c077e08c009140b3c0c160da90ddd0daa0d350d;
    inBuf[7468] = 256'h930ce80b540bac0ab3094b086a065f04c3020302530293033405aa06ab071008;
    inBuf[7469] = 256'h0408dd07b3079907ae07ef077a088309f70aa60c570e970f1510c80fb90e1f0d;
    inBuf[7470] = 256'h600bc5098808c0072f07840685050f046e0255015401c1028105c108810b100d;
    inBuf[7471] = 256'h1b0d010ca10aae098409190ae70a690b5f0bb90ab709ae08b407db063e06d105;
    inBuf[7472] = 256'hae050706cb06d307fb08ed09840ade0a0f0b3c0b910bf70b460c620c240c8d0b;
    inBuf[7473] = 256'hbb0abb09af08c407f5065606f5059e0524056a044c03f601e2006e00df004902;
    inBuf[7474] = 256'h4b04710682086b0a580c760e8910141282125911c50e910ba208be062f067b06;
    inBuf[7475] = 256'he606df061d06e204cd03430366031204d60456057f056505540593052406f406;
    inBuf[7476] = 256'hd3076e08a90898084c08fc07df07e707030825081608c7075c07e50683066b06;
    inBuf[7477] = 256'ha6063007f607bb0844096109e208cf075c06bc043b0320027c016601e801d702;
    inBuf[7478] = 256'h17048805de06e907a008fd08260955099a09ef09330a150a68092e088106b104;
    inBuf[7479] = 256'h1c03ef0146011b014101a1013d02f902c4038f042f059405db053306d306d807;
    inBuf[7480] = 256'h1109280ab70a6a0a4809a107d705520444038f021102af014e010a010c014901;
    inBuf[7481] = 256'hac01220291020803b803bb040b0670077c08d1084c080b07790513042b03db02;
    inBuf[7482] = 256'hf0020603d4024202610186001d006500790130030f0589062107910608051603;
    inBuf[7483] = 256'h67018e00bd00a201ab02470325036f0299010f011a01b30189024e03d7031504;
    inBuf[7484] = 256'h1e040004b303270358025201490075ff07ff1dffb3ffa500ca01e302af030d04;
    inBuf[7485] = 256'hfb0390030703950247020c02b001f600c9ff43fea2fc47fb90fabffaf3fb1afe;
    inBuf[7486] = 256'hee000604d906e308d309910951088506a2040403cc01d400d5ff8ffee6fcfafa;
    inBuf[7487] = 256'h29f9daf764f7f6f77ef9b5fb3dfea8009802d4034404f9032f032a022e017000;
    inBuf[7488] = 256'h0000d2ffc7ffb3ff71ffeffe32fe67fdd4fcbbfc44fd5ffeb1ffc2002701ab00;
    inBuf[7489] = 256'h78ff06fed3fc42fc6afc0bfdbdfd25fe08fe70fda3fceefb9cfbd4fb7cfc58fd;
    inBuf[7490] = 256'h1dfe84fe75fe0bfe7afd02fdc4fcb0fc99fc45fc89fb71fa3af937f8c7f71ef8;
    inBuf[7491] = 256'h2bf9b0fa47fc84fd3efe93fec2fe24ffe4ffcf007a016a014c0035fe9cfb17f9;
    inBuf[7492] = 256'h3af74cf631f6a3f64df7f4f79cf85ef944fa4bfb43fcdffcf8fc8cfcbafbd4fa;
    inBuf[7493] = 256'h26fad3f9e7f93ffa9bfad5fad6fa96fa3bfaecf9bef9cef917fa7bfaeffa62fb;
    inBuf[7494] = 256'hc0fb18fc6ffcabfcb7fc77fcccfbc6fa95f96df88ff713f7e3f6e2f6f4f613f7;
    inBuf[7495] = 256'h6ff735f879f933fb0efd82fe35ffeafea6fdd7fb04fa94f8d3f7b9f7eef723f8;
    inBuf[7496] = 256'h16f8a9f711f79bf681f6e9f6bcf7b4f899f93cfa8ffac9fa14fb79fbf4fb4cfc;
    inBuf[7497] = 256'h29fc70fb2ffaa2f840f765f628f67df612f77bf784f729f78ef618f616f6acf6;
    inBuf[7498] = 256'hecf79df955fbc4fc97fd92fdd0fc88fbf9f983f85cf784f6fbf5abf574f56af5;
    inBuf[7499] = 256'ha6f52bf6fdf6f1f7c3f84df978f954f930f93df97ff9f0f951fa4bfad1f9e8f8;
    inBuf[7500] = 256'hb0f785f6abf53af557f5f8f5e9f605f816f9e1f957fa77fa4afa02fabaf97ef9;
    inBuf[7501] = 256'h7af9b9f92cfac9fa51fb68fbe7fac2f91ff882f660f5f2f44ff542f666f77df8;
    inBuf[7502] = 256'h56f9dbf925fa40fa33fa28fa25fa1afa0cfadbf967f9d7f860f831f887f84ef9;
    inBuf[7503] = 256'h25fac0fae7fa90fa0efaaff988f989f964f9d7f8fcf718f786f6a2f662f775f8;
    inBuf[7504] = 256'h99f994fa56fb15fcddfc7afdb9fd54fd28fc82facef866f794f64ef65df6a7f6;
    inBuf[7505] = 256'h18f7a7f76bf851f927fae3fa76fbdafb30fc68fc4bfcc4fbccfa7ef945f873f7;
    inBuf[7506] = 256'h1ef73cf78bf7c8f7f7f736f8adf882f992fa84fb1ffc33fcbffb11fb6afaf0f9;
    inBuf[7507] = 256'hcaf9e0f9f4f9e7f98df9c8f8caf7dbf64df685f6a0f769f98bfb86fdedfeb7ff;
    inBuf[7508] = 256'h070011001100f7ff78ff58fe71fce3f92ff7dcf450f3c6f220f30cf450f5b4f6;
    inBuf[7509] = 256'h19f889f9fbfa53fc8bfd80fe04ff0cff8cfe91fd72fc9ffb76fb36fca5fd21ff;
    inBuf[7510] = 256'h0200cfff89fecbfc5bfbc4fa1ffbf1fb78fc37fc19fb7cf912f85ff782f755f8;
    inBuf[7511] = 256'h71f975fa3afbb7fbf8fb21fc3afc4bfc7cfce0fc80fd69fe86ffa900b9018e02;
    inBuf[7512] = 256'hf302c602e2012c00c9fd08fb4bf805f682f4ddf30ef4f0f45cf63df871fac8fc;
    inBuf[7513] = 256'h0bffea001f0297025d02a001b000c9ff09ff86fe39fe09feeffddafdb8fd82fd;
    inBuf[7514] = 256'h2ffdbdfc3ffcc3fb5cfb29fb39fb92fb34fc05fdd9fd8afe00ff34ff43ff4aff;
    inBuf[7515] = 256'h4eff3affe1fe21fe05fdcafbdbfa9ffa41fba9fc85fe5f00cd019b02be025302;
    inBuf[7516] = 256'h9f01ea0073005f00a200f400fb006c003affa7fd37fc70fb99fb97fc02fe4cff;
    inBuf[7517] = 256'h0b002700daff81ff74ffd7ff8d005e0111028a02da02260390032004b6041c05;
    inBuf[7518] = 256'h180585046103db013700bffeb1fd2cfd27fd81fd03fe89fe05ff7bff0900cc00;
    inBuf[7519] = 256'hbf01c602b8036204b204c104aa0488046c043f04e0034c039c020402c9010902;
    inBuf[7520] = 256'hb4029303460481042c0451032c0210014000edff340004013c02a303d4047005;
    inBuf[7521] = 256'h3905150445025700e6fe7efe68ff78013b04200789090d0b8d0b0c0bbb09f107;
    inBuf[7522] = 256'hf5050a0464020701e7ff06ff62fe18fe53fe17ff5200db01740304059a062e08;
    inBuf[7523] = 256'had09e10a5c0bd60a62095b07680542043a043d05ea069808bc09110a76090a08;
    inBuf[7524] = 256'h1b06f5030402c3007000170190025904f4052007c8071c087608f10887090f0a;
    inBuf[7525] = 256'h360ace09eb08a90754064e05cf0407050c06a6077909260b310c650ce00bd40a;
    inBuf[7526] = 256'h8f0954081307b5054d04fb0225024d029b03e805d0089e0bc80d1b0f7e0f150f;
    inBuf[7527] = 256'h1d0ea30cbe0ab108b406220564048d048405050785088b09d8094409ff078706;
    inBuf[7528] = 256'h4705a404e304d5052c07a208eb09f70af30bda0c9a0d0f0ee40d000da00b150a;
    inBuf[7529] = 256'hd008340823084d086208050839076306e1050d061307a708500aa20b260cbd0b;
    inBuf[7530] = 256'ha50a2c09c507e3069a06dd0686073a08c50832097a09b509070a4e0a750a8b0a;
    inBuf[7531] = 256'h8c0a9d0afb0a9a0b530cf60c260db80cc70b6f0af2089e078406b0053f052105;
    inBuf[7532] = 256'h5905ff05f30618086209970a990b6b0cf90c4b0d8d0dbc0de00df60db60de60c;
    inBuf[7533] = 256'h790b71092c07540560049604ea05c30773098e0ae30aba0aa70afe0aca0bc90c;
    inBuf[7534] = 256'h5f0d120dd20bcb09810795055504dc032104d304b905c106cd07e0081a0a6a0b;
    inBuf[7535] = 256'hc00c080ef40e490ff80ef30d6b0cbc0a15099d076f066b058504da036c035003;
    inBuf[7536] = 256'h9f033b040505f205e206cc07ba089509490ad30a190b1d0bfa0aa90a2d0a8809;
    inBuf[7537] = 256'h96085007da055004f602280207029a02cf035305cf060a08cb080b09f708b408;
    inBuf[7538] = 256'h72085d0866087008640817088c07f2066c061b0609060206ca05490579049303;
    inBuf[7539] = 256'hf602df0267037b04be05d6068607a3073e079206ce052305bb049304ab040a05;
    inBuf[7540] = 256'h9d054b06f7065f074807a20689055404800361030804360560060107d706e805;
    inBuf[7541] = 256'h920457038f026002b30234039703b60389033603fa02f30224037003a2039903;
    inBuf[7542] = 256'h5b030c03e702170395033904c4040105e50489041604b1036a032a03d6025402;
    inBuf[7543] = 256'h9701b600ddff46ff28ff9dff8a00a4017d02ad020502a400eefe6efd94fc95fc;
    inBuf[7544] = 256'h62fdb5fe34009801b5027e03fc0337043a0409049903da02be013c0072fea3fc;
    inBuf[7545] = 256'h25fb51fa5efa34fb84fcdcfdcafe19ffdcfe51fecdfd91fda6fdf8fd62feb8fe;
    inBuf[7546] = 256'heefe08ff06fff4fedafeadfe6efe1afe9dfdfefc53fcc0fb8afbedfbe3fc33fe;
    inBuf[7547] = 256'h6bfffbff93ff3bfe43fc3dfab7f8f0f7f3f790f86cf94dfa0ffb96fbf3fb44fc;
    inBuf[7548] = 256'h9bfc1cfdd3fd96fe32ff65ffebfec9fd3dfc95fa39f96cf823f841f897f8e8f8;
    inBuf[7549] = 256'h2df966f97bf960f9fff83af83df762f6fdf56af6bcf798f985fbfbfc85fd1bfd;
    inBuf[7550] = 256'hfbfb76fa04f9fef77cf78af708f897f8eef8caf8f8f7a6f62ef5dcf301f3b3f2;
    inBuf[7551] = 256'hbcf200f378f31ef426f59ff646f8cef9dafa11fb84fa7af933f80ef73ff6b5f5;
    inBuf[7552] = 256'h6cf54cf517f5bcf433f468f394f2fbf1bef10bf2d6f2caf3b1f45ff5aaf5b7f5;
    inBuf[7553] = 256'ha9f576f52cf5c5f421f46bf3d5f273f276f2e1f277f31ef4baf421f56bf5abf5;
    inBuf[7554] = 256'hc8f5cdf5adf53df593f4ccf3ebf21ef27bf1e5f06ef026f002f02df0baf089f1;
    inBuf[7555] = 256'h9df2e6f333f584f6bdf784f8a5f8ecf73df6faf3b8f1f2ef1def40efe3efa0f0;
    inBuf[7556] = 256'h25f140f13af15cf1a9f120f292f2b6f2abf2b0f2e6f27af34bf4eaf423f5ecf4;
    inBuf[7557] = 256'h54f4c3f384f389f3c8f305f4eaf371f3a3f27ef145f043efa9eedaeefbefc3f1;
    inBuf[7558] = 256'hd1f387f544f6f2f5d5f458f31df274f136f134f123f1c0f035f0bfef7eefadef;
    inBuf[7559] = 256'h56f048f17af2cff306f514f6e0f63ff749f712f793f6f4f541f562f46ef36bf2;
    inBuf[7560] = 256'h3ff10bf0e5eedbed40ed58ed2deec5efd1f1bbf329f5edf50bf6f5f50ef65ff6;
    inBuf[7561] = 256'hd4f611f7a3f695f538f401f385f2f9f209f446f52af653f6e8f545f5b3f480f4;
    inBuf[7562] = 256'ha2f4c3f4b8f464f4c3f325f3caf2c3f229f3e5f3b8f490f553f6ddf643f792f7;
    inBuf[7563] = 256'hc6f707f85bf8a4f8ddf8f2f8c4f878f831f8f7f7e3f7e0f7b1f750f7c0f617f6;
    inBuf[7564] = 256'h98f564f561f580f59ef5a7f5d2f557f640f783f8cef9acfaf1faa6fa03fa7df9;
    inBuf[7565] = 256'h58f98cf900fa6ffa9afa8afa57fa1cfa06fa16fa29fa2afaf1f95cf989f8acf7;
    inBuf[7566] = 256'h11f723f716f8c5f9d6fbaefdb3feb1fec2fd46fccffac2f943f95af9e1f9a8fa;
    inBuf[7567] = 256'h9afb90fc56fdc5fdb3fd0ffd08fce3faf3f990f9dcf9c4fa19fc81fda1fe4fff;
    inBuf[7568] = 256'h81ff5bff28ff16ff2cff4eff3cffc3feeefdeefc12fca9fbcefb67fc4dfd4efe;
    inBuf[7569] = 256'h54ff69008801930254037d03df028c01d0ff21fef2fc78fca6fc3cfde1fd5afe;
    inBuf[7570] = 256'ha1fecffe19ffb1ffa300e00144039604ac056d06c706c4067706e30513050304;
    inBuf[7571] = 256'hae02270198ff35fe48fd05fd78fd94fe2300d2015d038a043a05810590059a05;
    inBuf[7572] = 256'hd5054f06e6067807d907ed07c5076e07e606320643051604db02cd0123010d01;
    inBuf[7573] = 256'h830155025c036c046b0563064d071a08cc084d098a0987093009730862071506;
    inBuf[7574] = 256'hbe04c3036703d3031305e906f408e30a540c050df90c3e0c040baa096c087507;
    inBuf[7575] = 256'hee06c306d106ff061507e0065b0680057604a4035b03d6033e055d07de09800c;
    inBuf[7576] = 256'hed0eee107412491340136412ca10c40ee10c750b900a0a0a5c090d081106a103;
    inBuf[7577] = 256'h5401f8ff03008f0171040d08bd0b0f0f95111d13c513a713ff1234126a11a710;
    inBuf[7578] = 256'hee0ffc0eac0d250c8d0a300966082b085508c9084609bf09620a2c0b0d0cfd0c;
    inBuf[7579] = 256'hb70d190e500e6f0e9b0efc0e5b0f780f3c0f830e6d0d610c960b3c0b840b480c;
    inBuf[7580] = 256'h5c0daf0ef90f0011b211ce113d112b10b00e0a0d9e0b850acf099709b209080a;
    inBuf[7581] = 256'ha70a640b1f0cdd0c700ddb0d600e140f10106411b5129d13e4134513ce11e50f;
    inBuf[7582] = 256'hce0de10b7e0aac096909b709470add0a6e0bd60b2e0cc20c920d890e8c0f3910;
    inBuf[7583] = 256'h5f102a10b50f400f160f1a0f270f3b0f2a0ff40ebd0e5e0eb60dcd0c910b340a;
    inBuf[7584] = 256'h25098f0896085309850afb0ba50d390f81106811ac115311a910db0f190f850e;
    inBuf[7585] = 256'hd80ddb0ca00b430a2f09e9087809a20a090c120d790d6e0d240dee0c0b0d460d;
    inBuf[7586] = 256'h630d4c0de10c480cd60b900b6f0b680b340bc30a460ad2099509c509410af40a;
    inBuf[7587] = 256'hdc0bc80ca20d660ecd0ea50eea0d8b0ccc0a2909ee0757077707f5077d08e208;
    inBuf[7588] = 256'hf508d008bd08ce081a09b709730a370bf70b700c770c010cf10a7609fb07cb06;
    inBuf[7589] = 256'h340662061b071208050990098c090a090e08dd06dd05490559051d0641076708;
    inBuf[7590] = 256'h450990095609e40864080508db07b1076a070d0792061f06e605d805eb051006;
    inBuf[7591] = 256'h0c06d1057205f60492048504d40474053d06cc06e30679069f05af041104eb03;
    inBuf[7592] = 256'h3d04db046305a205990557051205f004d904ac044d04a203ce0214029d018c01;
    inBuf[7593] = 256'he0016402f3027a03e103330479049a0488043a04a103de02230295015d018601;
    inBuf[7594] = 256'he8015702a702ac0272021f02d701be01d301e201b60123011800c8fe85fda0fc;
    inBuf[7595] = 256'h63fce2fcf2fd54ffb400c1015f028d0262021102bb016e012f01f100a1003a00;
    inBuf[7596] = 256'hb3ff03ff3afe69fdabfc2efc00fc14fc4cfc78fc7cfc72fc80fccdfc63fd0dfe;
    inBuf[7597] = 256'h7cfe7cfefefd3cfd92fc43fc64fcdbfc64fdc9fdf6fde0fd92fd1efd84fcd7fb;
    inBuf[7598] = 256'h3cfbc9fa91fa93faa5faa8fa8ffa58fa19faecf9c8f9a9f990f979f97ef9b7f9;
    inBuf[7599] = 256'h18fa8cfaf3fa20fb18fbf9fad7facffadefad4fa93fa15fa5ef9aef846f839f8;
    inBuf[7600] = 256'h84f8f2f829f9fcf86ef8a5f702f7d4f61ff7c4f775f8cdf8b6f84cf8c0f762f7;
    inBuf[7601] = 256'h5cf78ef7dbf71cf82af81df811f8f8f7cff772f7acf68ef552f441f3cbf230f3;
    inBuf[7602] = 256'h51f4ecf58cf7a4f802f9b1f8e4f712f797f680f6c1f618f725f7d7f644f68ff5;
    inBuf[7603] = 256'h0af5d2f4b0f471f4dbf3c8f285f182f006f04cf028f118f2cef22bf344f391f3;
    inBuf[7604] = 256'h6cf4c6f569f7cff85cf9ecf8a7f7e8f557f468f327f380f30df43cf4d3f3ccf2;
    inBuf[7605] = 256'h52f1f7ef34ef29efd6efdaf0a2f1f6f1d0f14ff1e6f0d8f019f1a5f150f2dbf2;
    inBuf[7606] = 256'h5af3d4f334f48df4cff4d2f4b7f48ef44ef416f4d7f35ef3b5f2e2f1e6f00cf0;
    inBuf[7607] = 256'h86ef5cefb2ef72f046f105f26ff249f2c4f120f18ef063f0a0f0f7f041f151f1;
    inBuf[7608] = 256'h19f1f9f042f1fff12af35df403f5eef42df408f325f2e7f13ff2fff2a5f3a9f3;
    inBuf[7609] = 256'h06f3ebf1a9f0c8ef83efb2ef38f0cdf026f15ef189f1a8f1e4f130f25cf279f2;
    inBuf[7610] = 256'h85f26ff260f25af23ef22df22ff23cf281f2f9f26cf3d0f304f4e7f3b0f385f3;
    inBuf[7611] = 256'h64f36cf37af34ef3eef260f2acf120f1dcf0d6f024f1aff143f2e8f284f3eef3;
    inBuf[7612] = 256'h3cf46df472f46ef458f408f48af3dbf2fff14cf1fbf018f1bbf1aff29df36af4;
    inBuf[7613] = 256'hfff454f5a9f512f67af6e7f632f729f7e5f678f6eef585f545f509f5cef46cf4;
    inBuf[7614] = 256'hc5f308f367f208f229f2bbf272f321f48cf49af495f4c2f44bf556f6b4f701f9;
    inBuf[7615] = 256'h01fa79fa4bfaadf9c9f8c2f7dbf62bf6b0f580f58df5baf517f6a1f64ef737f8;
    inBuf[7616] = 256'h3ef923fac0faddfa61fa86f98af8a4f70df7b7f66ff624f6c7f568f551f5b0f5;
    inBuf[7617] = 256'h90f6f3f798f927fb6afc27fd47fdf1fc54fca7fb35fb1dfb5afbe3fb81fceffc;
    inBuf[7618] = 256'h0afda8fcc0fb87fa3cf928f899f79ff714f8c9f87af901fa70fae2fa6afb18fc;
    inBuf[7619] = 256'hcafc5bfdc7fd10fe48fe89febefec5fe8ffe1afe87fd1afdf6fc20fd86fdf8fd;
    inBuf[7620] = 256'h59feadfefafe43ff80ff83ff27ff6bfe68fd5efc9efb54fb8ffb41fc38fd4bfe;
    inBuf[7621] = 256'h5cff4a00030179019b016d010d01a1005e007000d90085014802e50237032a03;
    inBuf[7622] = 256'hb902ff0120014300a0ff63ff99ff3a001201d20144024c02f901880139013101;
    inBuf[7623] = 256'h86012502e702b0036304e2042a0534050605c70497049104cd043b05b0050406;
    inBuf[7624] = 256'h04068e05b40497037402a10150018c01470238031604c40436058805f6059006;
    inBuf[7625] = 256'h4a071208b40814093e093a090f09d1086808c307f5060e062e05900440043904;
    inBuf[7626] = 256'h7e04ee04710504068106c606d006920631060a0661065f070209e20a7d0c7d0d;
    inBuf[7627] = 256'ha50d0e0d1a0c0a0b0b0a37096b089807db063f06da05c505db05fc052c065f06;
    inBuf[7628] = 256'ha4062607d907ab089c097e0a370bcd0b220c320c240c040cf20b1b0c610c970c;
    inBuf[7629] = 256'ha00c440c7f0b960aaf09f8089a0866083208fd07b7078307b1074a0846098c0a;
    inBuf[7630] = 256'hb80b840ce80cdb0c8b0c4a0c220c140c220c170ce80bbb0b930b880bba0b010c;
    inBuf[7631] = 256'h430c7e0c850c4b0ce70b410b690a9909e6087d0892080709b509860a360bb10b;
    inBuf[7632] = 256'h180c660cb10c220d9f0d1a0e9b0ef00e020fe60e8a0e060e940d280db70c3a0c;
    inBuf[7633] = 256'h6a0b300abf083e0709069205e405ef068c08450ac50bf50cad0d030e3a0e5d0e;
    inBuf[7634] = 256'h820ec20eec0edf0e9f0e0e0e450d880ce30b680b250bdd0a720af90972090809;
    inBuf[7635] = 256'hfd0835098d09e709010adb09bb09c4091c0ad80aa90b4e0cb30cb60c780c400c;
    inBuf[7636] = 256'h0c0ce10bcc0baa0b880b940bc10b010c470c460ce30b3b0b560a5f099208e107;
    inBuf[7637] = 256'h51070607f5063607e207c608b409940a330b980bf60b4a0c930cd20ccb0c6e0c;
    inBuf[7638] = 256'hdb0b120b340a6a09a408ea076607180714076e07ea075a08ae08cd08d9081509;
    inBuf[7639] = 256'h7f09090a980adc0abf0a680af2098a0955091f09bf082e086707a7064d066e06;
    inBuf[7640] = 256'h0207d9078008b1086a08bc07fb0690069b0622070308d90855095709ca08e507;
    inBuf[7641] = 256'h090773064e069e0612075e075b07f1065106d00590059f05ee05360654065106;
    inBuf[7642] = 256'h2e060706f705e405c305a1057b056d059005c905ff0521061c0606060d063106;
    inBuf[7643] = 256'h640687065806c405e504dc03eb024f0212023a02bc0266030e048e04b3048104;
    inBuf[7644] = 256'h2504ce03b90303047e04ef042005f40493044604340461049b048604ed03dc02;
    inBuf[7645] = 256'h8a015e00b2ff9fff1700ee00de01c1028003010440043f040004a2034603f702;
    inBuf[7646] = 256'hb5026f0205027c01f30092008300d0004d01c6010a02ff01bc0165011201d000;
    inBuf[7647] = 256'h91003f00e2ff8eff60ff73ffc3ff3300a200ef000a01fc00ce0087003200d9ff;
    inBuf[7648] = 256'h8cff6aff87ffe6ff75000401610170012b01ad002700b9ff71ff46ff16ffc4fe;
    inBuf[7649] = 256'h4bfeb0fd11fd92fc45fc33fc5efcb6fc35fdddfda3fe7bff5500040165016001;
    inBuf[7650] = 256'he60010000eff0ffe40fdbafc6bfc3bfc15fceafbcbfbd7fb17fc89fc11fd7afd;
    inBuf[7651] = 256'ha9fda0fd6efd45fd4bfd7dfdcdfd1efe45fe3efe19fedffda3fd6cfd1cfda8fc;
    inBuf[7652] = 256'h12fc58fba4fa24faf0f91ffaadfa6dfb39fce8fc4bfd60fd38fde4fc90fc5ffc;
    inBuf[7653] = 256'h4bfc54fc69fc66fc47fc12fcbffb67fb19fbcffa9ffa9cfabdfa06fb67fbadfb;
    inBuf[7654] = 256'hc2fba6fb5bfb17fb08fb2afb73fbc2fbdcfbc0fb85fb3bfb0bfbfffaf3fadcfa;
    inBuf[7655] = 256'hb5fa72fa33fa12fafff9fdf908fa0afa1dfa5bfab7fa2ffba5fbdafbc0fb5cfb;
    inBuf[7656] = 256'hb4fa05fa84f93af940f992f905fa92fa27fb9afbe4fbf6fbaefb1afb52fa5ff9;
    inBuf[7657] = 256'h7af8cdf758f735f763f7bef744f8e7f87ff90efa90faeafa2dfb5efb65fb4ffb;
    inBuf[7658] = 256'h24fbd6fa85fa48fa11faedf9d1f996f948f9f6f897f84df821f8f3f7d0f7bdf7;
    inBuf[7659] = 256'hb0f7d0f730f8b5f85df90efa8efadafaeafaa6fa2cfa9bf9faf87ef847f842f8;
    inBuf[7660] = 256'h74f8c3f8f7f812f91bf90ef915f943f979f9b3f9d7f9b5f95ef9e8f85ef8f3f7;
    inBuf[7661] = 256'hc2f7aef7b7f7caf7c2f7bbf7d0f701f86bf807f9a0f92bfa94fab6faa5fa6dfa;
    inBuf[7662] = 256'hfff982f90cf997f83ef800f8b4f765f71bf7d8f6d0f619f791f727f8aff8edf8;
    inBuf[7663] = 256'hf1f8daf8b9f8c4f80df96ff9e3f947fa61fa2dfaa8f9cbf8d5f705f77cf66cf6;
    inBuf[7664] = 256'hcef658f7e3f742f855f84af84df866f8aaf802f934f93ef924f9e2f8a7f883f8;
    inBuf[7665] = 256'h5ff843f82ef811f814f84ef8aaf827f99df9cef9baf96bf9e8f86cf80ef8bcf7;
    inBuf[7666] = 256'h7df743f7f3f6a9f679f65ef676f6c4f627f7a7f737f8b4f82df9a4f90bfa7cfa;
    inBuf[7667] = 256'hf4fa46fb61fb28fb81fa9ef9baf8fbf78ef764f73ef706f7b8f663f64ff6a5f6;
    inBuf[7668] = 256'h49f71cf8d8f836f945f930f91ff953f9d3f96afaf2fa38fb0efb8afac5f9d3f8;
    inBuf[7669] = 256'hecf72df79cf65af66ff6c7f669f73bf809f9bcf92ffa43fa12fac3f976f96af9;
    inBuf[7670] = 256'hb2f92dfabcfa24fb29fbd0fa31fa6ef9c9f861f829f81ef82bf836f858f8a0f8;
    inBuf[7671] = 256'h05f987f907fa59fa80fa89fa81fa8cfaa6faa6fa7bfa1bfa8ef912f9d5f8dff8;
    inBuf[7672] = 256'h30f9a3f908fa5afa9dfacefafffa29fb35fb31fb26fb19fb1cfb21fb04fbc2fa;
    inBuf[7673] = 256'h5efae5f987f958f949f952f95af952f953f973f9b8f930fac7fa60fbf9fb8bfc;
    inBuf[7674] = 256'h0bfd7ffdd8fdfffdf3fdacfd29fd80fcbdfbebfa2dfa95f92ef90cf92af979f9;
    inBuf[7675] = 256'hfcf9acfa7cfb66fc45fde8fd32fe13fe98fdfafc67fcfcfbc0fb9afb69fb2cfb;
    inBuf[7676] = 256'hf1fadafa0ffb98fb59fc2efde2fd57fe96feb0febdfed0fedffed4fea3fe47fe;
    inBuf[7677] = 256'hcefd58fdf7fcb0fc7dfc47fcfefbabfb61fb3dfb64fbdcfb9efc92fd8dfe6aff;
    inBuf[7678] = 256'h110071008c0073003300e1ff91ff49ff09ffd0fe8dfe3cfedffd80fd36fd1bfd;
    inBuf[7679] = 256'h35fd82fdeefd59feb7fe07ff59ffc3ff5000ed007701c0019b010501170008ff;
    inBuf[7680] = 256'h1dfe93fd82fde4fd8ffe46ffe0ff4c009600e4005301e0017202d602de027f02;
    inBuf[7681] = 256'hd001fa003b00afff59ff2eff14fff7fee3fee7fe18ff91ff50003d013d022303;
    inBuf[7682] = 256'hc70323043a041a04e2039203190373029b01a600ccff39ff00ff28ff8afffeff;
    inBuf[7683] = 256'h80000e01b40185026b033e04e6044c057105790572055a052f05d4043e048a03;
    inBuf[7684] = 256'hcf022902b7016b0130010801eb00e40018018a0130020103d303830414057b05;
    inBuf[7685] = 256'hbf05fc052b063e063106e90559059c04c703050393028402da028c0361042305;
    inBuf[7686] = 256'hb90508061006fb05d505a9058b0560051705ba044604cb03760351036303bc03;
    inBuf[7687] = 256'h4504e804a80566060b079e070408340841082108d6077b070b078e062506cc05;
    inBuf[7688] = 256'h84055a053005f304b204660421040d042c047d040f05c605950685076f083309;
    inBuf[7689] = 256'hc409f809c6095409b40803086b07e0065e060106c905c3050d068206fa066207;
    inBuf[7690] = 256'h8f0782076c075a075f079507dd0722086a08920885084e08d9073c07b9066e06;
    inBuf[7691] = 256'h7506df067007f5076608b008ea084209a409f309220a0e0ac1097a093f090b09;
    inBuf[7692] = 256'hd208510872076d067705e4040305be05de0631085d09370acd0a0f0b030bd00a;
    inBuf[7693] = 256'h700af9099f095f0936092a090d09cb0881082c08e607d707eb0715085f08ac08;
    inBuf[7694] = 256'hf8085a09b209eb090a0aed0997093409c7086508380831085108ac081b098009;
    inBuf[7695] = 256'hd209df09a30952090009d608fc0849099009c009b1096e0933090809f6080609;
    inBuf[7696] = 256'h0b09ed08c708910861085e0874089b08dd081b094b097f099b099e09a709a909;
    inBuf[7697] = 256'hae09cc09de09cb099a093109a2082508c0077d076e07690760076e078e07d107;
    inBuf[7698] = 256'h5408ed087609df09fb09c90979091409b60885086f087208a308e50823095809;
    inBuf[7699] = 256'h4d09ee0859089e07f20698069206d0064707bd07190864088a08840863081408;
    inBuf[7700] = 256'ha6074d0714070c0740078107b207da07e907f007090817080308d3077b071807;
    inBuf[7701] = 256'he206db06f9062f0745072907f506b00675066206610663067206770672067606;
    inBuf[7702] = 256'h690643061306d2058e0568055a0561058a05c00504066506ca061e0751073d07;
    inBuf[7703] = 256'hde065c06d105690549055c057f05990580052e05c4045004e703a4037c036d03;
    inBuf[7704] = 256'h8603ba030104550491049f04890453041e0415043a048904f6045e05aa05d705;
    inBuf[7705] = 256'hcf058a0512056a04ac03050388023e0225021a020a02f701df01cf01d601ee01;
    inBuf[7706] = 256'h15025802bb024303e8037c04cd04ba0438046a039502ea018701660163015c01;
    inBuf[7707] = 256'h49012d011c0127014a017801a601c801e001f9011202280231021c02e1018401;
    inBuf[7708] = 256'h0d0188000b00a4ff67ff64ffa3ff1a00b3004501a901c301900122019c001f00;
    inBuf[7709] = 256'hc2ff89ff6fff6bff75ff87ff97ff97ff79ff3bffe7fe9bfe77fe90fee6fe65ff;
    inBuf[7710] = 256'hebff5c00a600bb009c004900c5ff26ff8afe10fed2fdd3fdf8fd20fe2afefefd;
    inBuf[7711] = 256'ha5fd32fdb5fc4bfc0dfc0bfc5bfc06fdeefdeefec8ff39002d00aeffddfefefd;
    inBuf[7712] = 256'h43fdbefc79fc69fc73fc92fcbefce0fcf3fceafcb3fc62fc0cfcc1fb9efba6fb;
    inBuf[7713] = 256'hbffbdbfbecfbdffbcafbbdfbbafbd1fb01fc33fc6bfca5fccdfce8fcf0fcd3fc;
    inBuf[7714] = 256'ha1fc60fc05fc9dfb28fb98fa0bfa9ff961f96df9b5f9fff929fa1bfacdf97af9;
    inBuf[7715] = 256'h5af984f907facafa8bfb30fca3fcc7fcabfc56fcbafbf9fa31fa6ef9daf882f8;
    inBuf[7716] = 256'h49f831f82ef826f82df84bf86bf89cf8def81ef970f9d6f92bfa6efa8afa63fa;
    inBuf[7717] = 256'h14fabdf962f92af917f905f9f6f8e2f8b1f87cf84cf80af8c4f780f72ef7f4f6;
    inBuf[7718] = 256'hedf60ef76af7f1f769f8c7f8fcf8edf8bcf884f83df806f8e7f7c4f7b4f7bff7;
    inBuf[7719] = 256'hcaf7e8f712f822f821f811f8daf797f756f700f7b5f683f65af657f67af699f6;
    inBuf[7720] = 256'hb8f6d1f6cff6dbf610f758f7baf71bf83df827f8e6f77bf71cf7e3f6b3f692f6;
    inBuf[7721] = 256'h77f63bf6fff5dcf5caf5edf54bf6b9f634f7a4f7d4f7cbf78ff714f791f62ef6;
    inBuf[7722] = 256'he7f5ddf50ef649f68cf6c9f6d5f6c4f69ff652f604f6d2f5b3f5cdf528f694f6;
    inBuf[7723] = 256'h0bf774f79df79af780f746f714f7f9f6d6f6c2f6c3f6bcf6c0f6c7f69ef64cf6;
    inBuf[7724] = 256'hdbf547f5d5f4b7f4e5f46ef535f6f0f68df7fff726f823f80bf8d2f7a0f78bf7;
    inBuf[7725] = 256'h7cf784f799f78af763f72cf7d7f68bf655f615f6daf5b1f58ff5a8f515f6b3f6;
    inBuf[7726] = 256'h75f730f89ff8c8f8bff884f844f811f8cef78bf754f719f7fbf607f718f734f7;
    inBuf[7727] = 256'h57f766f783f7c3f70ff873f8e0f826f948f94bf91ff9e5f8b0f86df82df8f4f7;
    inBuf[7728] = 256'ha5f758f720f7f6f6fcf640f79df70ef87ff8c5f8f2f81ef948f991f901fa6afa;
    inBuf[7729] = 256'hc2faf6fae2faa0fa48fadbf978f92ff9e3f89ef85df809f8b8f782f767f78bf7;
    inBuf[7730] = 256'h02f8b3f89af99dfa80fb31fca3fcc0fc9efc56fce3fb60fbddfa4efac9f960f9;
    inBuf[7731] = 256'h0cf9e3f8f0f81df971f9e6f959fac8fa29fb61fb7ffb95fba8fbd4fb23fc77fc;
    inBuf[7732] = 256'hbffce1fcbafc58fcd8fb4ffbe9fabcfabafaddfa1bfb58fb9dfbf0fb47fca7fc;
    inBuf[7733] = 256'h05fd42fd56fd43fd06fdbcfc83fc5ffc5afc6dfc7dfc87fc8dfc8efc9efccafc;
    inBuf[7734] = 256'h08fd57fdabfdeafd0efe18fe05fee6fdcffdc6fdd5fdf8fd1afe2ffe30fe19fe;
    inBuf[7735] = 256'hf6fdd3fdadfd88fd66fd4bfd51fd8bfdfcfd94fe2bff92ffaeff81ff29ffd3fe;
    inBuf[7736] = 256'ha4fea9fed9fe23ff6dffadffe0ff02000e00ffffd1ff89ff37fff1fed0fee5fe;
    inBuf[7737] = 256'h32ffa7ff25008800af0091003e00d8ff8bff75ff9affe4ff330069007c007c00;
    inBuf[7738] = 256'h7d009000be00fb00380170019d01c701f601230240023d020902a0011a019300;
    inBuf[7739] = 256'h2f0012004000a9003501b6010e02370234021a020e021c0246028b02d1020303;
    inBuf[7740] = 256'h1f031b03f902cc02990264023f022a02260243027602ae02eb0217032c034103;
    inBuf[7741] = 256'h5d038703cd0313043b0440041504ca038d036b036b038e03b103bb03b603a103;
    inBuf[7742] = 256'h8d039b03c203f50331045c046b0475047c048504a804d504fc04240537052d05;
    inBuf[7743] = 256'h1e050a05fa040c0532055c058a059c0580054e050905c504ac04b704d6040c05;
    inBuf[7744] = 256'h3a05520571059305ba05f7052d064a066006670668068506a906bf06ce06be06;
    inBuf[7745] = 256'h8c065d062e06fb05db05be05a705be0501066206e3064f0783078e076f073707;
    inBuf[7746] = 256'h1407fb06df06d206c306b406c706f0061e075c078d07a707c707dd07dd07d907;
    inBuf[7747] = 256'hb9077c074e072e0721073e0764077c079a07b107c207ec0717082f0846084908;
    inBuf[7748] = 256'h3a083f08480846084b083a081008f307e007d607f00712082b0850086a086c08;
    inBuf[7749] = 256'h6b0852081b08f107d907dd071c087108b608ec08f108c808a40886086f087508;
    inBuf[7750] = 256'h7e088008a208d80819096b0998097c092e09b3082d08dc07ba07b107c307cc07;
    inBuf[7751] = 256'hc407d707030841089c08e8080d0926092e0930094d096d0979097e0962091f09;
    inBuf[7752] = 256'hd3087208fe07a6076e076407aa0719088a08ed081709fe08d10896085b084008;
    inBuf[7753] = 256'h2e081c082408380856089008c508dd08e708cf089e087908570837082c081e08;
    inBuf[7754] = 256'h0608fb07eb07d207c907c007b507c507e30706083e086d0883088c0875083c08;
    inBuf[7755] = 256'hfe07b30761072a070607f9061c0754079007d50705081b0835084d0862088108;
    inBuf[7756] = 256'h82085008f7077507e10670062406fd0505061d063e067806bd0603074d077907;
    inBuf[7757] = 256'h7c0772075c0751076a079307b607cc07b90777071d07a7062106a90546050905;
    inBuf[7758] = 256'h0e0545059905020657068e06b706cd06d606de06cf06a4066d062b06e905b905;
    inBuf[7759] = 256'h88054d051105d004a104a504d7042a058e05db05030612060706ef05d505a705;
    inBuf[7760] = 256'h60051305c4048d0482049304ac04be04b1048c046504420429041c040904ed03;
    inBuf[7761] = 256'hda03d403e6031504490476049604a0049b048e046c043204e6038e0341031703;
    inBuf[7762] = 256'h0e031c032b032103fb02ca029b0281028902a702d6020f03420365036e034c03;
    inBuf[7763] = 256'h0103a0023e02fb01e401f0010d02280230022d02290223021a020202cf018b01;
    inBuf[7764] = 256'h4d0127012d0158018e01b601bd019b0162011d01d7009b006d004f004f006b00;
    inBuf[7765] = 256'h9d00d800060116010e01f700e000d400c6009d004d00d0ff3dffbdfe6efe5efe;
    inBuf[7766] = 256'h87fec7fefffe29ff41ff56ff7cffabffdbff020010000600f0ffc9ff96ff5cff;
    inBuf[7767] = 256'h12ffc0fe77fe34fefbfdccfd98fd62fd3bfd25fd29fd46fd63fd73fd76fd69fd;
    inBuf[7768] = 256'h60fd6ffd8efdb6fde0fdf3fdf4fdedfdd6fdb6fd8ffd54fd0dfdccfc8dfc5efc;
    inBuf[7769] = 256'h42fc25fc0afcf8fbeefbf8fb1efc47fc69fc7cfc70fc4ffc2cfcfffbcffba1fb;
    inBuf[7770] = 256'h65fb2afb03fbeafae8faf9fa00fbfbfaf3fae7faeffa19fb50fb8bfbc1fbd8fb;
    inBuf[7771] = 256'hdafbd4fbb9fb8cfb4cfbe5fa69faf5f98cf946f922f902f9e1f8c8f8b7f8d1f8;
    inBuf[7772] = 256'h2bf9aef94cfaeafa5dfba5fbc8fbb7fb7dfb1bfb7efac1f908f961f8f1f7c1f7;
    inBuf[7773] = 256'hb4f7c4f7eaf713f850f8a8f8fef84ef98df9a7f9b2f9c6f9daf9f8f91afa1cfa;
    inBuf[7774] = 256'h06fadcf991f93af9daf860f8e3f774f717f7e5f6e6f6faf621f756f789f7d0f7;
    inBuf[7775] = 256'h35f89bf8fdf84bf969f96ef970f969f96af968f93cf9ecf883f802f890f73cf7;
    inBuf[7776] = 256'hf5f6c4f6abf6a3f6c9f629f7a6f731f8abf8e3f8e3f8bcf876f838f813f8f4f7;
    inBuf[7777] = 256'he5f7e1f7cdf7b6f79af765f72ef706f7edf6fef63df788f7dcf72ef869f8a4f8;
    inBuf[7778] = 256'he8f818f933f922f9c9f843f8b6f735f7eef6e8f600f72ff762f77cf792f7a9f7;
    inBuf[7779] = 256'hb1f7baf7c4f7c0f7c5f7daf7ecf705f81bf818f80ef805f8f5f7f4f702f808f8;
    inBuf[7780] = 256'h19f838f857f888f8c3f8e6f8f2f8def89ff855f814f8dcf7c2f7c2f7c2f7caf7;
    inBuf[7781] = 256'hd7f7d7f7ddf7e7f7e6f7ecf7fcf70ff839f879f8b2f8e8f80df90ef905f9fff8;
    inBuf[7782] = 256'hfaf80bf92af93af942f93bf91af9f9f8ddf8b6f895f876f84ff83af83ef850f8;
    inBuf[7783] = 256'h80f8c6f809f952f994f9b8f9c7f9bdf992f966f949f93af947f961f96bf96af9;
    inBuf[7784] = 256'h60f94df951f96ff992f9baf9d5f9d5f9d2f9daf9e9f90efa3afa52fa5efa5cfa;
    inBuf[7785] = 256'h47fa37fa2cfa1afa0dfa01faedf9e2f9ddf9d4f9daf9f1f914fa56fab1fa0cfb;
    inBuf[7786] = 256'h62fb9ffbb2fbadfb97fb70fb4bfb20fbe2faa2fa64fa2cfa17fa24fa49fa8afa;
    inBuf[7787] = 256'hd8fa22fb6dfbb1fbe1fb08fc25fc38fc56fc80fcaafcd4fce9fcd5fca2fc55fc;
    inBuf[7788] = 256'hfcfbb2fb80fb62fb5efb67fb6ffb7afb82fb84fb92fbaffbdefb2cfc91fcfefc;
    inBuf[7789] = 256'h70fdd7fd26fe65fe8dfe97fe89fe5dfe12febefd6cfd29fd06fdfdfc00fd09fd;
    inBuf[7790] = 256'h0afdf9fce2fcc4fca9fca4fcbafcf1fc50fdc6fd41feb2fe01ff27ff2fff24ff;
    inBuf[7791] = 256'h18ff1eff36ff56ff77ff86ff7aff5bff2bfff6fecdfeb2fea7feb0fec5fee3fe;
    inBuf[7792] = 256'h0bff32ff4fff5eff55ff35ff0affdefec5fecffefefe50ffbcff2d009800f200;
    inBuf[7793] = 256'h300152015e0155013f0127010d01f700e800db00cd00bb009d0076004d002a00;
    inBuf[7794] = 256'h1c002f005e00a500f5003901690180017d0171016701640174019801c8010502;
    inBuf[7795] = 256'h47028102b202d202d902c902a3026b0232020402ea01f00110023b0267028802;
    inBuf[7796] = 256'h91028d0283027802780285029802b902e3020f03420373039603af03b803b103;
    inBuf[7797] = 256'hac03aa03ab03b603c103c303c303bf03b503b303b303b003b203b503b903cc03;
    inBuf[7798] = 256'heb03100440046a0482048c048604700462045c0462048004a904d004f5040a05;
    inBuf[7799] = 256'h09050305fb04f5040205150523052f052e0521051e052605370557056f057005;
    inBuf[7800] = 256'h620542051d050e051605300561059105b205cd05df05f00517064f068e06d406;
    inBuf[7801] = 256'h05070f07fc06c50675062a06e405a205720545051b0508050e0531057e05df05;
    inBuf[7802] = 256'h4006a006ea061e0752077e07a307cb07e307e507e207d107b207930763071b07;
    inBuf[7803] = 256'hce0679062a06fa05e205db05ec05ff0513063d067606bf0622078307d0070b08;
    inBuf[7804] = 256'h21081408ff07e207c907cb07da07ec0704080708ef07d007a80783077a077e07;
    inBuf[7805] = 256'h8407920791078007790772076d077707760764075107370722072f0755078f07;
    inBuf[7806] = 256'he30733087108a308b408a60890086f084e084908500860087d088a087f086708;
    inBuf[7807] = 256'h3708f507bb078307540744074307500776079c07ba07dd07f307ff0718082e08;
    inBuf[7808] = 256'h40085c086e0877088d08a408bc08e108f408ea08cd08910845080d08e307cc07;
    inBuf[7809] = 256'hd107d607d107cc07ba07a1079a0798079b07b207c807dc07fc07180830085608;
    inBuf[7810] = 256'h77089108ad08b3089e087e084a081208f207e107de07ec07ec07d507b4078207;
    inBuf[7811] = 256'h4b072b07170710072107380755078607b707e8071d08410852085c0850083308;
    inBuf[7812] = 256'h1408e807b6078f07650737070d07d606970666064106370653068106b406eb06;
    inBuf[7813] = 256'h100725073b0748074f075d0760075b075a074e0737071c07ee06b3067e064e06;
    inBuf[7814] = 256'h2e062806270623061d060906ef05e005d405cc05ce05c805b905ad059c058d05;
    inBuf[7815] = 256'h8c058a0589058e058c0585058405820585059905b105cc05e805f005e205c205;
    inBuf[7816] = 256'h8c0549050905c604860450041c04f003d203b803a4039603840373036f037603;
    inBuf[7817] = 256'h8f03bb03ea03180441045b046c04780478046b044e041804d00382033203ef02;
    inBuf[7818] = 256'hbe02960276025a02390219020102f101ee01fb010f022a0247025b0266026402;
    inBuf[7819] = 256'h4f022d020302d301a90189016f015b0148012e011301f700db00c700ba00af00;
    inBuf[7820] = 256'ha700a1009a009a00a100ad00be00c500b80091004e00f7ffa3ff5fff39ff37ff;
    inBuf[7821] = 256'h4bff62ff6dff5cff30fff5feb8fe86fe6bfe61fe68fe7efe99feb5fecffeddfe;
    inBuf[7822] = 256'hdcfed0feb4fe8ffe6afe3efe10fee7fdbefd9dfd8efd83fd78fd63fd32fdebfc;
    inBuf[7823] = 256'ha1fc5dfc38fc3efc5ffc8ffcbffcd6fcd3fcbbfc8cfc57fc2efc0cfcfdfb03fc;
    inBuf[7824] = 256'h0afc11fc14fc01fce0fbbcfb8dfb5efb37fb0bfbe6fad3fac7facefae5faf6fa;
    inBuf[7825] = 256'hfdfaf9fadafaaefa83fa54fa31fa23fa1bfa1dfa25fa1cfa05fae8f9b9f98af9;
    inBuf[7826] = 256'h69f947f92df91ef909f9fbf802f911f932f961f980f98cf984f958f920f9f0f8;
    inBuf[7827] = 256'hc0f8a6f8a5f8a1f89ff899f875f841f809f8c6f78ff773f760f762f777f784f7;
    inBuf[7828] = 256'h96f7b1f7c1f7d5f7eef7f3f7ebf7d8f7a5f769f734f7fef6e2f6e7f6f5f610f7;
    inBuf[7829] = 256'h2ff733f727f716f7f3f6d8f6cff6c5f6c5f6cef6c2f6b3f6a5f685f668f657f6;
    inBuf[7830] = 256'h3cf628f61ff60bf6fcf5f4f5def5d2f5d8f5ddf5f2f513f61ff61ff616f6f5f5;
    inBuf[7831] = 256'hdbf5d7f5daf5f4f520f63af64af652f639f618f6f7f5c3f592f56af539f515f5;
    inBuf[7832] = 256'h09f5fef409f52af543f560f577f56af550f539f51cf51cf542f571f5abf5e2f5;
    inBuf[7833] = 256'hf4f5f3f5e6f5bef596f574f541f515f5faf4e4f4edf416f53cf568f58ff590f5;
    inBuf[7834] = 256'h82f56df546f52af523f520f536f565f58bf5b0f5c9f5b9f596f56df537f518f5;
    inBuf[7835] = 256'h1af525f547f577f596f5b3f5cef5d2f5d5f5dcf5d1f5cdf5d4f5d6f5e9f50cf6;
    inBuf[7836] = 256'h26f643f65af651f63bf61ef6eef5caf5b9f5abf5b6f5d5f5ebf506f622f62cf6;
    inBuf[7837] = 256'h37f64af656f66ef693f6b1f6d9f60af72df752f772f773f765f74ff725f707f7;
    inBuf[7838] = 256'hfbf6f3f600f71cf731f74ef76ff77df786f788f774f767f76cf77cf7a9f7e9f7;
    inBuf[7839] = 256'h1bf843f85bf857f853f85af860f876f896f8acf8c8f8e8f8fdf815f92af92bf9;
    inBuf[7840] = 256'h27f920f90ff90cf918f928f949f973f995f9b7f9d1f9d5f9d0f9c9f9c0f9cef9;
    inBuf[7841] = 256'hf8f92ffa74fab3fad7fae9faecfadefad6fad7fad8fae1faeffafafa15fb3dfb;
    inBuf[7842] = 256'h6afba1fbd5fbf5fb08fc0bfcfefbf1fbe9fbe9fbfffb27fc53fc81fca4fcb0fc;
    inBuf[7843] = 256'hb2fcb2fcb5fccdfcf7fc27fd5bfd88fda4fdbafdc8fdd0fdd9fde0fde5fdf0fd;
    inBuf[7844] = 256'hfdfd0bfe20fe35fe46fe5dfe78fe94feb3fecbfedbfeedfe02ff22ff54ff8eff;
    inBuf[7845] = 256'hc8fffaff140016000a00f6ffe9ffe9fff3ff0900280044005800660069006800;
    inBuf[7846] = 256'h6a0074008f00be00f60037017801ae01dd0102021902280230022d0229022602;
    inBuf[7847] = 256'h1f022102270229022c022b02250224022b0239025b028f02ca0212035b039603;
    inBuf[7848] = 256'hc703e703ef03f003eb03e003e003e603ec03f9030504090414041b0417041a04;
    inBuf[7849] = 256'h1e041f04300450047704b304f304260554056f056f056c056205530556056305;
    inBuf[7850] = 256'h73059205ad05ba05c605c505b305ab05a505a005b305d205f305250658068106;
    inBuf[7851] = 256'hae06d006e206f406fa06ee06e806df06cf06d606e406f1060907180713071207;
    inBuf[7852] = 256'h0907fc0607071d07340760078907a107bf07d407db07ed07f707f50700080508;
    inBuf[7853] = 256'h01081208260832084b085808530853084a0839083d084308420852085b085708;
    inBuf[7854] = 256'h63086c086f0887089e08ac08cb08e408f0080c09200928093d09490943094609;
    inBuf[7855] = 256'h3e092809220918090909100912090a0915091a091709270936093d0959097009;
    inBuf[7856] = 256'h7c099609a709aa09bb09c109b809bb09b4099e099909910985099509a509ab09;
    inBuf[7857] = 256'hbc09bd09ac09a909a1099609a809b909c109dd09f309fc09120a1a0a100a0f0a;
    inBuf[7858] = 256'hfd09dd09d209c509b709c609d509da09f009f909ef09ef09e109c909c809c609;
    inBuf[7859] = 256'hc209d609e509ed09080a190a190a230a1b0aff09ed09d309b509b409b709b909;
    inBuf[7860] = 256'hd109e309e709f809fa09ed09ed09df09c709c409be09b309b909b3099f099809;
    inBuf[7861] = 256'h84096909660960095509600968096c0986099a09a409b809bb09ac09a7099409;
    inBuf[7862] = 256'h78096a0950092c091d090d09fe0808090e0909090b09fb08dd08ce08bc08ad08;
    inBuf[7863] = 256'hb808c208c708d908e008d908dc08cf08b608a9089208730864084f0839083908;
    inBuf[7864] = 256'h3b083e0853085a0852084a082f080508e907cc07b407b207ae07aa07b407b407;
    inBuf[7865] = 256'ha907a70797077a0765074b07310728071d0712071607120709070a070007ec06;
    inBuf[7866] = 256'hdc06c106a20690067e0672067a067e067b067b066e065706450629060806ee05;
    inBuf[7867] = 256'hce05b305aa05a1059a059d0593057e056b054e0530051d050705f104e504d704;
    inBuf[7868] = 256'hce04d104cf04cb04ca04be04ab049a047f0464044e0434041d0411040504fa03;
    inBuf[7869] = 256'hf103db03bb03960368033b031a03fd02ea02e402e202e602f002f302f302ea02;
    inBuf[7870] = 256'hce02ab0288026402470237022c0224021a020b02fc01e901cd01af0193017401;
    inBuf[7871] = 256'h5b01470136012a011e010d01ff00f000db00c600ae008f007000520035002200;
    inBuf[7872] = 256'h13000400faffeaffd7ffc7ffb3ff9cff89ff72ff57ff41ff2cff1bff13ff09ff;
    inBuf[7873] = 256'hfdfef5fee6fed3fec3feaffe98fe81fe60fe40fe27fe07fee6fdd1fdb8fd9ffd;
    inBuf[7874] = 256'h8dfd79fd65fd56fd41fd2efd25fd17fd0ffd0ffd06fdf8fce9fccdfcaefc96fc;
    inBuf[7875] = 256'h79fc60fc50fc39fc25fc1bfc0bfcfdfbf6fbe2fbcbfbb7fb97fb7bfb6cfb59fb;
    inBuf[7876] = 256'h48fb3cfb21fb05fbf0fad3fabafaadfa98fa88fa83fa75fa6cfa6dfa64fa5cfa;
    inBuf[7877] = 256'h58fa48fa3cfa36fa21fa0bfaf9f9d7f9b5f99ef97cf95ff94ff93af92df92cf9;
    inBuf[7878] = 256'h1ff914f90ff9f7f8dff8cff8b5f8a5f8a4f89cf89bf8a2f896f88af885f86df8;
    inBuf[7879] = 256'h53f841f822f808f8f9f7e2f7d4f7d3f7c4f7bbf7bcf7aaf79af793f77ff772f7;
    inBuf[7880] = 256'h73f768f763f767f757f747f73df721f70af703f7f2f6ebf6edf6ddf6cef6c6f6;
    inBuf[7881] = 256'haaf693f68af676f66ff675f66ef670f67ef67af67cf686f67af66df667f651f6;
    inBuf[7882] = 256'h42f63ff62ef626f62bf61ef616f615f6fdf5e8f5dbf5bbf5a7f5a6f59ef5a4f5;
    inBuf[7883] = 256'hbaf5bff5c8f5d4f5c9f5c1f5c2f5b2f5abf5b2f5abf5aef5b9f5b2f5aff5b4f5;
    inBuf[7884] = 256'ha4f59cf59ef590f588f588f577f56ff575f570f578f58bf58af586f582f56af5;
    inBuf[7885] = 256'h5df562f55ef568f57df582f58ff5a4f5a5f5adf5bef5b9f5b5f5b7f5aaf5a5f5;
    inBuf[7886] = 256'haaf5a2f5a4f5aff5aaf5aff5bcf5b2f5acf5aef5a2f5a3f5b3f5baf5cef5e7f5;
    inBuf[7887] = 256'hedf5fbf511f617f623f634f631f631f636f62df631f641f644f64df65af654f6;
    inBuf[7888] = 256'h57f664f665f66ff680f682f68cf69df6a1f6adf6c4f6cff6e2f6fbf607f71af7;
    inBuf[7889] = 256'h2ef72ff732f73bf737f73bf748f74cf75af76ff776f784f798f79df7a9f7b8f7;
    inBuf[7890] = 256'hbaf7c5f7d8f7e6f702f827f83ff85af872f877f87ef889f889f893f8a6f8aff8;
    inBuf[7891] = 256'hbff8d8f8e9f8fdf811f918f924f92ff92df935f944f94cf95df977f98df9abf9;
    inBuf[7892] = 256'hcef9e5f9fbf90bfa0efa1afa2efa3efa5bfa80fa9dfabbfad7fae6faf6fa00fb;
    inBuf[7893] = 256'hfcfafafaf7faedfaf1fa02fb15fb34fb5afb7afb9cfbbdfbd4fbecfbfefb08fc;
    inBuf[7894] = 256'h17fc2bfc3dfc5bfc7cfc95fcabfcbafcbcfcc0fcc4fcc7fcd4fce7fcfafc19fd;
    inBuf[7895] = 256'h3cfd5bfd7afd96fda8fdb6fdc0fdc9fddefdf5fd09fe21fe36fe44fe54fe63fe;
    inBuf[7896] = 256'h6ffe7efe8bfe97fea8febdfed3fef0fe0dff29ff44ff59ff6aff7fff90ff9dff;
    inBuf[7897] = 256'hadffbfffd5fff1ff0a001e00300039003c0042004a00560067007a009000a900;
    inBuf[7898] = 256'hbf00d700f100040116012a013d014f016201730185019601a201b201c701d901;
    inBuf[7899] = 256'hec01fd010802170226023102400250025c026b0279027f028b029d02ac02be02;
    inBuf[7900] = 256'hcf02dc02ee0201031103250338034403540364036e037d038d039903ab03bc03;
    inBuf[7901] = 256'hc403ce03d703d903e203ed03f203fd030904130426043704430458046d047a04;
    inBuf[7902] = 256'h8b049a04a104ad04b904bd04c804d004d004d904e204e304eb04f304fa040a05;
    inBuf[7903] = 256'h17051e052f053e05440553056205670574057f0582058e0599059c05a705af05;
    inBuf[7904] = 256'haf05b605ba05ba05c705d705df05f005fc05fd05080610060f0619061f061e06;
    inBuf[7905] = 256'h2806310636064706530654065a065a0653065b06620664067006780678068606;
    inBuf[7906] = 256'h91069506a206a806a306aa06af06ad06b506bb06ba06c206c906cb06db06e506;
    inBuf[7907] = 256'he406ea06e706d706d906de06de06eb06f606fa060407070700070307ff06f306;
    inBuf[7908] = 256'hf606fa06fb060a071607190726072c0729073107320728072807220716071c07;
    inBuf[7909] = 256'h2507280735073b07340735072d071e071b07150707070a070e07110725073307;
    inBuf[7910] = 256'h34073d073d072f072a0725071f07230720071507180718071007150716070d07;
    inBuf[7911] = 256'h0d070707ff0607070b07080710071007040703070107f906f706ee06e106e106;
    inBuf[7912] = 256'hdf06d706dd06de06d606d906d606cc06d006cf06c406c206bc06b106b406b506;
    inBuf[7913] = 256'hb106b306a80694068d06840678067c067f067b067e067d0677067c0679066f06;
    inBuf[7914] = 256'h6f066706560652064f06460645064106360633062d06240623061606ff05f305;
    inBuf[7915] = 256'he605d905df05e505e505ec05ed05e605e305dd05d205cf05c505b705b705b605;
    inBuf[7916] = 256'hb105b305ad059c058b0574055c055005410530052a052505200526052d052f05;
    inBuf[7917] = 256'h3405300523051e0517050f050d050705fc04f804ef04df04d204bb049c048304;
    inBuf[7918] = 256'h6b045a045b045d045c04600460045f04630463045f04590447042f0421041604;
    inBuf[7919] = 256'h0d040f040c04ff03f003d903be03aa03980386037a036f0367036a036c036a03;
    inBuf[7920] = 256'h6903610355034f03490344034503400335032b031d030f030703fc02eb02d802;
    inBuf[7921] = 256'hc102aa029b028d02810278026a025c0254024d02480248024802460247024502;
    inBuf[7922] = 256'h42023e02340229021e020f02fd01f001e401d701c501af019c01900182017601;
    inBuf[7923] = 256'h6f0167015c01550150014e014c01480143013b01310127011e0113010901ff00;
    inBuf[7924] = 256'hf200e800e300dd00d600ca00b800a4008f007e0072006a0062005c0059005800;
    inBuf[7925] = 256'h5800560052004c0042003200230016000c0007000200fbfff4ffebffdfffd1ff;
    inBuf[7926] = 256'hc0ffadff9aff86ff74ff6aff65ff66ff6fff74ff73ff73ff6eff62ff55ff45ff;
    inBuf[7927] = 256'h36ff28ff1cff17ff17ff15ff11ff0cff00ffeefeddfeccfebefeb7feb1feaefe;
    inBuf[7928] = 256'haefeabfea5fe9ffe93fe83fe75fe66fe5cfe58fe54fe52fe53fe4ffe4bfe4bfe;
    inBuf[7929] = 256'h4afe46fe43fe37fe2afe20fe15fe0cfe0afe04fefafdeffdddfdcafdbbfdaefd;
    inBuf[7930] = 256'ha6fda4fd9ffd9ffda6fda8fdaafdaefdaafda3fd9dfd92fd89fd87fd83fd7efd;
    inBuf[7931] = 256'h79fd71fd6afd65fd5afd50fd49fd39fd29fd23fd1cfd1bfd21fd24fd23fd21fd;
    inBuf[7932] = 256'h16fd0efd0bfd04fdfefcfdfcf9fcf6fcfbfcfcfcfdfcfdfcf3fce7fcddfccdfc;
    inBuf[7933] = 256'hc0fcb9fcadfca6fca7fca3fca1fca5fca3fca0fc9ffc98fc94fc96fc97fc9efc;
    inBuf[7934] = 256'ha9fcabfcadfcb2fcadfca4fc9afc86fc6ffc5efc4efc46fc48fc47fc48fc4cfc;
    inBuf[7935] = 256'h47fc44fc49fc4cfc54fc5dfc5dfc5efc64fc66fc6dfc78fc78fc6ffc67fc58fc;
    inBuf[7936] = 256'h49fc3efc2efc21fc19fc0efc0afc12fc18fc22fc2dfc2cfc2bfc2ffc30fc36fc;
    inBuf[7937] = 256'h3ffc3ffc3cfc3bfc37fc3afc43fc44fc42fc3efc2ffc1ffc17fc0ffc0cfc0cfc;
    inBuf[7938] = 256'h06fc07fc0ffc15fc1ffc2cfc2dfc28fc27fc22fc23fc29fc2bfc2dfc2ffc2efc;
    inBuf[7939] = 256'h31fc39fc39fc3afc38fc2afc1bfc13fc0bfc0dfc17fc1afc21fc2cfc34fc3bfc;
    inBuf[7940] = 256'h43fc40fc38fc2ffc22fc1cfc22fc29fc36fc43fc46fc4afc53fc55fc56fc54fc;
    inBuf[7941] = 256'h45fc36fc2bfc23fc2bfc41fc54fc65fc71fc70fc6afc62fc51fc40fc32fc26fc;
    inBuf[7942] = 256'h2afc3cfc4ffc67fc80fc87fc85fc81fc76fc6efc6bfc64fc60fc63fc6afc7afc;
    inBuf[7943] = 256'h8efc99fca1fca3fc94fc81fc77fc72fc74fc7dfc82fc8bfc98fc9ffca9fcb3fc;
    inBuf[7944] = 256'haffca7fca1fc98fc94fc99fca2fcb3fcc5fccffcdbfce9fce9fce3fcdafcc6fc;
    inBuf[7945] = 256'hb3fca8fca3fcabfcbdfccbfcd8fce4fce8fcebfceffcebfce9fce8fce5fcecfc;
    inBuf[7946] = 256'hfdfc0dfd20fd30fd2ffd24fd17fd06fdfafcf2fce7fce3fceafcf2fc02fd18fd;
    inBuf[7947] = 256'h2bfd38fd3cfd34fd2efd30fd30fd35fd3dfd41fd46fd4dfd4dfd4dfd4cfd43fd;
    inBuf[7948] = 256'h39fd32fd2efd32fd3afd40fd48fd52fd54fd5afd63fd67fd68fd6afd66fd64fd;
    inBuf[7949] = 256'h67fd6afd75fd82fd86fd85fd85fd80fd7ffd80fd7efd7dfd7efd7afd7afd7efd;
    inBuf[7950] = 256'h80fd87fd8ffd90fd93fd9afda2fdabfdb6fdbbfdc0fdc7fdcbfdd0fdd5fdd2fd;
    inBuf[7951] = 256'hccfdc3fdb5fdaefdb0fdb5fdbffdcbfdd0fdd2fdd7fddafdddfde3fde8fdeefd;
    inBuf[7952] = 256'hf5fdfbfd06fe12fe19fe1afe19fe13fe10fe10fe10fe15fe1efe22fe25fe2afe;
    inBuf[7953] = 256'h2ffe35fe3cfe3ffe40fe41fe41fe45fe4bfe4ffe54fe5afe5efe62fe65fe67fe;
    inBuf[7954] = 256'h6dfe75fe7bfe82fe8dfe97fe9ffea4fea5fea2fe9dfe99fe9bfea4feaefeb7fe;
    inBuf[7955] = 256'hbefec2fec5fecafecdfed1fed4fed4fed5fedefee8fef4fefffe07ff09ff09ff;
    inBuf[7956] = 256'h06ff06ff0cff12ff17ff1dff26ff36ff47ff51ff55ff51ff45ff37ff32ff35ff;
    inBuf[7957] = 256'h3eff4eff5fff6fff7dff88ff92ff97ff95ff8fff88ff83ff86ff93ffa6ffbcff;
    inBuf[7958] = 256'hceffd9ffdfffe2ffdeffd3ffc5ffb8ffafffb0ffbbffd1fff1ff0e0021002700;
    inBuf[7959] = 256'h26001e0015000f000e0014001d002e00480062007700840087007d006c005e00;
    inBuf[7960] = 256'h5500500052005c006d0081009400a700b800bd00b500a600970093009e00b200;
    inBuf[7961] = 256'hcd00ea0002011501210123011b010e01fc00eb00e200e200ed00000116012a01;
    inBuf[7962] = 256'h3a0145014a014c0147013f013901380142015b0179019501ac01b701b501ab01;
    inBuf[7963] = 256'h9901860177016c0168016f0180019901b501cd01de01e601e201da01d601d301;
    inBuf[7964] = 256'hd301db01e501f00101021402250231023102270218020502f801f901fe010602;
    inBuf[7965] = 256'h1502250236024a025a026402690260025202490246024a025602650273028302;
    inBuf[7966] = 256'h8e0295029d029d02940288027a027202760281028e029f02ad02b602c102c802;
    inBuf[7967] = 256'hca02cb02c602ba02b202af02b502c502d602e502f202f402f102ef02e802df02;
    inBuf[7968] = 256'hdd02dd02df02e902f80208031a03240328032a0325031d03180312030a030903;
    inBuf[7969] = 256'h09030c031a03290334033e033e03370332032c0327032b0333033b0348035603;
    inBuf[7970] = 256'h62036e036f03640359034a033d033b033e0344034f0357035d036a0373037503;
    inBuf[7971] = 256'h75036f0362035a0358035c03690374037a03810382037d037c0378036f036e03;
    inBuf[7972] = 256'h6d036c03710376037a03810383037e037d037b037703770374036e0370037303;
    inBuf[7973] = 256'h76038303910398039f039f039803910389038103820384038303870388038303;
    inBuf[7974] = 256'h81037a036e036603620363036e037a03840393039c039e03a303a20398038f03;
    inBuf[7975] = 256'h840377037103700372037d038603870386037e0371036b0365035f0362036a03;
    inBuf[7976] = 256'h720383039403990398038f037f03740368035f036203670369036f0373037203;
    inBuf[7977] = 256'h730371036703600356034b034b034d034e035803610366036d0370036c036903;
    inBuf[7978] = 256'h63035803500347033d033e033f033d03420345033f033a0335032b0325031f03;
    inBuf[7979] = 256'h160318031f03260333033c0340034503430337032b031c030903fd02f402ee02;
    inBuf[7980] = 256'hf502000306030c030c030303fd02f602ec02e702e302dd02e102e602e802ee02;
    inBuf[7981] = 256'hee02e402dd02d402c402b902b102a802a602a802aa02b302be02c202c502bf02;
    inBuf[7982] = 256'had029f02930284027e027b0278027d02820285028c028c028102760267025202;
    inBuf[7983] = 256'h4202390235023a02450250025b025f025c0259024c02350226021b0211021202;
    inBuf[7984] = 256'h18021e0225022802210218020802f101de01cb01b801b201b601bf01d201e301;
    inBuf[7985] = 256'hec01ef01e701d501c301b0019d0194019101910198019f019d0197018a017701;
    inBuf[7986] = 256'h660155014301380130012c0132013c014701540159015001430132011b010801;
    inBuf[7987] = 256'hfa00f200f100f300f500fa00fa00f200ea00da00c300ae009b008b0081007d00;
    inBuf[7988] = 256'h80008a009400970096008e0080006f005f005000470043004200440045004100;
    inBuf[7989] = 256'h3c00310020000e00fcffe9ffdaffd0ffcaffc7ffc8ffcdffd3ffd6ffd5ffd0ff;
    inBuf[7990] = 256'hc5ffb6ffa9ff9eff94ff8cff87ff83ff7dff74ff68ff5dff50ff43ff38ff30ff;
    inBuf[7991] = 256'h2bff25ff21ff1fff1eff1dff1dff1dff1aff14ff0afffcfeedfedffed1fec6fe;
    inBuf[7992] = 256'hbdfeb9feb7feb4feb1feaefea5fe98fe8cfe7ffe73fe6bfe69fe6bfe6efe6dfe;
    inBuf[7993] = 256'h68fe62fe59fe4ffe48fe3dfe32fe29fe21fe1afe16fe11fe0cfe08fefdfdf1fd;
    inBuf[7994] = 256'heafde2fdd7fdcdfdc3fdbcfdb8fdb5fdb5fdb8fdb6fdb1fdabfda0fd96fd8ffd;
    inBuf[7995] = 256'h86fd7ffd79fd70fd68fd65fd5efd55fd4efd46fd3ffd37fd2afd21fd1ffd1cfd;
    inBuf[7996] = 256'h1dfd23fd24fd24fd22fd17fd0bfdfffceefce0fcd8fccffccbfccdfccbfcc9fc;
    inBuf[7997] = 256'hcbfcc7fcc3fcbffcb8fcb6fcb7fcb1fcacfcacfca6fca2fca0fc96fc89fc80fc;
    inBuf[7998] = 256'h73fc68fc61fc57fc54fc59fc5bfc60fc68fc66fc62fc5dfc52fc4cfc4efc4cfc;
    inBuf[7999] = 256'h4ffc55fc51fc4dfc4cfc42fc37fc30fc23fc18fc13fc0dfc0ffc18fc18fc1afc;
    inBuf[8000] = 256'h20fc20fc20fc21fc17fc11fc0ffc06fc02fc07fc0afc10fc18fc17fc14fc11fc;
    inBuf[8001] = 256'h03fcf9fbf3fbe9fbe5fbeafbebfbf1fbfcfbfffb02fc06fcfffbfafbfafbf2fb;
    inBuf[8002] = 256'heffbf5fbf5fbfafb00fcfffbfdfbfcfbf1fbe8fbe3fbd8fbd8fbe0fbe0fbe4fb;
    inBuf[8003] = 256'hecfbeffbf4fbfcfbfbfbfbfbfcfbf4fbf0fbf1fbecfbedfbf3fbf4fbf9fb02fc;
    inBuf[8004] = 256'h03fc05fc05fcfbfbf5fbf3fbebfbedfbfafb01fc08fc0efc0dfc0ffc14fc11fc;
    inBuf[8005] = 256'h13fc17fc14fc15fc1afc19fc1cfc25fc28fc2ffc37fc36fc36fc39fc33fc2ffc;
    inBuf[8006] = 256'h30fc2ffc34fc3cfc3efc46fc51fc55fc5cfc66fc68fc6cfc71fc6ffc72fc78fc;
    inBuf[8007] = 256'h79fc7ffc89fc8cfc94fc9dfc9cfc98fc97fc91fc91fc97fc9efcadfcc0fccbfc;
    inBuf[8008] = 256'hd9fce6fce6fce7fceafce9fcecfcf2fcf3fcf8fcfffc02fd09fd14fd19fd21fd;
    inBuf[8009] = 256'h28fd28fd2cfd32fd34fd39fd43fd4bfd57fd65fd70fd7cfd85fd83fd81fd82fd;
    inBuf[8010] = 256'h81fd86fd91fd9afda5fdb1fdb9fdc4fdcefdd2fdd7fddbfdd8fdd6fdd8fdd9fd;
    inBuf[8011] = 256'he0fdeffdfefd11fe23fe2efe35fe37fe33fe32fe36fe3cfe4afe5bfe67fe71fe;
    inBuf[8012] = 256'h78fe7bfe7dfe7efe7dfe80fe87fe8cfe95fea2feaffebdfeccfed9fee4feebfe;
    inBuf[8013] = 256'heefef1fef1feeffef1fef8fe00ff09ff15ff1fff27ff2fff35ff3cff44ff4cff;
    inBuf[8014] = 256'h56ff5fff67ff6fff78ff81ff8cff98ffa2ffa7ffa9ffa9ffa9ffabffb1ffbaff;
    inBuf[8015] = 256'hc6ffd5ffe4fff3ffffff08000e001100130016001c0022002900300037003c00;
    inBuf[8016] = 256'h43004b0053005a0062006b007300790080008b0093009b00a500ae00b500bb00;
    inBuf[8017] = 256'hc000c200c500cb00d400e100eb00f400fc00fe00ff00020106010b0114011c01;
    inBuf[8018] = 256'h24012c012f01310138013e0145014f0156015b0165016c01720178017c018001;
    inBuf[8019] = 256'h87018b018e019401970198019e01a201a801b301bb01c001c501c601c801d101;
    inBuf[8020] = 256'hda01e501f201f701f801fc01fc01fc010102030206020d021002120216021902;
    inBuf[8021] = 256'h1b022302290230023d0246024b0250025002510258025d0263026d0272027302;
    inBuf[8022] = 256'h7802780276027902780278027e02820285028b028c028b02910294029802a202;
    inBuf[8023] = 256'ha802ad02b602bb02bf02c802cd02d202da02db02d802da02da02da02de02df02;
    inBuf[8024] = 256'hdf02e302e102df02e302e402e602ed02ee02ee02f502fb0201030d0314031603;
    inBuf[8025] = 256'h1b031d031d0322032303210322031e0319031b031a0317031c031e031f032703;
    inBuf[8026] = 256'h2c03310338033b033a033d033c033b033e033d0338033b033d033f0348034b03;
    inBuf[8027] = 256'h4b034c03460340034203410341034603490349034d03500352035b035f035e03;
    inBuf[8028] = 256'h5e03590350034c034603420347034d03540360036503640364035f0356035403;
    inBuf[8029] = 256'h530352035603570355035903590358035c035c03590358035603540359035c03;
    inBuf[8030] = 256'h5d03620362035e035e035c0359035a03560350034f034e034d03500352035003;
    inBuf[8031] = 256'h510351034f0352035303510352034f03480345033f03360331032f032d033203;
    inBuf[8032] = 256'h37033a033e033d033603340331032d032e032d032803260323031e031c031a03;
    inBuf[8033] = 256'h150312030c030103fb02f802f602fb020003020305030303fc02f802f302ec02;
    inBuf[8034] = 256'he802e202d902d402d002ca02c702c402be02bb02b802b302b302b002a802a202;
    inBuf[8035] = 256'h9e029a029c029f029e029c02940286027b027202690266026502630262026202;
    inBuf[8036] = 256'h5d025902520245023a022f0223021e021c021a021b021d021b021a0218021102;
    inBuf[8037] = 256'h0a020202f601ed01e601dd01d701d201cb01c401be01b401ab01a3019a019501;
    inBuf[8038] = 256'h92018d018901870182017e017b0174016e0168015e01530148013a012f012701;
    inBuf[8039] = 256'h1e01180112010b0105010001fa00f400ef00e900e200dd00d600d100cf00ca00;
    inBuf[8040] = 256'hc100b700a9009b00900086007f007a0072006a0063005a0052004e0049004400;
    inBuf[8041] = 256'h3f0037002b00200015000e000d000c000b0007000000f5ffe9ffddffd1ffc8ff;
    inBuf[8042] = 256'hbdffb2ffa9ffa0ff98ff91ff89ff7fff77ff6fff68ff63ff5eff57ff53ff50ff;
    inBuf[8043] = 256'h4eff4dff4bff44ff38ff28ff16ff07fffafeedfee3fedafed0fec8fec4fec2fe;
    inBuf[8044] = 256'hc4fec7fec6fec3febefeb4feaafea0fe94fe8afe82fe77fe6efe66fe5bfe52fe;
    inBuf[8045] = 256'h4bfe43fe3cfe37fe30fe2cfe2afe26fe23fe21fe1afe12fe0afefefdf4fdebfd;
    inBuf[8046] = 256'he1fddafdd6fdcffdcbfdc9fdc4fdbffdbbfdb4fdaefdabfda4fd9dfd98fd90fd;
    inBuf[8047] = 256'h89fd85fd7dfd75fd6ffd64fd5dfd5bfd58fd58fd5dfd5cfd59fd58fd51fd4bfd;
    inBuf[8048] = 256'h48fd41fd3bfd36fd2afd1efd16fd0cfd05fd04fd01fd00fd03fd01fd02fd06fd;
    inBuf[8049] = 256'h06fd06fd08fd05fd01fd00fdf9fceffce6fcd6fcc7fcc1fcbcfcbdfcc5fcc9fc;
    inBuf[8050] = 256'hccfcd0fccffccefcd3fcd3fcd4fcd6fcd1fccafcc6fcbcfcb3fcaffca7fca2fc;
    inBuf[8051] = 256'ha2fc9dfc9bfc9efc9ffca4fcaffcb4fcb7fcbbfcb5fcaefcacfca5fca1fca3fc;
    inBuf[8052] = 256'h9ffc9dfca0fc9dfc9bfc9dfc99fc97fc9afc9bfca0fcaafcaefcb2fcb8fcb7fc;
    inBuf[8053] = 256'hb5fcb6fcb0fca8fca4fc9afc94fc95fc94fc97fca3fcaafcb4fcc1fcc6fccafc;
    inBuf[8054] = 256'hd0fccefccdfcd1fccffccffcd3fcd2fcd1fcd5fcd3fcd3fcd7fcd7fcdafce5fc;
    inBuf[8055] = 256'hecfcf4fc00fd04fd07fd0efd10fd15fd1cfd1cfd19fd18fd12fd0ffd16fd1efd;
    inBuf[8056] = 256'h29fd39fd42fd4afd52fd55fd58fd60fd62fd64fd69fd68fd68fd6ffd75fd7efd;
    inBuf[8057] = 256'h8cfd91fd95fd9afd9afd9cfda5fdaafdaffdb7fdbafdbffdc9fdd1fddbfde9fd;
    inBuf[8058] = 256'hf1fdf9fd03fe07fe09fe0cfe08fe05fe07fe0afe12fe21fe2dfe3afe48fe50fe;
    inBuf[8059] = 256'h57fe5ffe62fe63fe66fe64fe63fe67fe69fe71fe7ffe8efe9ffeb3fec1feccfe;
    inBuf[8060] = 256'hd4fed3fed0fecdfec6fec2fec4fec6fecdfed7fedffee7fef1fefbfe09ff1cff;
    inBuf[8061] = 256'h2bff38ff41ff43ff43ff45ff44ff44ff44ff40ff3cff3cff3eff46ff55ff65ff;
    inBuf[8062] = 256'h76ff89ff97ffa2ffaaffadffadffadffadffaeffb0ffb0ffb0ffb0ffb0ffb5ff;
    inBuf[8063] = 256'hbeffc9ffd5ffe1ffebfff4ffffff0b00170022002b0032003600390039003700;
    inBuf[8064] = 256'h33002c00260021001f001e002100290036004a00610079008e009e00a900af00;
    inBuf[8065] = 256'hb000ae00a900a000940088007d00750076007e008d00a000b400c400d200db00;
    inBuf[8066] = 256'he000e300e200dd00d600cf00c900c700ca00cd00d400db00e200ee00fb000901;
    inBuf[8067] = 256'h170122012601270125011d0114010801f900ef00ea00ec00f9000a011c012e01;
    inBuf[8068] = 256'h3c014401480146013c01320126011b0119011d012601350143014c0150014c01;
    inBuf[8069] = 256'h40013401280120012201280131013e014b01560163016d0170016f0167015701;
    inBuf[8070] = 256'h48013c0131012e012c012b01300136013f014d015c01680174017c017d017d01;
    inBuf[8071] = 256'h750165015501430130012601220121012b013b0150016a018201900196018f01;
    inBuf[8072] = 256'h7b01660150013c0132012c0129012e01370140014e015b0164016e0175017801;
    inBuf[8073] = 256'h7b017b0174016c0160014e013f012e011d0115011301170127013c014f016201;
    inBuf[8074] = 256'h6f017401790179017601760173016a01620158014b0144013b012e0122011201;
    inBuf[8075] = 256'h0001f500f100f60008011f013901590176018e01a201aa01a2018f0170014901;
    inBuf[8076] = 256'h25010201e000c800b600ad00b600cc00eb0014013b015d017d0192019a019801;
    inBuf[8077] = 256'h8501610136010701dd00c200b500b400c300d800f0000c012501370145014901;
    inBuf[8078] = 256'h41013601270116010e010a010701090109010601070109010e0116011c011a01;
    inBuf[8079] = 256'h1701100108010301ff00f600ef00e700e200ea00fa000e012301300132012f01;
    inBuf[8080] = 256'h260117010701f300dd00d100d400e7000b01330150015c01530137011101e600;
    inBuf[8081] = 256'hbb009a00850082009800c200f9003401640180018a018101670144011c01f000;
    inBuf[8082] = 256'hcc00b200a600ac00bf00d800f4000b011a0125012b012c012c012a0124011f01;
    inBuf[8083] = 256'h1a0113010e010a010301000100010501140129013f0153015e015c014f013801;
    inBuf[8084] = 256'h1801f800d800bd00ae00ae00bd00dd0005012d0152016c0179017f017d017401;
    inBuf[8085] = 256'h69015d014f014101330120010c01f700e000d000c800c800d300e500f9001301;
    inBuf[8086] = 256'h30014c016b0187019b01aa01b301b401b101a7019101700143010b01d400a700;
    inBuf[8087] = 256'h87007e008b00aa00dc001b016101a901e90115022c0228020b02df01a8016901;
    inBuf[8088] = 256'h2d01f500c600ab00a800ba00e000100142017401a301cc01ed01fd01f301d101;
    inBuf[8089] = 256'h9c015e012b010b01ff000a012301450170019d01c101d901da01c1019b017001;
    inBuf[8090] = 256'h4a0135012c012b0136014801610181019e01ae01b201a80197018f018f019401;
    inBuf[8091] = 256'h9b0199018c017d01710169016a016c016a0168016501620167016a0167016101;
    inBuf[8092] = 256'h55014a014d015f017b01a201c701e101f201f301df01ba0182013a01f400bd00;
    inBuf[8093] = 256'ha000ac00d9001c016b01b201e70108020e02f701cb0189013e010001d800cd00;
    inBuf[8094] = 256'he1000501290148015c01660171017a017d017e0178016e016a0166015a014301;
    inBuf[8095] = 256'h1701dd00a9008a008b00b300f20038017d01b301d601e601d701a4015601f400;
    inBuf[8096] = 256'h940054003b0049007700af00e2000e01290131012b010f01e500c000aa00b300;
    inBuf[8097] = 256'he40029016e01a201af0193015601fc0090002000b3ff5aff2bff2fff68ffd3ff;
    inBuf[8098] = 256'h5300d20042019401c401d801c90197014e01ee0087002b00d9ff96ff65ff42ff;
    inBuf[8099] = 256'h33ff45ff74ffbeff19006c00ac00d800ec00ef00e700ca009a005e001700d5ff;
    inBuf[8100] = 256'ha8ff8aff7aff75ff71ff72ff81ff99ffb9ffdefff6ff00000300fcfff1ffe7ff;
    inBuf[8101] = 256'hd4ffbaffa0ff83ff6fff69ff69ff6aff6bff62ff56ff4dff46ff44ff4aff4fff;
    inBuf[8102] = 256'h58ff68ff77ff84ff8bff7dff59ff26ffe6feadfe87fe76fe7efe9cfec7fefefe;
    inBuf[8103] = 256'h3cff73ff9affa5ff86ff45ffeffe96fe51fe2dfe25fe36fe55fe74fe90fea7fe;
    inBuf[8104] = 256'hb1feaefea0fe88fe74fe6ffe77fe89fe9afe9cfe8efe77fe5bfe44fe35fe25fe;
    inBuf[8105] = 256'h16fe0afe04fe0efe27fe41fe55fe57fe41fe1efef5fdc8fd9cfd71fd4afd32fd;
    inBuf[8106] = 256'h36fd59fd9ffdf9fd56feaafee9fe0aff0affe1fe88fe07fe6bfdcbfc45fcebfb;
    inBuf[8107] = 256'hc5fbd2fb07fc5bfccbfc51fde2fd71fee2fe21ff23ffe9fe81fe03fe83fd10fd;
    inBuf[8108] = 256'hbafc85fc74fc83fca3fcbffcc5fca7fc69fc24fcf1fbeefb2bfca2fc41fdf2fd;
    inBuf[8109] = 256'h96fe15ff5bff51fff2fe46fe61fd6cfc93fbf4faa3faa0fad8fa3cfbbdfb48fc;
    inBuf[8110] = 256'hd2fc51fdb4fdf5fd15fe14fefcfdd7fda1fd60fd16fdc4fc75fc32fcf9fbcefb;
    inBuf[8111] = 256'haffb99fb95fbacfbdffb30fc94fcf2fc3bfd65fd68fd52fd30fd05fddefcbcfc;
    inBuf[8112] = 256'h9cfc83fc74fc69fc64fc5ffc4ffc38fc1efc05fcfafb02fc15fc35fc5ffc89fc;
    inBuf[8113] = 256'hbafcecfc10fd23fd1cfdf2fcb3fc6ffc2bfcfafbe2fbdefbf7fb2dfc75fccbfc;
    inBuf[8114] = 256'h19fd3ffd35fdf5fc86fc0bfca1fb57fb45fb6dfbc3fb42fcd3fc54fdb2fdd5fd;
    inBuf[8115] = 256'hb0fd55fdddfc5dfcf8fbb8fb9bfba4fbcbfb01fc47fc8efcc3fce5fceefcdafc;
    inBuf[8116] = 256'hc0fca9fc96fc95fca0fcadfcc0fcd3fcd8fcd3fcbdfc8cfc53fc1efcfafb02fc;
    inBuf[8117] = 256'h3afc93fc02fd69fda8fdb8fd94fd39fdc2fc42fccafb7bfb67fb90fbfcfb9afc;
    inBuf[8118] = 256'h43fde5fd5dfe94fe8efe4efedcfd53fdc5fc3cfcd3fb93fb7efb9efbecfb54fc;
    inBuf[8119] = 256'hd4fc56fdc1fd0efe2dfe12feccfd68fdf9fca5fc80fc91fce0fc59fddbfd54fe;
    inBuf[8120] = 256'ha3feaefe74fef4fd36fd61fc98fbfffac4faf9fa96fb91fcbffde9fee8ff9100;
    inBuf[8121] = 256'hc3007e00c9ffb9fe84fd5afc69fbe0facffa29fbddfbbefc9afd55fed4fe0cff;
    inBuf[8122] = 256'h10fff4fecbfeb3feb1feb9fec6febffe8efe38fec0fd33fdb4fc5bfc38fc5cfc;
    inBuf[8123] = 256'hc2fc51fdf9fd9afe16ff6cff9affa3ff9eff8fff75ff54ff24ffdafe81fe19fe;
    inBuf[8124] = 256'ha9fd45fdf7fcc4fcbbfcdafc1dfd86fd11feb4fe6eff3000e3007501ca01c401;
    inBuf[8125] = 256'h5d0195007cff3efe0bfd13fc87fb80fb00fcf6fc38fe8bffb9009001eb01c701;
    inBuf[8126] = 256'h3901650086ffd0fe61fe4cfe88fef8fe7dfff5ff43005a003300d3ff50ffc4fe;
    inBuf[8127] = 256'h4bfe06fe0afe5bfef5fec3ffa0006d0107024e023902c8010f0132005effbcfe;
    inBuf[8128] = 256'h70fe89fef9fea4ff5a00e600250104018900d8ff22ff99fe6afeaffe63ff6f00;
    inBuf[8129] = 256'ha501cb02ab031b04020464035f022101e3ffdffe3cfe12fe5bfefafec4ff8c00;
    inBuf[8130] = 256'h290185019f018501530127011a013b018a01f8016c02c902f202d6027402db01;
    inBuf[8131] = 256'h27017b00faffb8ffc2ff10008c001a019f0107024b026f027a0278026d025902;
    inBuf[8132] = 256'h3e021e02fc01e401e101f601230262029d02c402c302890218027c01cd003000;
    inBuf[8133] = 256'hcdffc2ff2600fb0028028303d004ca053c060d0640050404a1025f0181002f00;
    inBuf[8134] = 256'h65000a01eb01ca027603ce03c2036103ca0220029101410142019e014d023003;
    inBuf[8135] = 256'h230401059d05de05bd053c0575049003b002fd0196017e01ae0111027b02ce02;
    inBuf[8136] = 256'hf602ec02c2029b029302cb025503260425052b06f8065d073a0781064905ca03;
    inBuf[8137] = 256'h3a02e100fcffa7ffefffc300ef013b036f045605dd050f06fd05cb05a0058305;
    inBuf[8138] = 256'h7d058805860561050805660482037d027d01ba006d00ad008101d70275041e06;
    inBuf[8139] = 256'h93079008ee08a908c7077806ff0491036502a40152016f01f301bb02af03b804;
    inBuf[8140] = 256'hab056c06e706fb06a406f305f904e603fa0263024d02d402e3035105e5064508;
    inBuf[8141] = 256'h25095209a70836074905360373016e005a003f01ee02f504da063508b2084008;
    inBuf[8142] = 256'h14077a05de03af0226025c024703a5042d06a007b1083909320998088b074006;
    inBuf[8143] = 256'he004a303c302580275021f032b046f05be06da079a08ee08c2081e082607f605;
    inBuf[8144] = 256'hc104c8032903fe0251030104e704e405c4066b07d407f407d7079e0756071407;
    inBuf[8145] = 256'hec06cf06b3069906730648062f062a063a0665068b0696067d062b06ac052405;
    inBuf[8146] = 256'haf047704a2042b05fa05f006ce076808b308a8085f080708b20772074f072e07;
    inBuf[8147] = 256'hfe06be0665060206b60589058405b105ff056406e0065807b607ed07de078507;
    inBuf[8148] = 256'h00076f060206ed053806d906b1077f0806092109ab08af0765060b05f3036a03;
    inBuf[8149] = 256'h8c035504a6053a07c808150adc0af20a520a0c096107b8056904bc03d1038104;
    inBuf[8150] = 256'h87059b067107e407f507b1073c07c7066b06410655069306e406330760075e07;
    inBuf[8151] = 256'h3407e4067e061e06d005a405a805ce05ff0526062006e1057e051205ca04d204;
    inBuf[8152] = 256'h3305e205c306a4075a08ca08db088608d607d806a90579047203bc0273029002;
    inBuf[8153] = 256'h0103aa0364041405a9050e0636061e06cb055305db047f0454045b047f04a904;
    inBuf[8154] = 256'hc904d804db04dd04dd04d504bc0480041b049003e9023e02b10166017d010302;
    inBuf[8155] = 256'he80203041405d9052006d305fc04bf034d02da0098ffaefe37fe42fec9feb6ff;
    inBuf[8156] = 256'he2001b023103fd0367046a0413047903bd02060270011101ef00f200f800d800;
    inBuf[8157] = 256'h6f00bdffe1fe0bfe7bfd58fda3fd42fefefe93ffd4ffabff1bff50fe86fdf7fc;
    inBuf[8158] = 256'hddfc52fd42fe86ffde00f901a102aa02f7019700b5fe93fc9dfa37f99af8daf8;
    inBuf[8159] = 256'hc3f9ecfafafbacfceffcf2fcf4fc1bfd80fd08fe6efe7dfe04fee8fc4efb7bf9;
    inBuf[8160] = 256'hbff785f613f670f687f70df99dfaf2fbe0fc49fd42fde3fc3bfc75fbb4fa06fa;
    inBuf[8161] = 256'h88f934f9e1f876f8dbf705f725f678f526f55bf50ff608f713f8f7f877f98df9;
    inBuf[8162] = 256'h3bf983f893f79cf6bff53ef53bf5a6f56ef65af713f86ff850f8a5f799f65cf5;
    inBuf[8163] = 256'h13f403f35ff234f29df28af3b7f4eef5e6f64cf70ff732f6c8f429f3b3f1acf0;
    inBuf[8164] = 256'h73f02ff1b9f2d6f40cf7b5f866f9d7f8f6f624f4f2f0f0edd2eb08eba5eb93ed;
    inBuf[8165] = 256'h62f058f3dcf562f785f768f668f409f204f0deeec1eeb2ef5af123f3a0f46bf5;
    inBuf[8166] = 256'h3af52af473f25ef06eee0aed60ec9eeca7ed1befb3f015f2ecf237f303f362f2;
    inBuf[8167] = 256'h9cf1def02bf0a4ef44efe3ee8dee42eefaedeaed36eedaeeebef47f196f2a6f3;
    inBuf[8168] = 256'h33f401f431f3f6f187f052ef94ee4cee7beeefee4fef83ef75ef11ef8bee07ee;
    inBuf[8169] = 256'h8bed42ed38ed5aedc8ed85ee7aefb1f006f22cf3fdf345f4d9f3ebf2baf17ef0;
    inBuf[8170] = 256'h94ef1deffaee22ef6cefa7efe3ef23f048f05df049f0eaef67efe9ee91eea8ee;
    inBuf[8171] = 256'h3fef2af052f175f241f3a1f383f3d9f2e6f1ebf01cf0ccef0af09ff05cf1f3f1;
    inBuf[8172] = 256'h1ef2f4f19ff148f137f17ff102f2c1f2a5f382f44ef5d9f5daf54bf539f4d9f2;
    inBuf[8173] = 256'ha4f1f2f0ccf027f1aff105f21df20af2f1f11ff2a5f267f35ef471f584f6a0f7;
    inBuf[8174] = 256'ha9f859f98af913f9e9f756f6a5f411f3e0f12df1faf073f1a5f27af4cef635f9;
    inBuf[8175] = 256'h21fb3efc5efc8bfb26fa86f8e4f683f580f4ecf3f9f3b0f4e9f570f7def8d2f9;
    inBuf[8176] = 256'h38fa26fad3f998f9a0f9e4f95ffaecfa60fbaffbb4fb40fb57fa14f9c5f7f0f6;
    inBuf[8177] = 256'hf8f6f2f7b2f9b5fb6afd8cfe11ff22ff09ffdafe73febbfd9cfc30fbd3f9dbf8;
    inBuf[8178] = 256'h7af8c5f897f9b9fa0cfc6bfdb6fed5ffa5000d012001fa00bd0086004c00edff;
    inBuf[8179] = 256'h5bff92feabfdddfc4dfc11fc3efcdffc00feaeffc501eb03a6056f06ff057404;
    inBuf[8180] = 256'h42020b0066fe9bfdaafd65fe8affe8005f02bc03bb04110583041e0339015bff;
    inBuf[8181] = 256'h18fed8fdb6fe8d000803b6052908fb09da0aaa0a8009a8079405af0339025401;
    inBuf[8182] = 256'hfc002b01e9012f03d0047c06ba072408a2076b06f304c0031703f3022d039403;
    inBuf[8183] = 256'h1d04f3043706e107be09620b6a0cb60c4c0c580b1b0aac081607830527045403;
    inBuf[8184] = 256'h67036e0432064d082c0a610bcc0b730b830a4c09fe07cc060206c7052e063507;
    inBuf[8185] = 256'h8b08ce09c20a390b3f0b140bd30a870a460a040ad509f2095e0af90a8b0ba50b;
    inBuf[8186] = 256'h0c0bed09a108ad0793075f08ce09830bf80cd20d030e780d460cb70a09099e07;
    inBuf[8187] = 256'hf40633074708ed098b0ba80c270d0a0d930c290cdf0bb50bb20bb20bb90bf00b;
    inBuf[8188] = 256'h470ca60c020d160dca0c420c890bc50a300ac7099109b8092e0aed0af70b010d;
    inBuf[8189] = 256'hd00d5b0e840e5e0e2b0ee10d790d010d5d0ca50b290bf10af50a200b0c0b8e0a;
    inBuf[8190] = 256'he50959096709810a780cd30e0611571275129311f00ffe0d4b0c020b4e0a640a;
    inBuf[8191] = 256'h1a0b420caa0dc50e2f0fd20e9f0de90b570a4d092709250af30b170e1e105511;
    inBuf[8192] = 256'h601164109e0ea80c490bc70a290b450c7c0d640ef50e240f250f470f660f590f;
    inBuf[8193] = 256'h1c0f8d0edc0d840d9f0d290ef70e6d0f230f2a0ea70c220b4d0a570a3c0bd60c;
    inBuf[8194] = 256'h960e10102211861137117310450feb0dd60c210cf10b740c6f0db70e3d109c11;
    inBuf[8195] = 256'h8a12e6125c12ef100c0f090d690bb10acb0a7b0b890c800d440e150ff40fee10;
    inBuf[8196] = 256'hfd11ac12ac120412b810240fd50de90c660c4e0c4d0c4a0c7b0cdc0c890da50e;
    inBuf[8197] = 256'he40f11112212d9122d134313f31235123011d50f4d0ef70ce20b390b390bc90b;
    inBuf[8198] = 256'he40c8f0e5e10e611d712b8128211ac0fac0d270cb40b490ca10d620fed10ea11;
    inBuf[8199] = 256'h63124c12d5114c11a910ed0f310f4c0e480d680cc10b8a0b090c1b0d920e4510;
    inBuf[8200] = 256'hc211ca125f135613b812a7110f100b0ef90b1e0af008e908010afc0b6a0e8310;
    inBuf[8201] = 256'hb811e8110f11970f230e0c0d990cef0cc10dc30eb60f2f1004104f0f210ecb0c;
    inBuf[8202] = 256'hbe0b210b160ba70b8a0c790d410e7f0e080eef0c480b790915087307c8071009;
    inBuf[8203] = 256'hd40aaa0c540ea00f9f10791105120b1255119e0fff0ce609bc06fe030a02e900;
    inBuf[8204] = 256'h9f003301870289041e07e7098e0cd40e73106411c3119111da10ac0ff40dbb0b;
    inBuf[8205] = 256'h24093a062f034b00d2fd2ffcd5fbeafc5affbb024a065a09820b990cd30c7f0c;
    inBuf[8206] = 256'hb70b830ae008d906c7042a0356025f02fc029503ba034e038002bd0158014c01;
    inBuf[8207] = 256'h65015f011e01d600e10078019a02f203ff046305fa04da035002a7001bffe5fd;
    inBuf[8208] = 256'h2ffd0efd86fd66fe54fffeff2500c9ff25ff7dfe00febdfd9afd7dfd6cfd79fd;
    inBuf[8209] = 256'hbdfd3bfec2fe10fff6fe5ffe68fd50fc3ffb52fa95f902f9a7f89af8cff829f9;
    inBuf[8210] = 256'h7af989f956f91af915f981f956fa32fbabfb84fbbbfab1f9e0f87af87af892f8;
    inBuf[8211] = 256'h58f8a7f7a3f686f5a3f425f4ecf3def3e8f3f5f31ff479f4f0f489f54bf61ff7;
    inBuf[8212] = 256'h09f8e5f854f916f911f856f660f4aef269f189f0c2efb0ee6bed6bec38ec55ed;
    inBuf[8213] = 256'hbbefb4f271f53ff7c3f756f78bf6b2f5f3f41af4c1f2f1f003ef66eda9ecf3ec;
    inBuf[8214] = 256'hd4edd2ee6bef3cef75ee76ed88ec14ec4aec08ed4deeeaef76f1c0f294f3bcf3;
    inBuf[8215] = 256'h63f3b1f292f114f025eeafeb2ae940e772e62fe742e9c2ebe1ed0aef11ef9dee;
    inBuf[8216] = 256'h6deecbeec3efd0f026f184f008ef01ed18ebafe9ade815e8cfe7b8e70fe8f5e8;
    inBuf[8217] = 256'h34eab4eb2bed2ceebeeeefeeaeee37eea0edcfecffeb57ebc5ea6fea4aea0cea;
    inBuf[8218] = 256'hc8e98fe953e954e995e9c7e9e7e9ede9cce9eee995ea9eebefec20ee99ee55ee;
    inBuf[8219] = 256'h7aed31ecfaea0cea37e986e8f1e75de71fe767e710e821e968ea85eb83ec62ed;
    inBuf[8220] = 256'hf2ed4dee66eef8ed2bed1eeccbea89e986e8afe741e74de79fe749e829e9ece9;
    inBuf[8221] = 256'haaea72eb2eec1ded38ee1cefb1efc7ef1feffeed98ecefea51e9e2e79be6dfe5;
    inBuf[8222] = 256'hf1e5c5e672e8b2eae8ecddee5df02ef18df186f1d9f099efc7ed6deb29e98ce7;
    inBuf[8223] = 256'hd6e657e7dce8c5eac4ec85eeb4ef82f002f113f1e5f07df0bcefddeef4eddbec;
    inBuf[8224] = 256'hcbebe2ea26eafbe984ea83ebdbec2eee0def9fef21f0b5f0b2f101f320f4cff4;
    inBuf[8225] = 256'hc6f4cbf32af21cf0afed42eb1ee97ae7f2e6dbe713ea69ed3df1abf450f7ecf8;
    inBuf[8226] = 256'h61f90cf927f8acf6daf4caf27ff061eeb8ec9ceb5deb01ec43ed09eff6f085f2;
    inBuf[8227] = 256'h90f304f4e3f3aff3ccf350f457f592f673f7caf779f77df640f5fff3bff2b7f1;
    inBuf[8228] = 256'hfaf08bf0c0f0b5f131f3fef49cf679f78af7f5f6fef535f5daf4d1f410f55df5;
    inBuf[8229] = 256'h75f575f570f565f58df5f2f57af636f701f88ff8d0f8b2f83af8cef7bcf714f8;
    inBuf[8230] = 256'he0f8cff962fa71fae9f9d4f88cf73ff6f6f4e8f341f32bf305f4e8f595f8b4fb;
    inBuf[8231] = 256'ha2feb800b2017a01280022febdfb35f9e8f610f5cbf352f3aef3c5f499f602f9;
    inBuf[8232] = 256'hbcfb8bfeff009a0227039b0239019aff38fe41fda9fc08fcf4fa68f9aaf739f6;
    inBuf[8233] = 256'ha6f520f675f753f957fb4dfd4bff5b015203df048105d804fe025d00a5fd8ffb;
    inBuf[8234] = 256'h7efa7bfa55fba4fc00fe20ffc1ffc6ff50ff9ffe17fe1dfed1fe080062016002;
    inBuf[8235] = 256'hb8027102c40102016400e2ff64ffdcfe59fe19fe5afe2fff7800ec0134032704;
    inBuf[8236] = 256'hc7041f053e050f0561041f0361017afff4fd46fda3fdfffefa001403ea043c06;
    inBuf[8237] = 256'hf30631071a07d00679061a069d05f7041004e702bc01d4007400c900aa01ba02;
    inBuf[8238] = 256'ha90338046e04a5042a0524068e0716095d0a390b8d0b570bb30a9109e507dd05;
    inBuf[8239] = 256'hb803e501f1001601420230044a060a083b09c409c30990095b0947098609040a;
    inBuf[8240] = 256'ha50a5b0be10b030cbe0bfb0ac4095b08d80667055704ca03e803e904af06fd08;
    inBuf[8241] = 256'h9c0b1a0e2410ac119512de12ac12e0116710690ef60b4d09e706f904a9032803;
    inBuf[8242] = 256'h55032104a805cb07680a680d5e10e712db14fa153816cf15c01424133d11130f;
    inBuf[8243] = 256'hce0cc50a0c09c10727073207e70766096f0bba0d1310fa1121139c136d13cc12;
    inBuf[8244] = 256'h25128211e9107610f90f690fff0eb00e8b0ec00e250fa60f5b100e11a1111f12;
    inBuf[8245] = 256'h461204129311fb1071104d106e10a010c7108610d60f260fc00e0e0f70109f12;
    inBuf[8246] = 256'h231594174919ef19a51964185e16fc135411a10e620cc50a080a760ad40be00d;
    inBuf[8247] = 256'h751017137f15af175f19721afb1ac01ab4191b18fd159f138711df0fdc0ec20e;
    inBuf[8248] = 256'h500f421076117a121e138f13cb13021488143815f015b0162a174d1755172c17;
    inBuf[8249] = 256'hcf1650166315f3134e1297102d0f890e950e250f251038115512c81389158c17;
    inBuf[8250] = 256'hb7196b1b2c1ce01b611af5173b157b120710400e120d800cb20c710da20e5510;
    inBuf[8251] = 256'h3d122d142416c517e018791955197718261760154b133e11420f950da90c8e0c;
    inBuf[8252] = 256'h570d070f161104138e14551565152715c01458141414a713e612f411d210ca0f;
    inBuf[8253] = 256'h4c0f560fd20fa8106511c811de118b11ef105610bd0f3b0f0e0f260f860f4810;
    inBuf[8254] = 256'h2111d7114c1222123f11de0f200e6c0c570b180bca0b650d5c0f291180120913;
    inBuf[8255] = 256'hd41244127e11ad10f20f100fec0dab0c5a0b3a0aa5099209f209b80a900b500c;
    inBuf[8256] = 256'h030d850dd30d070ef80da40d2e0d920cf20b930b740b980b060c7c0ccd0cf20c;
    inBuf[8257] = 256'hc20c460cb00b000b4b0ab2092209a30864086608bc0879095a0a1b0b880b560b;
    inBuf[8258] = 256'h800a4b09e907a006b4052305ec042505be05bf062e08c509310b270c4e0c990b;
    inBuf[8259] = 256'h440a9308ee06b5050105cf040d057105c305e805bf055905ea0491047404aa04;
    inBuf[8260] = 256'h12058a05f50527061206bf052c056f04ad0300038e027802ac020b036e039b03;
    inBuf[8261] = 256'h7f032d03c80287029902ff02a3035a04e6041f05ff048d04eb0334036c028901;
    inBuf[8262] = 256'h7c003effecfdcafc1ffc30fc11fd98fe730039028d033e044904ce0304031902;
    inBuf[8263] = 256'h27013a004dff62fe84fdc1fc2bfcd3fbb3fbc6fb09fc7dfc35fd3ffe90ff0401;
    inBuf[8264] = 256'h5c023a035f03b402510187ffb6fd24fcfcfa38faa7f92af9baf868f86cf8f3f8;
    inBuf[8265] = 256'hf5f94cfba5fc9cfd02fed9fd42fd8dfcf8fb8dfb51fb36fb1ffb1bfb39fb6ffb;
    inBuf[8266] = 256'hbdfb03fc09fcc3fb3bfb78faacf9fbf861f8e8f78ef737f7f8f6dff6e1f611f7;
    inBuf[8267] = 256'h70f7e0f765f8f0f856f990f990f93cf9b4f81cf880f711f7e3f6daf6fdf647f7;
    inBuf[8268] = 256'h96f7f3f74df865f82ff89ff7b0f6b1f5f4f49bf4cbf462f5fcf565f677f61af6;
    inBuf[8269] = 256'h8ef511f5abf479f46df450f425f4f2f3abf386f39cf3cff32af495f4d3f4edf4;
    inBuf[8270] = 256'heef4c5f4a3f499f488f487f49af4a4f4caf40df52bf507f56bf41bf356f183ef;
    inBuf[8271] = 256'h07ee7bed21eeb5efe2f116f49df53af6eaf5c6f459f319f234f1eef03af1b6f1;
    inBuf[8272] = 256'h3af28af260f2dbf118f118f020ef5aeebeed8fedeaedb3eefcef9ff131f38bf4;
    inBuf[8273] = 256'h76f5aff55df5a3f47ef333f2dff06def15eefdec24eccdeb0eecafecaaedcdee;
    inBuf[8274] = 256'hb1ef4ff09af073f01af0c1ef6def67efc2ef49f0fbf0acf103f208f2bdf10af1;
    inBuf[8275] = 256'h30f052ef60ee94ed0bedb5eccfec66ed3dee4fef68f026f18af18ff11af166f0;
    inBuf[8276] = 256'h90ef83ee7beda2ecfaebd1eb45ec1ced42ee6bef22f064f03cf0b1ef27efdaee;
    inBuf[8277] = 256'hbaeeedee69eff5efa5f06bf1fbf14ef23bf282f151f0e3ee62ed45ecd0ebebeb;
    inBuf[8278] = 256'h9beca2ed8eee49efc1efdeefeeef23f06cf0ddf04ef163f11ff188f0a6efe0ee;
    inBuf[8279] = 256'h7eee7deef8eec6ef82f014f161f149f10ef1dcf0a6f08cf07ef042f0f8efc5ef;
    inBuf[8280] = 256'hb4ef0cf0d4f0bdf19ef235f33ef3edf27cf2fef1b0f189f142f1d9f049f093ef;
    inBuf[8281] = 256'h0cefecee2cefdcefd3f0b3f167f2def207f329f373f3dff37ff42ef593f5a2f5;
    inBuf[8282] = 256'h57f5b4f40af48bf330f30ff314f30ef319f341f374f3c9f325f445f425f4c4f3;
    inBuf[8283] = 256'h27f399f24bf242f299f23ef3f7f3c2f48cf52ef6b4f611f726f70ef7dcf699f6;
    inBuf[8284] = 256'h85f6c2f647f71af80ef9d0f934fa09fa2df9d2f73bf6a4f469f3b8f286f2e1f2;
    inBuf[8285] = 256'hbef308f5caf6e4f8f8faa6fc73fd00fd6afb1df9b2f6e6f42ef499f402f608f8;
    inBuf[8286] = 256'h33fa45fc06fe43ffeffff7ff49ff02fe4cfc5dfa90f82ff769f668f61ef74bf8;
    inBuf[8287] = 256'ha6f9d8faa4fb15fc5afcb0fc50fd32fe10ff99ff85ffc4fe9efd78fcaffb75fb;
    inBuf[8288] = 256'hb2fb1afc73fc9efcb0fceffc89fd7cfe97ff8100f100d9005900beff5dff66ff;
    inBuf[8289] = 256'hd6ff8600320198018c0101011a001bff4cfee7fdf4fd48fea2fed3fedffe08ff;
    inBuf[8290] = 256'h9dffc800680211043c0599052b0548046903db0299026b02040248017400f4ff;
    inBuf[8291] = 256'h2a004a0124033d050e071e08350873071e0690042f033202ab019601ce012d02;
    inBuf[8292] = 256'ha9023603cf0381043305c5052a065506550660069406f3067007ca07cd077e07;
    inBuf[8293] = 256'hf70676064e0691062007cb0742085b083008dd07870756073007ef0692061606;
    inBuf[8294] = 256'ha0057e05c8057a06840792085f09da09f909db09c809d309f8092f0a380aec09;
    inBuf[8295] = 256'h6c09d90879089e084109220afc0a650b340ba30af4097b098009de09460a8a0a;
    inBuf[8296] = 256'h6d0afa098209360934098f090a0a730ad70a370bae0b710c550d100e620ef00d;
    inBuf[8297] = 256'hab0cf40a3409e80788070a082709930ace0b940cfe0c1a0d160d380d710da60d;
    inBuf[8298] = 256'hd60dcd0d7a0d090d7a0cdb0b560bd70a5f0a210a230a760a3f0b400c2a0dce0d;
    inBuf[8299] = 256'he40d730dde0c610c340c7d0cea0c1d0df60c4c0c490b630ad109bf09530a500b;
    inBuf[8300] = 256'h770cb10db60e610fc70fcf0f810f0c0f690ea20de90c340c930b350b020be40a;
    inBuf[8301] = 256'he60ada0abc0abe0adb0a1a0b900bfb0b300c3d0c160cdd0bde0b170c7d0c140d;
    inBuf[8302] = 256'h9d0dfe0d580e970ebf0ee80ee00e850ee70dec0cac0b770a6909ae088708da08;
    inBuf[8303] = 256'h8a098a0a7f0b2f0c960c970c4c0cff0bb90b870b880b8f0b8a0b980baf0bdd0b;
    inBuf[8304] = 256'h430cb30c080d3c0d180d8f0ccf0bd40abc09cb081208c0071608fd084f0adc0b;
    inBuf[8305] = 256'h2f0dff0d4f0e150e7d0dc80ce80bd00a92092b08d7060a06ee059106d9074709;
    inBuf[8306] = 256'h6a0a190b380bfb0ac60aaf0ac30a010b2b0b250b0c0bdc0aa60a830a460ad309;
    inBuf[8307] = 256'h3c097808b107320705073007b6075908ef087409c109da09e509d909c209b009;
    inBuf[8308] = 256'h7609f7083e08420739067d0535057d0551065f0762083d09c509f809ef099709;
    inBuf[8309] = 256'hfe085208b5076707a5074b080f099609740992083b07ca05b1043f045304ad04;
    inBuf[8310] = 256'h1005410550058105f605c206ce07ba08390929097d086b0750065c05b8047b04;
    inBuf[8311] = 256'h8e04e60489055a064a073908d708eb085e082d0799050b04d5023f026002f702;
    inBuf[8312] = 256'hb60352048c0472044b045904d704c305cb068c07c20752078006b1052505ec04;
    inBuf[8313] = 256'hcf04680483033902e20005000700e5005802eb032605e5054a068d06e8065707;
    inBuf[8314] = 256'h950750074f06890453023300a5fe07fe67fe7dffe400310218039503cc03e903;
    inBuf[8315] = 256'h11043c043e04f4035b039702fb01ca011202a8022a033303a00294016b0093ff;
    inBuf[8316] = 256'h4aff86ff0d009200e70021017101fd01c70292030304d603f3028a010400c1fe;
    inBuf[8317] = 256'hfbfdbafdd0fdfffd2afe4bfe82fe01ffd3ffde00e901a002c50253026a015600;
    inBuf[8318] = 256'h6affd3fe98fe9cfea7fe96fe69fe28fef0fdd8fdd1fdc3fd99fd42fdd9fc93fc;
    inBuf[8319] = 256'h97fc01fdcefdc7feb4ff6600ba00b6006e00e2ff18ff15fed7fc80fb4dfa6cf9;
    inBuf[8320] = 256'h0cf93ef9d8f9b7fab6fbadfc8cfd48febcfed4fe87fecbfdc7fcaefbabfaf2f9;
    inBuf[8321] = 256'ha3f9b5f928fae9fac0fb83fc0afd2dfdf5fc82fce9fb55fbd7fa59faddf969f9;
    inBuf[8322] = 256'h01f9c5f8c4f8e0f800f9fff8b9f847f8dcf7a5f7daf78cf893f9c9faf9fbe2fc;
    inBuf[8323] = 256'h6ffd96fd48fda0fcb5fb89fa3ef9e8f78af646f53ef48cf366f3e5f3f5f47af6;
    inBuf[8324] = 256'h36f8c7f9f7faa3fbb5fb4efb8ffa82f94af8fbf6a0f572f4aff379f3fff339f5;
    inBuf[8325] = 256'he2f6b8f864fa8ffb24fc1ffc7dfb68fafcf844f772f5bff356f27ff15df1e1f1;
    inBuf[8326] = 256'hfaf26ff4e6f52ef720f895f8a1f860f8e5f76bf714f7dff6ddf602f729f749f7;
    inBuf[8327] = 256'h54f72af7d3f64af685f5abf4e5f34ff323f371f319f404f5fdf5c4f651f79ef7;
    inBuf[8328] = 256'ha4f783f73ff7ccf63ff6a9f517f5bcf4b9f403f595f53df6b2f6daf6aaf624f6;
    inBuf[8329] = 256'h81f5eff47df445f448f474f4dbf478f52cf6e6f677f7a6f778f707f776f60cf6;
    inBuf[8330] = 256'he2f5e0f5eff5eaf5b5f577f55df57cf5ebf58af610f758f744f7d3f63df6b3f5;
    inBuf[8331] = 256'h4bf525f53bf56bf5b4f50ff671f6f0f687f713f886f8b7f87af8daf7faf606f6;
    inBuf[8332] = 256'h53f513f54df5fbf5e7f6c9f785f808f94af965f95cf917f992f8c3f7adf68cf5;
    inBuf[8333] = 256'ha2f41ef434f4e1f4f4f546f7a0f8cdf9c0fa68fbb0fba1fb3cfb88fab5f9e6f8;
    inBuf[8334] = 256'h2ef8a6f74bf709f7ecf6fdf645f7ddf7b6f89bf95efacbfac0fa5afac5f931f9;
    inBuf[8335] = 256'hd6f8cbf805f980f923facbfa66fbcffbdffb95fbfdfa31fa70f9e9f8b4f8e9f8;
    inBuf[8336] = 256'h80f95ffa6ffb85fc5bfdbffd85fda7fc64fb15fa17f9baf80ff9e7f901fb14fc;
    inBuf[8337] = 256'he7fc70fdb4fdbefda5fd71fd23fdcffc87fc5cfc69fcb0fc19fd86fdc7fdaefd;
    inBuf[8338] = 256'h2ffd5bfc5dfb83fa10fa24fac7fad8fb1efd6afe92ff7e002b0190019e015601;
    inBuf[8339] = 256'hb900caffa6fe70fd4efc6cfbe6facafa24fbe6fbf0fc22fe51ff52000c017301;
    inBuf[8340] = 256'h85015101ec006500d1ff44ffcffe86fe70fe84feaefed2fedcfecffec4feddfe;
    inBuf[8341] = 256'h3affdbff9d004e01c201df01b0015301e4007700060086fff8fe6ffe0bfef1fd;
    inBuf[8342] = 256'h37fedcfecbffdd00e401ba0242036e034203d8024e02c1013f01c5004600bbff;
    inBuf[8343] = 256'h2dffbafe88feaafe1effc3ff6d00f200450175019901c8010c025f02b302f902;
    inBuf[8344] = 256'h260338032503e3026c02cc0118017200f3ffa2ff71ff4bff24ff08ff21ff92ff;
    inBuf[8345] = 256'h7000a601f5021004b904ca04500470035c0242014a008eff23ff1eff83ff4400;
    inBuf[8346] = 256'h43014a022803b403d60399031c038302f0017c012701e500a5005500f4ff96ff;
    inBuf[8347] = 256'h4eff39ff6effedffa90083015002f1025d039403b203d8030a043b044604f603;
    inBuf[8348] = 256'h2c03f401790006ffe9fd50fd4dfdd2fdb2fec5fff10015021c03f3037f04ad04;
    inBuf[8349] = 256'h7604d903f002e901f1003900e6fffbff6500ff009601050243024d0234020c02;
    inBuf[8350] = 256'hd80198014b01eb0086003800180039009f002d01be0134027302800277026a02;
    inBuf[8351] = 256'h6402600244020402ac015401260142019b010c02690283025002e7016101dd00;
    inBuf[8352] = 256'h73002000e6ffd0ffe3ff2a00ad005c012a020803db038c0405051f05c004e803;
    inBuf[8353] = 256'ha5022b01c7ffb7fe2dfe3ffed6feccfff50014020203ad0303040404c1034503;
    inBuf[8354] = 256'ha70208027a011501ef0000013a018f01e30124024f025b02510245023c024102;
    inBuf[8355] = 256'h62029102ba02ce02b0025e02f3018f015b017001bf0122027702980285026102;
    inBuf[8356] = 256'h4b0257028b02c602ef02070313032e037003c603ff03eb035f0366024c016600;
    inBuf[8357] = 256'h04005600370158026503160452043e040404d503d003e503f903fc03db03a003;
    inBuf[8358] = 256'h710360037203a103c503bd037e030a0381021c02fc013002b50266031604af04;
    inBuf[8359] = 256'h19055605770578054b05ee0458049603da025602360297025e03570457052906;
    inBuf[8360] = 256'hb90610072a0700079006c905b20477034b02680105012c01d501f3025e04ec05;
    inBuf[8361] = 256'h7107aa085c096a09ce08ab0753060b0505046b0339036303de0385043605dc05;
    inBuf[8362] = 256'h4e0678066e063f060106cf05a70582056a0565058105d7055c06f1067707c207;
    inBuf[8363] = 256'hb9076f07f3066106de057805350525053e057805d5054406b40622077c07ae07;
    inBuf[8364] = 256'hb1076f07e9064306a0052d051a0569050206c5067e070608570866083008c407;
    inBuf[8365] = 256'h26076506b20531050b055e051206ee06b70727081a08a407ea06240697055b05;
    inBuf[8366] = 256'h7205d4055b06e10656079f07b307a70781074b071807dc0689062806be056605;
    inBuf[8367] = 256'h50058405ef057106cc06dc06b306740650066d06b406f106fc06bb063e06c405;
    inBuf[8368] = 256'h730555055e055c053105ea04a3048604bc043a05de058c061907680774073307;
    inBuf[8369] = 256'ha906f60535058d042404f703eb03ee03ed03ee0315047104f7048905eb05f605;
    inBuf[8370] = 256'hb5054105c50469042a04f703cf03b603c50319049e042005660538059304b103;
    inBuf[8371] = 256'hdc02530235026302ab02f3022a035f03b30326049d04f204f4049104e5031703;
    inBuf[8372] = 256'h5b02ea01d10106027302ea02410366034e030503ae025d021c02ef01c1018901;
    inBuf[8373] = 256'h5a0148017001dd017102f8023f031d039f0202028101440153018601a901a001;
    inBuf[8374] = 256'h67011d01ed00e400f5000c010e01f900e400e600090143016e016a013401dc00;
    inBuf[8375] = 256'h86005200450050005b004f002800f7ffcdffb8ffc2ffe5ff1900530080008d00;
    inBuf[8376] = 256'h71002900ccff7cff53ff58ff7fffa7ffb7ffadff9cff9fffbbffd7ffd0ff89ff;
    inBuf[8377] = 256'hfdfe50febafd65fd5dfd8afdccfd0ffe57feaffe22ffa6ff170050003d00e6ff;
    inBuf[8378] = 256'h6affe6fe6efe03fe98fd24fdabfc36fcdafbaffbcbfb40fc11fd29fe57ff5700;
    inBuf[8379] = 256'he000ce002f0036ff2afe44fd8efcf7fb64fbcffa5bfa45fab4faacfbf4fc29fe;
    inBuf[8380] = 256'hf1fe1fffb9fefdfd38fd99fc35fcfffbdbfbc0fbb8fbd1fb1bfc94fc19fd87fd;
    inBuf[8381] = 256'hc3fdb9fd73fd09fd8bfc10fca7fb4efb0cfbe2fac0faa3fa8ffa86faa1faf7fa;
    inBuf[8382] = 256'h84fb34fcdafc39fd35fdd5fc39fca4fb4dfb40fb75fbcffb1dfc45fc3efcfafb;
    inBuf[8383] = 256'h88fbf7fa55faccf982f97ff9c8f94dfae2fa72fbf3fb56fca0fcc5fca1fc2afc;
    inBuf[8384] = 256'h6ffb89fabbf942f930f97ff90bfa95fa07fb5bfb8dfbb1fbc9fbbdfb8afb38fb;
    inBuf[8385] = 256'hcafa65fa28fa0ffa20fa50fa81fab5faedfa0ffb1dfb0ffbd3fa79fa1bfac1f9;
    inBuf[8386] = 256'h90f998f9c7f91bfa8afaf3fa50fb94fba1fb80fb36fbbbfa2cfaaaf939f9f6f8;
    inBuf[8387] = 256'hf2f822f98ff92cfacbfa5efbcefbf7fbe5fbaafb45fbd4fa66faedf97af91bf9;
    inBuf[8388] = 256'hccf8b3f8e4f84cf9e4f990fa12fb56fb59fb18fbbefa6cfa22faeff9d0f9a3f9;
    inBuf[8389] = 256'h78f963f965f997f9fef970faddfa2afb2efbf9faa2fa31fad7f9aef9a5f9c0f9;
    inBuf[8390] = 256'he6f9e9f9d3f9b8f9a1f9b9f906fa5bfa9afaa2fa56fae8f993f96df994f9f4f9;
    inBuf[8391] = 256'h45fa6ffa6afa32faf7f9d5f9b9f9a9f99df97ef96bf977f98ff9b7f9e1f9eef9;
    inBuf[8392] = 256'hf2f9fef909fa23fa43fa45fa37fa2ffa27fa37fa55fa4dfa15faacf91af9a7f8;
    inBuf[8393] = 256'h84f8abf819f9a3f904fa2efa26faecf9adf986f971f989f9d3f934faa9fa15fb;
    inBuf[8394] = 256'h37fb06fb82fab2f9def843f8f0f7f9f751f8c7f85bf907fab5fa68fb02fc40fc;
    inBuf[8395] = 256'h0ffc6bfb61fa3ef948f89bf75af77df7dbf772f838f90bfae2fa9bfbfcfb00fc;
    inBuf[8396] = 256'habfb09fb59fac8f95ff939f955f998f905fa8afaf6fa36fb30fbcdfa31fa8bf9;
    inBuf[8397] = 256'hfcf8bdf8dcf838f9c6f965fae9fa50fb92fba1fb94fb7bfb53fb32fb16fbe5fa;
    inBuf[8398] = 256'ha4fa56fafbf9c3f9c6f9f6f94efaaefaecfa0cfb20fb3afb80fbedfb55fc9efc;
    inBuf[8399] = 256'habfc66fcf4fb7efb20fb00fb1bfb51fb8efbb8fbb3fb91fb68fb4cfb63fbb1fb;
    inBuf[8400] = 256'h16fc78fcb0fc9efc5bfc0ffcdafbe6fb2efc88fcdafc0dfd1cfd26fd3efd5cfd;
    inBuf[8401] = 256'h78fd72fd30fdc9fc61fc20fc2cfc87fc0bfd98fd06fe37fe38fe1bfeeffdcffd;
    inBuf[8402] = 256'hc4fdcdfdedfd10fe20fe15feedfdadfd79fd70fd9dfdfbfd65feb3fed0febbfe;
    inBuf[8403] = 256'h8ffe7efea2fef7fe6bffd2ff0f001d000700e0ffb9ff8bff4eff03ffb6fe80fe;
    inBuf[8404] = 256'h7dfeaffe05ff5fff9dffb4ffb7ffbfffe3ff2d008c00ec003901620166014101;
    inBuf[8405] = 256'hec007100e6ff6eff39ff65ffeaffa8005f01d401f401cb017c0139011e012b01;
    inBuf[8406] = 256'h5e01a201e901330275029602850232029e01ea003e00c4ffa1ffd1ff4200e900;
    inBuf[8407] = 256'hb001840261032e04c4040705db04410464037602ab0136011a014701b1013602;
    inBuf[8408] = 256'hbd024703bf030e042f040d04a803230396022202ef0101024c02cc026103ec03;
    inBuf[8409] = 256'h6804bb04db04db04c1049504720450041f04e60390032003bd027a026e02b902;
    inBuf[8410] = 256'h4703ff03d5049805270684069b066406fb056605bc042b04be0382038d03c003;
    inBuf[8411] = 256'h010451049204be04f20429055f05a705e50509061c061306f305de05c705aa05;
    inBuf[8412] = 256'h98057a054b052d05220534057e05e8055c06d9063b0771078a076d0715079e06;
    inBuf[8413] = 256'h02065605d70494049b0401059c054406ec066607a507c907cf07c307cf07e507;
    inBuf[8414] = 256'hfb0716080808b90740079c06f20595059c051106f106f107c70855096b091109;
    inBuf[8415] = 256'h8c08f4076d0726070607fd061a073f076507a607ea07230865089608b408e008;
    inBuf[8416] = 256'h020914092c092f091a0910090009e108c0087f081708b507640741077507d707;
    inBuf[8417] = 256'h4708c5082a097b09e2094b0a9a0abf0a820ade091a096208f5070d087d080409;
    inBuf[8418] = 256'h7c09a20972092309c60877085c085208480852085b0867089808de083809c209;
    inBuf[8419] = 256'h5f0a000ba40b080cfe0b860b8f0a3f09f507df062806fa052c069f064d071108;
    inBuf[8420] = 256'he108cc099f0a350b860b670bdc0a210a4b097908dd0766070e07e806e106fc06;
    inBuf[8421] = 256'h5007c2074a08f5089b09270a9c0acc0a9c0a1a0a41093708430780060606ed05;
    inBuf[8422] = 256'h0c0645069c06f8065d07df075b08b208e008c2086108f7079f0776079007bb07;
    inBuf[8423] = 256'hcd07b6075b07ce064806dd05a305b205e8052d068606d2060807390757075f07;
    inBuf[8424] = 256'h600744070507af0632069a0511059e04570456048504cf0432059205e7054006;
    inBuf[8425] = 256'h8e06cd06fc06f606ae0633068305bc0411049103490343036a03b3032404ab04;
    inBuf[8426] = 256'h3b05c60520062a06e10546058204d303550316031a033d0366038d03a403ad03;
    inBuf[8427] = 256'hb003a3038a0375036a037903af03f503330451042f04cf035003d10274025202;
    inBuf[8428] = 256'h63028e02bb02ce02c202a5027a0250022d020502d901b801aa01bb01f5014c02;
    inBuf[8429] = 256'had0202033b03540349030f03a302070244017c00dbff83ff80ffc2ff25008300;
    inBuf[8430] = 256'hc700ee0006011d013b0163018e01ba01ea011d0242023e02f10148014b0019ff;
    inBuf[8431] = 256'hf1fd13fda6fcb8fc3dfd12fe15ff28002901fc01810292021d022d01e6ff88fe;
    inBuf[8432] = 256'h53fd6efceffbd0fbfafb66fc15fdf6fdf9fefcffc2001c01f5004f0054ff37fe;
    inBuf[8433] = 256'h1ffd39fc98fb39fb21fb51fbadfb25fca8fc18fd71fdaffdc5fdb8fd85fd20fd;
    inBuf[8434] = 256'ha2fc29fcc9fba6fbc2fbf3fb18fc0dfcb5fb2dfbabfa5bfa64fac3fa40fbb5fb;
    inBuf[8435] = 256'hf9fbf4fbc9fb9efb7bfb67fb4afbf5fa66fab2f9f1f85ff822f82ff87df8eef8;
    inBuf[8436] = 256'h59f9bef91dfa69fab1faf3fa10fb0dfbe1fa71fac8f9f8f807f82bf796f665f6;
    inBuf[8437] = 256'hb7f67df774f86ef92dfa72fa4afad5f927f974f8dbf74ef7ddf68ff662f67bf6;
    inBuf[8438] = 256'he6f680f72df8b1f8bdf853f88ff79cf6dcf59af5def5aaf6d0f7f9f8f0f983fa;
    inBuf[8439] = 256'h81fafff91cf9eaf7aef693f59bf4e8f38af378f3d2f3a5f4c5f516f756f826f9;
    inBuf[8440] = 256'h71f939f997f8e2f759f7fdf6d8f6c7f68ff63df6f1f5bdf5d9f552f6e7f666f7;
    inBuf[8441] = 256'h92f734f773f689f5acf432f441f4baf498f5bcf6e3f7faf8def94cfa3bfaa7f9;
    inBuf[8442] = 256'h8ef830f7c6f56df461f3baf26af28df224f305f431f596f6fff765f9b0faa7fb;
    inBuf[8443] = 256'h2efc17fc2bfb87f962f7fdf4dcf260f1a9f0d7f0d5f155f32cf525f7edf868fa;
    inBuf[8444] = 256'h73fbddfbb8fb13fbf8f9a4f848f7f6f5e9f444f4fef330f4cef496f565f60af7;
    inBuf[8445] = 256'h47f728f7d3f670f659f6bcf682f795f8aff96cfab0fa77fac4f9d8f8ebf709f7;
    inBuf[8446] = 256'h5bf6f7f5cef5f6f564f6eaf674f7d6f7ddf7a6f759f70ef708f761f7eef791f8;
    inBuf[8447] = 256'h1bf95af960f949f928f929f94bf95ef953f90ff975f8a7f7d2f612f6a9f5c3f5;
    inBuf[8448] = 256'h5ff680f7fef882fad1fbb1fcecfc98fcd2fbabfa5ff911f8cdf6cbf537f51df5;
    inBuf[8449] = 256'h9bf5acf61df8c6f96efbccfcbdfd1bfebcfdb1fc1efb38f974f73ff6ddf57ef6;
    inBuf[8450] = 256'h04f800fafcfb82fd36fe14fe48fd19fce7faebf92ef9c4f8a7f8bff816f9aef9;
    inBuf[8451] = 256'h6afa3efb16fcd3fc72fde3fd06fecffd2bfd15fcc8fa8df9a6f85df8ccf8d0f9;
    inBuf[8452] = 256'h40fbe1fc70fec1ffa700f30095008dfff8fd29fc7dfa3ff9b6f8f4f8d7f934fb;
    inBuf[8453] = 256'hd0fc68fecfffe00075017a01e100aeff0ffe47fca7fa90f944f9d4f92ffb10fd;
    inBuf[8454] = 256'h0dffcb00010280025602b301d90008005dffd4fe55febbfdfefc4bfce9fb15fc;
    inBuf[8455] = 256'hf2fc67fe1b00a201a302f502a702eb01fe00120041ff96fe23fef2fd0afe6dfe;
    inBuf[8456] = 256'h11ffd7ffa2005901ea01460261023a02d2013a0193000600aeff96ffb9ff0100;
    inBuf[8457] = 256'h5500ab000a017b01fd018802090363037b034703c402f801f900e4ffe3fe2cfe;
    inBuf[8458] = 256'heefd48fe3dffb0006c022f04aa059e06dd064506dd04e302b900d8feb4fd8ffd;
    inBuf[8459] = 256'h66fef0ffb40142034d04b8049f044904ed03b403b103c803ca0393030d034502;
    inBuf[8460] = 256'h6d01c4008200c1006301340201039703ea031604280424040b04c3033a038302;
    inBuf[8461] = 256'hc5013e012d01ac01b60223049905be06580735075706f6045103b8017f00d1ff;
    inBuf[8462] = 256'hc4ff5c007601df026704c705c606420715074306040591033c0263012d019301;
    inBuf[8463] = 256'h6e026b034304d604150517050705e704ba049004600438043c046804ad04fd04;
    inBuf[8464] = 256'h3405430534050605be046804fa03880348034e03a4033804b404c6046104a303;
    inBuf[8465] = 256'hee02c5026103af045406ae074b080f081507bf058f04c7037b039f03ee032a04;
    inBuf[8466] = 256'h3c040f04bc038903a50337044a059e06e207d0081e09c208e707a40611054f03;
    inBuf[8467] = 256'h69019aff5ffe33fe77ff3b02ed05a109630c690d900c5e0a990712055d037902;
    inBuf[8468] = 256'h1b02f901da01d5013e024b03fe0419070109220a300a12091e07fe0446036402;
    inBuf[8469] = 256'h8c027a03af04a805ef056d057304740300038403ed04d606b408df09f209f108;
    inBuf[8470] = 256'h1707da04cd024d019900d600e8019b03b005ba075e09680aa20a060ac7080807;
    inBuf[8471] = 256'h0105100380019f00ae0098011003ab04e0056d0674063e063906bb06a3078f08;
    inBuf[8472] = 256'h1509c9089107c305cf03330255014501df01e9020404f804c3056406f906ab07;
    inBuf[8473] = 256'h5b08c808b608e9076d06a9041e034802660234033404ef040a0596040b04d503;
    inBuf[8474] = 256'h3f045305b206e00782085d08760713067e040e031b02ca012902250363048005;
    inBuf[8475] = 256'h3b0669061a069d052a05e104cb04c604c104da042c05d305c3069b07e6075207;
    inBuf[8476] = 256'hc50592036a01eeff83ff4300d701bd038805e206ac07f007ad07f706f205b404;
    inBuf[8477] = 256'h70037402ec01f501a102ca03280565061607f60607068e0419034b0271027003;
    inBuf[8478] = 256'hd004d205ed051705af0354029f01b601540204035e034c031603100377034c04;
    inBuf[8479] = 256'h3205c805e1058005e00457040704e603d3039a0325038a02f1018b017e01ca01;
    inBuf[8480] = 256'h560201039003dd03ec03d203b803d3032a049304ce049204c403870227010500;
    inBuf[8481] = 256'h6bff64ffdbffc000f90175032305b906c207ca0790063c046d01f6fe97fdabfd;
    inBuf[8482] = 256'hf7fed7009402a403e703ae03640352038403b5038403bd0276011b003fff4cff;
    inBuf[8483] = 256'h55000c02cb03e604ff0419049c0222012600d5ff07005b007a00510011001700;
    inBuf[8484] = 256'hb300e5015a038d04fc04720428039e016700eaff2b00d30064017501e200deff;
    inBuf[8485] = 256'hd4fe3efe6ffe6fff0401cb025104340547058e0432037e01c5ff55fe66fd14fd;
    inBuf[8486] = 256'h5efd29fe3eff60005401f0012a021c02f501e001f201210243022602ad01e700;
    inBuf[8487] = 256'h01003affc7fec2fe21ffb9ff5a00de0025012201d9005c00c6ff41fff5fefefe;
    inBuf[8488] = 256'h62ff0e00d8008b01f101e5015a015f0027fffffd38fd10fd99fdaefefaff2401;
    inBuf[8489] = 256'he8012e020e02be0166011a01cc006400d1ff11ff37fe6bfdcefc78fc7afcd7fc;
    inBuf[8490] = 256'h77fd39fef5fe83ffdeff1b006200d8007b011c02720235024701d4ff37fecffc;
    inBuf[8491] = 256'hebfba4fbd7fb4efcd8fc5cfde1fd75fe1effd7ff8300f7001601d10023002cff;
    inBuf[8492] = 256'h1afe1cfd67fc20fc47fccdfc85fd35feb1fedbfeaafe36fea8fd2afdf2fc1cfd;
    inBuf[8493] = 256'ha0fd64fe2dffafffbaff47ff73fe89fdd3fc79fc7dfcacfcb7fc72fcd7fb14fb;
    inBuf[8494] = 256'h8efaa8fa92fb49fd7cff9a0118038e03d00209019efe0bfcccf92af83af702f7;
    inBuf[8495] = 256'h72f76ff8f0f9d7fbd6fd8dff9b00bd001000fcfe06fea1fde1fd67fea9fe27fe;
    inBuf[8496] = 256'hb3fca8fab1f874f75ff772f83dfa36fce9fd09ff96ffadff66ffdffe2afe54fd;
    inBuf[8497] = 256'h83fcd7fb58fb0ffbf1fad9fac2fab1faaafac3fa0dfb80fb16fcb7fc37fd77fd;
    inBuf[8498] = 256'h60fdedfc55fcddfbbefb28fc04fdedfd7dfe64fe84fd15fc81fa2cf968f847f8;
    inBuf[8499] = 256'haef88df9c9fa3cfccafd2efff4ffc8ff87fe5dfce9f9fef745f714f82afab8fc;
    inBuf[8500] = 256'hcdfe98ffc2feb2fc42fa62f8d5f7ccf8cdfa1bfdf2fec9ff95ff9ffe44fde6fb;
    inBuf[8501] = 256'hb6fac1f925f9fef851f924fa3dfb2cfc98fc53fc71fb65fab9f9c5f9a1fa09fc;
    inBuf[8502] = 256'h74fd65fe89fecefd80fc04fbb4f9e8f8c0f814f9bdf98bfa49fbeefb82fc04fd;
    inBuf[8503] = 256'h7bfdcefdcbfd62fd90fc6afb3dfa52f9c9f8baf814f9a8f967fa49fb3bfc2ffd;
    inBuf[8504] = 256'hf4fd3bfed4fdb2fc07fb5af939f8f7f7acf80afa74fb6efcb6fc53fca1fb0dfb;
    inBuf[8505] = 256'hd1fafafa52fb7cfb47fba9fabef9e5f878f8acf8a0f934fb05fdaffec4ffebff;
    inBuf[8506] = 256'h17ff77fd5bfb37f967f71cf67df58cf533f673f73bf94dfb69fd3aff5e00a300;
    inBuf[8507] = 256'hffff90feb1fcc3fa18f900f89bf7d0f77cf860f92ffad1fa46fb9dfb00fc80fc;
    inBuf[8508] = 256'h00fd5bfd5cfdd8fce6fbb2fa73f977f8eef7e3f76af882f90dfbe2fcacfef1ff;
    inBuf[8509] = 256'h49006cff5cfd8dfaabf76bf571f402f5eef6c3f9d5fc6fff1b01a0010801abff;
    inBuf[8510] = 256'hf6fd42fcdafad9f92ef9cbf89ef89bf8dcf86df944fa5efba3fce5fd03ffd3ff;
    inBuf[8511] = 256'h2300d4ffd0fe22fd17fb1af999f7faf65cf788f822fab8fbeefcb4fd30fe98fe;
    inBuf[8512] = 256'h1bffb7ff33004a00c1ff8dfeeffc47fbf0f93cf942f9dcf9d6faf5fbfafcc5fd;
    inBuf[8513] = 256'h44fe70fe55fe01fe85fd0afdabfc79fc8bfcdffc57fdd9fd43fe79fe80fe70fe;
    inBuf[8514] = 256'h65fe79fea5fec5feaffe4afea8fd10fdccfc07fdbdfda3fe44ff52ffc6fee0fd;
    inBuf[8515] = 256'h16fdd4fc46fd44fe66ff39007f0038009eff0affb2fe94fe8cfe64fef7fd5dfd;
    inBuf[8516] = 256'hd8fcb3fc1bfd06fe32ff4000da00e50089000c00b6ffb5fffeff550085007800;
    inBuf[8517] = 256'h3b000100f9ff33008900b4007700c6ffccfee9fd8bfdecfdf9fe6000a4015a02;
    inBuf[8518] = 256'h5702bd01e4003100edff2c00c5007101f0011602cf01210129000afff0fd20fd;
    inBuf[8519] = 256'he7fc84fd0cff5501f2034206ad07d407ad068604f20184ff9ffd6dfce0fbcefb;
    inBuf[8520] = 256'h1cfcd1fc13fefeff73021d057207d408de089a0772050a030b01d5ff62ff62ff;
    inBuf[8521] = 256'h74ff60ff36ff36ffabffb60025029f03cf047a059a055a05de042f044a032902;
    inBuf[8522] = 256'he200baff01ff00ffcbff2c01c9024404410590053b055304020389012b002cff;
    inBuf[8523] = 256'hcafe1dff1b0099014c03f1045a065c07e507f30776076f0602055803ab014500;
    inBuf[8524] = 256'h59ff04ff4eff23006701fc02a30423064707d407b3070407f705cb04c503fa02;
    inBuf[8525] = 256'h6502f60198014e0139016201d1017e023703df038404340507060707f9078208;
    inBuf[8526] = 256'h5108390762054b037f017a0073003201530279034c04bc04f104080511051505;
    inBuf[8527] = 256'hf904b7046c043b045504e204c805d306c3073d0812084a07fd056804e602b601;
    inBuf[8528] = 256'h0a0105019a01ac0218049705f9062008e20832092309b008ec07030707061005;
    inBuf[8529] = 256'h3b048103d8024102b30150015401db01f50295045e06eb07020977095c09ee08;
    inBuf[8530] = 256'h4b087e0788065305ff03e40252029202b4035105e306ff075608f90742078106;
    inBuf[8531] = 256'he70584053405e604b004ab040505dd05f8060508b608b508f407b70654053304;
    inBuf[8532] = 256'haf03d1036c043505c305e905c5058b0590051306e2069d07e2075c071d06a904;
    inBuf[8533] = 256'h93034c03f70332056b06240715076e06af0537053d05c0055f06bd06c4067d06;
    inBuf[8534] = 256'h26060f064306a006e306b60605060b052104c2034d04a8056a070c09e6099d09;
    inBuf[8535] = 256'h55087906a90477031b0380035e044505fe058c06ed062f0759073b07b506db05;
    inBuf[8536] = 256'hd404e803610350039a0316048504d7041d0554058505b505c405b105a905c305;
    inBuf[8537] = 256'h1206920606072207bd06d605ae04b203310365035204a705fe0600085408dd07;
    inBuf[8538] = 256'hcf06770538047203340357039803b303a803bc0334044105bf061a08ab082108;
    inBuf[8539] = 256'h89067404b802eb012902160308047f046304ef039d03d1038604760542068d06;
    inBuf[8540] = 256'h3d067e0586049303db0275026902b9024803f0038a04f0042505450559055d05;
    inBuf[8541] = 256'h3c05c204df03c702d3016801c601d00226044f05e805df056d05db0464041e04;
    inBuf[8542] = 256'he8039d033503b9024a020b02fb01010207020202fd0113025002b60232039b03;
    inBuf[8543] = 256'hd303d50399031f036f028f019800b9ff2cff25ffbcffd1001b024203f9032804;
    inBuf[8544] = 256'hea0377030f03d502bc0294022a025f0143001bff47fe23fed8fe48001102ad03;
    inBuf[8545] = 256'ha004aa04e1039f025d018000300052009d00be008000deff02ff2efea4fd93fd;
    inBuf[8546] = 256'h05fed9fed5ffb7004901770151010101b0006b001c00a3ffedfefffd0afd48fc;
    inBuf[8547] = 256'he1fbdafb17fc7afc05fdd3fdfdfe82001d024d039203a402a60026fee5fb84fa;
    inBuf[8548] = 256'h54fa2bfb83fcc4fd7afe78fef4fd53fd00fd57fd69fefaff9b01c202ee02e501;
    inBuf[8549] = 256'hbfffe0fcebf97df707f6cef5cdf6bbf83ffbe0fd12006901a301ba000cff21fd;
    inBuf[8550] = 256'h83fb8ffa45fa47fa2cfaaaf9c3f8e7f7a2f759f82cfac1fc5aff4101ee013001;
    inBuf[8551] = 256'h52ffe3fc83fac3f8e1f7d1f76af866f97ffa9ffbb9fcaafd56fe8ffe24fe1ffd;
    inBuf[8552] = 256'hb2fb2bfaeff83cf810f851f8c4f833f9a6f92efacefa94fb60fce6fcfbfc89fc;
    inBuf[8553] = 256'h96fb60fa2cf930f897f75bf74ff759f759f740f744f7a4f787f807faf6fbd5fd;
    inBuf[8554] = 256'h22ff6dff7cfe8bfc15faa9f7d2f5cff48ff4f7f4d1f5e9f645f8dbf97bfbf7fc;
    inBuf[8555] = 256'h0efe77fe26fe32fdcffb54fa04f905f881f775f7b4f71df871f868f803f86bf7;
    inBuf[8556] = 256'he3f6d9f690f7f0f8acfa3efc17fdfcfcedfb25fa28f861f60ff574f49ff46bf5;
    inBuf[8557] = 256'hb6f63ef89cf987facffa65fa88f985f89bf710f7f5f62bf7aef768f833f90bfa;
    inBuf[8558] = 256'hd7fa60fb93fb67fbd7fa12fa40f96bf8a7f7edf62df698f564f5bdf5daf6a9f8;
    inBuf[8559] = 256'hc0faa7fcdffd04fe21fd85fba0f902f800f79df6c1f61ff758f751f70bf79df6;
    inBuf[8560] = 256'h59f67ff61df735f892f9cdfa9bfbc3fb2efb17fad2f8acf701f7f3f65df71df8;
    inBuf[8561] = 256'hf2f88af9cef9b1f934f989f8e9f77ff78ff733f84af9a8faf9fbd5fc16fdbbfc;
    inBuf[8562] = 256'he4fbebfa17fa7ff92ff908f9d2f880f815f89cf750f760f7ddf7ddf849fadafb;
    inBuf[8563] = 256'h4afd43fe73fec5fd4cfc3afafcf7faf582f4e1f332f456f521f741f947fbe2fc;
    inBuf[8564] = 256'hd4fdf9fd6dfd61fc11fbd2f9e3f861f867f8e7f8a9f985fa48fbc2fbf7fbfbfb;
    inBuf[8565] = 256'he1fbcdfbd2fbe6fb07fc23fc1ffcfefbb7fb41fbb9fa43fafbf917fab3fab6fb;
    inBuf[8566] = 256'hf5fc23fee6fe0eff8ffe83fd35fce8faccf90cf9b2f8aef803f9a7f97ffa75fb;
    inBuf[8567] = 256'h6afc36fdc7fd1afe38fe37fe1cfed7fd61fda6fca7fb94faaff932f959f931fa;
    inBuf[8568] = 256'h89fb19fd88fe87fff6ffe0ff74fff9fe9cfe66fe46fe0cfe89fdc5fcf0fb58fb;
    inBuf[8569] = 256'h56fb1bfc8ffd59fffa00fa0117025301f5ff6afe0efd1bfca8fb9ffbdbfb45fc;
    inBuf[8570] = 256'hcdfc68fd11fec4fe75ff17009600df00d900690088ff4ffef2fcbefb0afb14fb;
    inBuf[8571] = 256'heafb6cfd53ff3b01be0291039103ca027e011500f8fe6afe77feeefe73ffb8ff;
    inBuf[8572] = 256'ha0ff50ff17ff41fff2ff150156025a03e303dd035f039b02bc01dd00120067ff;
    inBuf[8573] = 256'he9feabfeb3fefbfe73ff03009a003601cd015202b902e302ba0247029c01d800;
    inBuf[8574] = 256'h22008eff29ff04ff2bffb3ffa900ee013b034204ab04560470034e025d01f500;
    inBuf[8575] = 256'h1f01ac015802d9020a030003da02bb02c102e1020e034b038f03dc033e04a104;
    inBuf[8576] = 256'hea040805e4047904e5033d03a402430222023d028b02e5022b03570359034003;
    inBuf[8577] = 256'h3103360357039d03f0033b047c04a504b804c804cb04bb0499044704b503f702;
    inBuf[8578] = 256'h1f026101100159014e02de03a9053e074b08940824084c075b06990537051705;
    inBuf[8579] = 256'h10050705da048c044d0437046004d8047e0522069f06bd066d06da053405c504;
    inBuf[8580] = 256'hd9046a05450620078f075c07ad06bd05e50478047404aa04e704f004c3049404;
    inBuf[8581] = 256'h8604bc044505ee058a060f077407cf074908d608500989093309260888069a04;
    inBuf[8582] = 256'hd702cf01d201f20202056a0790090b0b960b4d0b9f0ae8096b093a090b098c08;
    inBuf[8583] = 256'h9407180666040b036d02ce022f0424062508bb09790a410a5009ef0783067605;
    inBuf[8584] = 256'hf004f3046b051206b5064307a607e90731086b08840870080708440752065605;
    inBuf[8585] = 256'h8b0432045404e904e60514074e088809980a6f0b060c2f0ccf0bee0a8709be07;
    inBuf[8586] = 256'he505400411039202c3029403eb0488063b08e309420b2a0c850c290c0f0b6209;
    inBuf[8587] = 256'h490715053403ee017a01e90102037404ec051307d10749089308d30821095009;
    inBuf[8588] = 256'h2d09a208a60765062e053a04b403ab03f8037e043205f805cb06ab077008f808;
    inBuf[8589] = 256'h330906097508a307a7069e05b004f10383038203e7039f048a055d06e9062d07;
    inBuf[8590] = 256'h2a07ff06d706ae066e06fa053205270416033e02e50135020a032c0455053406;
    inBuf[8591] = 256'ha0069e0632067905a104c40303037f0242025302ab022b03c2036704fa046e05;
    inBuf[8592] = 256'hba05bf057305e8043a049a033603180331035c036a0350032803110333039503;
    inBuf[8593] = 256'h06044c043b04be03f7022d029a0164018a01e4014c02a502da02f002f002cf02;
    inBuf[8594] = 256'h8d022f02bd0153010e01f000f5000301fb00d900af009800b4000d018201ea01;
    inBuf[8595] = 256'h1502e2015c01a600eeff65ff2dff52ffdaffbb00ce01e602be030f04b803c402;
    inBuf[8596] = 256'h6801feffd8fe22fee3fdfbfd44feb3fe4bff12000a011302ed025b0334037602;
    inBuf[8597] = 256'h4a01ebff99fe8afdddfca0fcdbfc80fd72fe85ff7c0016012e01ba00d4ffb9fe;
    inBuf[8598] = 256'hacfdeefca2fccafc4ffd0bfec8fe5dffbaffd7ffb8ff78ff2affdefe9afe5afe;
    inBuf[8599] = 256'h15fec5fd65fd05fdc2fcaefce3fc6bfd33fe1dff0900c90038013f01ce00eaff;
    inBuf[8600] = 256'ha9fe35fdd2fbc2fa31fa3cfad7fac1fbbbfc93fd22fe69fe83fe88fe81fe6bfe;
    inBuf[8601] = 256'h2cfebdfd26fd80fcfcfbbcfbbdfbebfb21fc30fc17fcfdfb0dfc72fc36fd28fe;
    inBuf[8602] = 256'hf8fe53fffefe04fea8fc4dfb66fa44fae8fa27fcaafdf4feabffa4ffe8febafd;
    inBuf[8603] = 256'h79fc79fbf3faeafa2cfb89fbd3fbf3fb00fc21fc63fccdfc4efdbafdf4fdf3fd;
    inBuf[8604] = 256'hb5fd4efdcefc3bfca3fb0dfb77faf6f99bf965f968f9b4f946fa1bfb24fc31fd;
    inBuf[8605] = 256'h15fea8fecffe99fe1dfe70fdaffce2fb06fb35fa94f944f970f921fa30fb66fc;
    inBuf[8606] = 256'h80fd3cfe82fe56feccfd19fd69fcdbfb90fb89fba4fbc6fbcffbacfb7bfb6ffb;
    inBuf[8607] = 256'hadfb4ffc34fd09fe7afe47fe61fd0ffcb3faaaf93ff979f925fa0efb00fcd7fc;
    inBuf[8608] = 256'h98fd43fec3fe02ffd8fe24fefafc8ffb2afa29f9c4f8fef8c3f9d8faf2fbebfc;
    inBuf[8609] = 256'habfd25fe71fe9dfea7fe94fe50fec1fdebfcdffbc5fae6f97cf99ef94afa45fb;
    inBuf[8610] = 256'h3afcf8fc65fd88fd95fdb5fde9fd1ffe1ffebafdf5fcf6fbfffa6bfa69faeffa;
    inBuf[8611] = 256'hd7fbd0fc87fdd9fdbefd45fda8fc18fcacfb7cfb85fbb4fb01fc5afcaffc04fd;
    inBuf[8612] = 256'h50fd84fda2fd9dfd6afd1cfdc6fc7bfc5cfc73fca9fce6fc04fde8fca1fc4dfc;
    inBuf[8613] = 256'h18fc38fcb4fc70fd43feeafe2cff00ff75feaffdeefc63fc23fc33fc74fcbcfc;
    inBuf[8614] = 256'hf0fcf4fcc1fc76fc2bfcf1fbe1fbfefb41fcaefc37fdc9fd5dfed1fefdfed3fe;
    inBuf[8615] = 256'h4cfe7afd89fca2fbeffa98faa2fa05fbbafb9ffc7dfd2dfe82fe6efe0bfe8afd;
    inBuf[8616] = 256'h24fd0dfd3efd8bfdc6fdbbfd62fdebfc8ffc7afcc2fc41fdbefd0afe07febbfd;
    inBuf[8617] = 256'h51fdedfcb0fcb4fcf2fc56fdd0fd34fe61fe50fe00fe87fd16fdccfcb5fcd1fc;
    inBuf[8618] = 256'h05fd38fd66fd8dfdadfdcbfdd6fdc0fd8dfd43fdfefce4fcfcfc36fd82fdc7fd;
    inBuf[8619] = 256'hf3fd13fe35fe66fea5fed4fed5fe9bfe1bfe6bfdbafc2dfcdffbebfb4afce9fc;
    inBuf[8620] = 256'hb6fd8bfe42ffc5fffcffe1ff7effdffe1cfe54fd9dfc14fcd9fbeffb4bfcdffc;
    inBuf[8621] = 256'h88fd28feb2fe21ff72ffa2ff9aff47ffa4fec2fdd4fc24fcdffb15fcb6fc85fd;
    inBuf[8622] = 256'h4cfef1fe6dffc8ff0f0035002800d5ff35ff66fe94fde2fc6ffc4ffc7bfce9fc;
    inBuf[8623] = 256'h94fd6afe4eff1b00a600dc00be005900d1ff46ffbffe3ffed1fd7cfd57fd73fd;
    inBuf[8624] = 256'hc5fd35fea0fee8fe0eff2fff6fffe2ff7500ee001201bd00f2fff0fe0bfe7dfd;
    inBuf[8625] = 256'h5cfd9bfd09fe79fed9fe2aff77ffc6ff070022000700acff2cffb1fe5ffe53fe;
    inBuf[8626] = 256'h95fe0bff93ff0f005c00710057001f00e0ffadff87ff64ff3afffdfeb6fe82fe;
    inBuf[8627] = 256'h7afeb6fe38ffe7ff9a002b017a01820157011001c900950071004f002400e3ff;
    inBuf[8628] = 256'h8fff35ffebfec7fedafe26ffa4ff4900fe00b1014902ac02c3027e02d701e500;
    inBuf[8629] = 256'hd5ffe3fe4dfe3cfeb6fe97ff9d00820118024f023602ec018f012901b9003b00;
    inBuf[8630] = 256'hbcff5cff44ff92ff4e005c0181027d0313041f04a203b002740129000eff58fe;
    inBuf[8631] = 256'h24fe70fe28ff2700380138021403bc031e043004e703420353023e01370072ff;
    inBuf[8632] = 256'h13ff2bffaeff750057012a02c3020e031103da027f021d02c801880162015b01;
    inBuf[8633] = 256'h7801ba011b028a02ee0223031703d60273021002d601d50100023b0263026602;
    inBuf[8634] = 256'h45021102ec01f30130029e022903b00310043004fc037b03ca020e0272011501;
    inBuf[8635] = 256'h000129017901da014602bf023d03b6031404360406048e03ee025a020102f701;
    inBuf[8636] = 256'h3b02ae0227038503b1039f035303d9024202ae0148012c016901fc01c0028603;
    inBuf[8637] = 256'h1c0463045f042204c50369031e03e302bb02a802a902c202f102220344034303;
    inBuf[8638] = 256'h1503c80277023f023a027102d5025903e5036204c8040c051805e1046704ae03;
    inBuf[8639] = 256'hd302050272013f017401f901a9025903df0333045e04680463045a0440041304;
    inBuf[8640] = 256'hd1037203020395023402f201de01f9014602c1025103e5036904c104de04be04;
    inBuf[8641] = 256'h5e04d2033703a70241021a0223024b027b029d02b402dc022f03c2038e045e05;
    inBuf[8642] = 256'hf1050a067e056004f40291018f002b0062000e01f201cd027e0305046704b104;
    inBuf[8643] = 256'he604eb04ac042d048103d60263023d025c029d02cc02cb02a102680251027f02;
    inBuf[8644] = 256'heb02790300044c044a040a04a5033f03fb02e202f1021c034b036f0383038203;
    inBuf[8645] = 256'h7b0377036e035d033a03f00285021802c801b90101028d023403c1030604ff03;
    inBuf[8646] = 256'hc80383035403490343032303d1024702a4011701c000b600ff0084012e02e802;
    inBuf[8647] = 256'h98032e049a04c304a5044c04c30324038b020002930149011d01130130016501;
    inBuf[8648] = 256'hab01fd015102aa020b036803b903f5030304d8037603df022d028201f700af00;
    inBuf[8649] = 256'hc3002701c1016b02ef022d031c03c8025702f301ae019201a001c501fa013e02;
    inBuf[8650] = 256'h8402c302f302fe02d902850202026701d500630030005c00df009f0178022f03;
    inBuf[8651] = 256'h950399034003af02180294012b01d9008e004d002b004000a100490105029802;
    inBuf[8652] = 256'hd5029f02060244019b003a0033007500dd0049019801c401d501d001bf01a801;
    inBuf[8653] = 256'h860158012301de008b003500e6ffaaff94ffb2ff0c0099004501fc019f020703;
    inBuf[8654] = 256'h1703c2020402f300c4ffb1fef6fdbafd00feb2fea3ff9c007401150274029202;
    inBuf[8655] = 256'h79022d02b80127018100d1ff29ff96fe2afef8fd14fe88fe49ff35002401e501;
    inBuf[8656] = 256'h48023d02d1011e014b0089fff4fe9afe76fe79fe92feb4fed8fe0dff5fffcdff;
    inBuf[8657] = 256'h4f00d10028013001dd0032004dff59fe86fdfbfccdfc02fd95fd6dfe63ff5500;
    inBuf[8658] = 256'h2501b301e801b9011e011f00dafe81fd56fca1fb8afb1afc2ffd88fed7ffe000;
    inBuf[8659] = 256'h8001b0017901eb00160013fffefdfdfc3dfce2fbfcfb81fc54fd47fe25ffc2ff;
    inBuf[8660] = 256'h0300e9ff8dff11ffa0fe5afe3ffe3afe2efe05feb9fd5dfd19fd0cfd45fdb4fd;
    inBuf[8661] = 256'h38fea7fee5feebfec7fe8dfe4ffe19feeafdbafd88fd5afd33fd23fd32fd61fd;
    inBuf[8662] = 256'ha9fdfefd4efe8cfeacfea4fe77fe2bfec3fd50fde2fc83fc44fc31fc54fcb3fc;
    inBuf[8663] = 256'h3efdd4fd57fea8feacfe68fef2fd67fde6fc86fc51fc4efc7cfcc8fc26fd83fd;
    inBuf[8664] = 256'hc4fddefdd2fda7fd79fd5dfd56fd64fd7dfd89fd87fd78fd57fd2efd08fdeafc;
    inBuf[8665] = 256'hdafcdffcf9fc24fd4cfd5afd52fd3bfd20fd19fd3bfd77fdb7fde0fdd2fd89fd;
    inBuf[8666] = 256'h18fd97fc2bfcf3fbf8fb39fca4fc19fd82fdccfde4fdd3fdb0fd8afd75fd75fd;
    inBuf[8667] = 256'h75fd60fd22fdb3fc2efcbcfb83fb9ffb0bfca4fc47fdcefd1bfe2ffe1cfeeefd;
    inBuf[8668] = 256'hb9fd8dfd6cfd58fd42fd13fdc9fc63fceffb96fb80fbb9fb3ffcebfc81fddcfd;
    inBuf[8669] = 256'hebfdb8fd6cfd2efd14fd29fd57fd83fda4fdb0fd98fd66fd23fdcdfc72fc25fc;
    inBuf[8670] = 256'hf2fbeefb1bfc6dfcdefc5bfdcbfd2afe64fe63fe2afec2fd3efdccfc91fc97fc;
    inBuf[8671] = 256'hd9fc32fd69fd67fd29fdc1fc63fc36fc49fc9afc0afd76fdd2fd17fe3afe4cfe;
    inBuf[8672] = 256'h54fe44fe1bfedafd76fd00fd8cfc2cfc05fc22fc6ffcd6fc33fd5efd56fd30fd;
    inBuf[8673] = 256'h09fd0efd50fdb8fd2ffe8efeadfe8cfe39fec4fd4dfde6fc8bfc44fc15fcf5fb;
    inBuf[8674] = 256'heefb0bfc4dfcbdfc55fdfbfd99fe13ff46ff30ffdafe51feb8fd2bfdb3fc61fc;
    inBuf[8675] = 256'h39fc2ffc45fc79fcc3fc1cfd79fdc8fd0afe42fe77febafe09ff4aff63ff35ff;
    inBuf[8676] = 256'haafed5fde3fc08fc79fb55fb91fb1dfcd3fc8bfd34febefe18ff40ff34fff3fe;
    inBuf[8677] = 256'h96fe2bfebcfd5bfd0efdd7fcc2fcd5fc0efd6afdd3fd24fe4ffe4afe19fedafd;
    inBuf[8678] = 256'haffdadfde2fd3cfe99feddfee8feabfe3dfebcfd45fdfffcf6fc1ffd67fdb6fd;
    inBuf[8679] = 256'hf8fd32fe68fe9cfed2fef8fef4febffe59fedafd72fd44fd5bfdb6fd2efe8dfe;
    inBuf[8680] = 256'hb4fe9bfe4efef8fdbdfdb0fdd8fd1afe4efe61fe4afe15feebfdedfd29fe9dfe;
    inBuf[8681] = 256'h26ff95ffcbffbdff73ff14ffbffe81fe56fe2efef4fdaafd5ffd2cfd37fd90fd;
    inBuf[8682] = 256'h2bfef0feb8ff5300a2009b004800ccff48ffd0fe70fe25fedefd9efd71fd6bfd;
    inBuf[8683] = 256'ha2fd1afebefe6dff00005c00790060002400d8ff84ff2dffd9fe8dfe4bfe18fe;
    inBuf[8684] = 256'hfffd05fe2ffe7ffef1fe73ffedff4800710064002f00e2ff8bff3bfffffed6fe;
    inBuf[8685] = 256'hc4fed4fe0cff69ffd8ff3f00870098006a000e009eff2fffdbfeb0feb2fee1fe;
    inBuf[8686] = 256'h3affadff29009800e3000001ec00b10066002000e2ffb0ff8aff6eff63ff74ff;
    inBuf[8687] = 256'ha4fff2ff5000a900f300220130012101f500ac005200f8ffadff86ff8affb9ff;
    inBuf[8688] = 256'h0a006800bf0008013a01500150013c011701ee00c700a50091008c009200a500;
    inBuf[8689] = 256'hc600ed00170136014501430132011a010c010d011a013701590172017b016d01;
    inBuf[8690] = 256'h4a011d01f100d000cb00e5001a015f019f01cb01df01d501ba01a5019b019d01;
    inBuf[8691] = 256'ha601a901a401a001a301b201d501f601fd01e0019f0151011b0113014301a801;
    inBuf[8692] = 256'h20028e02e90225033e033b031303c4025d02e6017901370129014e01a1010902;
    inBuf[8693] = 256'h7402dd0233036f038b0370031b03a0020e02850130011c014501a20113028202;
    inBuf[8694] = 256'hea0242038903c803ef03f303d503890313038e020502920158016201b1014102;
    inBuf[8695] = 256'he7027803da03f703d903a80378035b03580355033c031203de02b602b502d602;
    inBuf[8696] = 256'h070334033a031203d902a902a102dd024d03cc03340455041c04a6031b03ae02;
    inBuf[8697] = 256'h9102c5023503b90312041d04e5037b030303ae0289028a02a702c502e1020a03;
    inBuf[8698] = 256'h4d03b8035004f5048205d305c20546057704710364028701fa00d7002f01e901;
    inBuf[8699] = 256'he302f703ea049205e205d2057305e4043a0492030903a4026702570267029002;
    inBuf[8700] = 256'hd7022d038f03fd0359048e04960468041104b203610335033c0361039603d403;
    inBuf[8701] = 256'h030419041604e6038f032b03cb028e029702e2025b03e203420460044004ec03;
    inBuf[8702] = 256'h8d0358035e039c03fd03470455041d049e030103880255027902e5025f03b703;
    inBuf[8703] = 256'hdb03c5039103710377039b03cb03e203d603b303850361035a0357033c030703;
    inBuf[8704] = 256'hb702680245025f02b10228039403d103d903b00370033f032a03330352036803;
    inBuf[8705] = 256'h5a032303c2025002fc01db01f8015202c6022a036b037e037203640364037a03;
    inBuf[8706] = 256'ha003b4039d035803e7025b02d9017d0158017301bd0121028a02dd020c031e03;
    inBuf[8707] = 256'h16030003ed02dd02d102c802b20288024c02fb01a4015b012b01250150019c01;
    inBuf[8708] = 256'hf1013c026702700268025d0261027b029902a4028a024702ef019e0166015401;
    inBuf[8709] = 256'h60016d0169015901470146016601a001e1011a023e0251025e0266026a025c02;
    inBuf[8710] = 256'h2602ca015901e10075002900fdfff0ff0a004e00c0005201e40155028c027902;
    inBuf[8711] = 256'h2702b5013801bf0058000a00ddffdaff02005000b10006013d0154014b013001;
    inBuf[8712] = 256'h1201f300cd00a40080006b006e008800ab00c300c300ad0090007a0077008700;
    inBuf[8713] = 256'h9b00a200900062001d00d6ff9fff84ff8fffc2ff10006500ac00d500d200a300;
    inBuf[8714] = 256'h5a000d00c8ff91ff6dff5eff5dff66ff7cff97ffa8ffa8ff99ff85ff80ff94ff;
    inBuf[8715] = 256'hc6ff0a00450057003700e9ff82ff24ffe9fedafef4fe28ff62ff98ffbfffd0ff;
    inBuf[8716] = 256'hcfffbcff95ff64ff33ff05ffe6fedafedcfef0fe13ff37ff59ff77ff89ff8bff;
    inBuf[8717] = 256'h7bff5aff32ff02ffc6fe82fe3bfef5fdc6fdc1fdebfd47fec2fe38ff92ffc2ff;
    inBuf[8718] = 256'hbbff83ff2cffc1fe51fee8fd90fd59fd4bfd60fd9bfdf3fd4ffea5feedfe17ff;
    inBuf[8719] = 256'h21ff11ffedfec3fe9dfe79fe5cfe3ffe15fee5fdb9fd97fd89fd93fda8fdc8fd;
    inBuf[8720] = 256'hf0fd1bfe4dfe83feabfeb7fe9dfe57fef6fd94fd41fd10fd05fd14fd38fd67fd;
    inBuf[8721] = 256'h95fdc0fdddfdddfdc0fd88fd3cfdf9fcd3fccdfceefc29fd65fd98fdc0fdd7fd;
    inBuf[8722] = 256'he4fdeefdedfddffdb5fd64fdf8fc7afcfefbabfb9ffbddfb65fc1cfdd3fd6afe;
    inBuf[8723] = 256'hc4fed0fea1fe4afeddfd6ffd07fd9efc3cfcddfb84fb4cfb46fb71fbd8fb6cfc;
    inBuf[8724] = 256'h07fd8efde3fdeffdc3fd73fd0efdb2fc69fc27fceefbc1fb9efb97fbb4fbe7fb;
    inBuf[8725] = 256'h28fc5dfc67fc4dfc1ffcf3fbeefb21fc71fccafc0dfd1cfdfefcc7fc82fc4bfc;
    inBuf[8726] = 256'h29fc12fc0cfc18fc27fc39fc40fc25fcf2fbb8fb8afb8dfbcdfb2efc92fcd8fc;
    inBuf[8727] = 256'he0fcb7fc7cfc41fc1ffc17fc13fc0afcf2fbbcfb74fb1ffbbdfa6dfa4dfa69fa;
    inBuf[8728] = 256'hd1fa7bfb38fcddfc42fd4afd0afda5fc32fcd3fb92fb5efb30fbfdfabdfa85fa;
    inBuf[8729] = 256'h69fa73fab8fa3cfbe4fb95fc2afd79fd7dfd3cfdc3fc41fcd3fb82fb58fb4bfb;
    inBuf[8730] = 256'h41fb36fb23fb09fb00fb15fb45fb9afb03fc63fca8fcc4fcaafc69fc16fcc3fb;
    inBuf[8731] = 256'h8cfb75fb6ffb6ffb65fb40fb0efbdcfabdfacdfa09fb57fbb1fb06fc44fc76fc;
    inBuf[8732] = 256'h9ffcb4fcb5fc95fc49fce5fb7bfb1cfbeafaeefa17fb64fbc5fb20fc70fca9fc;
    inBuf[8733] = 256'hc0fcc7fcc5fcbffccafcddfcdbfcb8fc6cfcfdfb95fb5afb5bfb9ffb0afc6bfc;
    inBuf[8734] = 256'haafcb9fc9dfc76fc55fc43fc4bfc65fc7afc8bfc91fc82fc69fc4afc28fc12fc;
    inBuf[8735] = 256'h11fc1bfc32fc4ffc68fc83fc9bfcacfcbcfcc2fcb7fca7fc9dfc9cfcb5fce6fc;
    inBuf[8736] = 256'h20fd61fd9efdcbfdebfdf6fde0fda7fd4ffde4fc8efc6ffc94fcfbfc83fdfcfd;
    inBuf[8737] = 256'h45fe50fe25feebfdc4fdbefddcfd09fe26fe1efee6fd89fd23fdcffca3fcb3fc;
    inBuf[8738] = 256'hf8fc5afdc5fd1bfe47fe4ffe3efe25fe16fe1afe2afe40fe4dfe49fe39fe20fe;
    inBuf[8739] = 256'h08fefbfdfbfd03fe12fe2afe56fea3fe0aff78ffd9ff0a00fcffbfff6dff25ff;
    inBuf[8740] = 256'h00fffbfe02ff02ffecfec7feadfeb2fee8fe52ffd5ff5200af00d100a8004100;
    inBuf[8741] = 256'hb2ff17ff98fe4cfe3afe61feb3fe1eff96ff0c007200bc00da00cb009b005400;
    inBuf[8742] = 256'h0000aeff62ff2cff24ff51ffb3ff3600b30009012a011a01f700e700f8002901;
    inBuf[8743] = 256'h66019001970178013b01f800c600ac00af00d100010133015b0175018d01b101;
    inBuf[8744] = 256'hea013b028f02bf02b0025802bb01040169001500250090003101db016002a202;
    inBuf[8745] = 256'ha8028a026402480236021e02f501b4016601300127015601bb013a02b4021b03;
    inBuf[8746] = 256'h64038c039a038f036b033203e5028e0248021c0219025202bf024c03e7036b04;
    inBuf[8747] = 256'hb304b5046f04f80378030c03cd02d10204034c039a03cc03d103b80388035403;
    inBuf[8748] = 256'h3f0350038003cb0314043b043d041404c703770336030b030603230353039303;
    inBuf[8749] = 256'hd4030b043904510455045704590467049004c204ea0406050605e304ae047104;
    inBuf[8750] = 256'h36041404100436048d04fb046405bb05e405dc05bd05980574055d0541050e05;
    inBuf[8751] = 256'hcf0488044604210416041e043a045f048e04d6042e058805dd050e060606c505;
    inBuf[8752] = 256'h4805a104fc0379033c036203da037d042705a705e605f305dd05bb05ab05a705;
    inBuf[8753] = 256'ha405a20591056a053c050c05ea04f4042905870505067906c406dc06b0064a06;
    inBuf[8754] = 256'hca054005cb048d048604b6041d059205f5054006600652062606d6056805f204;
    inBuf[8755] = 256'h7d042204060421046204b804fd0422053a05470557057c059d05ab05af059705;
    inBuf[8756] = 256'h63052905e0048d04570448046d04cf044805b005f405ff05d705a6057d056c05;
    inBuf[8757] = 256'h8105a205c005dc05e205cc05aa0573052a05e10497045a04400445046c04bd04;
    inBuf[8758] = 256'h160563059805980564051b05c604760440041204e103b4037e034f0345036103;
    inBuf[8759] = 256'ha7031e04a60422057f0597056005f1045a04bf034d03100312035503bb032d04;
    inBuf[8760] = 256'h9d04ec0413051f050b05df04ac0468041a04d4039b0380039403c203f6032104;
    inBuf[8761] = 256'h2a041304f303d703d303e903f403d9039203180388021902eb0114028d022603;
    inBuf[8762] = 256'hb3030504f9039a030f037602ff01cd01d6010b02530287029702890268025802;
    inBuf[8763] = 256'h7402b102fd023c0340030603a9024702070201022302570287029e02a2029e02;
    inBuf[8764] = 256'h90027e0270025b02400224020102db01bd01a5019d01b101d101eb01f301d601;
    inBuf[8765] = 256'h96014a010401d800cf00d900e800f200ec00d300b0008600670063007a00a900;
    inBuf[8766] = 256'hd900e800cc009100470012000f00330069009b00b000a7009000780069006e00;
    inBuf[8767] = 256'h81009800a700a100890066003f0028002e0044005a005a003800fdffc0ff92ff;
    inBuf[8768] = 256'h86ff94ffa4ffa0ff84ff58ff2bff0afffbfefefe08ff0cff08fff3fec6fe8cfe;
    inBuf[8769] = 256'h51fe29fe25fe48fe7efeb0fec9febefe9dfe77fe5bfe4efe46fe3efe35fe2bfe;
    inBuf[8770] = 256'h2bfe42fe65fe88fea2fea8fe9afe82fe66fe50fe49fe48fe49fe47fe32fe09fe;
    inBuf[8771] = 256'hdcfdaffd8efd8afd9cfdb8fdd7fdeafdebfdd6fda8fd65fd16fdbbfc6cfc41fc;
    inBuf[8772] = 256'h40fc6efcbffc0efd43fd53fd32fdeffca5fc60fc2ffc15fc02fcf3fbecfbe9fb;
    inBuf[8773] = 256'hfefb35fc86fce1fc2afd40fd22fddafc77fc20fcedfbd6fbd8fbe9fbf2fbf7fb;
    inBuf[8774] = 256'h03fc14fc39fc73fca9fcccfccdfc9afc47fcebfb94fb60fb57fb64fb81fb9dfb;
    inBuf[8775] = 256'h9ffb8ffb79fb5dfb4dfb52fb61fb76fb81fb6ffb49fb12fbccfa97fa7ffa77fa;
    inBuf[8776] = 256'h84faa1fabdfae1fa0afb24fb30fb26fbf8fabffa93fa74fa72fa89faa0fab7fa;
    inBuf[8777] = 256'hcbfad6fae3faf0faeffaf2faf6faedfae9fae8fad8fac4fab6faa7faa4faabfa;
    inBuf[8778] = 256'habfaabfaa5fa96fa9afaabfaaafa9cfa7ffa46fa14fa02fa09fa27fa47fa45fa;
    inBuf[8779] = 256'h29fa01fad1f9b7f9bcf9c7f9d7f9e6f9e5f9e2f9e7f9eaf9fbf919fa35fa4ffa;
    inBuf[8780] = 256'h58fa3afa04fac8f996f991f9c1f90bfa5ffaa1fab5faaffa9efa86fa7ffa85fa;
    inBuf[8781] = 256'h7efa6dfa51fa1cfae7f9c6f9bcf9dcf922fa6bfaacfacefabbfa88fa4ffa18fa;
    inBuf[8782] = 256'hfdf9fdf901fa07fa02fae6f9cef9c1f9b6f9c0f9e3f909fa35fa5efa64fa4efa;
    inBuf[8783] = 256'h27faf6f9dbf9e1f9f8f91cfa3dfa4afa52fa5bfa62fa79fa97faa6fab8facafa;
    inBuf[8784] = 256'hc9fac0fab6faa0fa90fa8bfa8efaa8facafadbfae7faf2faf8fa0efb33fb4afb;
    inBuf[8785] = 256'h4efb30fbebfaa3fa76fa6bfa90facffa07fb32fb42fb2ffb19fb0bfbfcfafbfa;
    inBuf[8786] = 256'h02fb00fb01fb03fbfdfa00fb0cfb16fb2cfb47fb58fb6afb76fb70fb70fb7cfb;
    inBuf[8787] = 256'h88fb9efbaefba6fb96fb8dfb8ffbb3fbf5fb3afc71fc8bfc7efc5efc38fc13fc;
    inBuf[8788] = 256'h02fc08fc1afc37fc57fc71fc87fc8ffc8cfc92fc9dfca4fcacfcaafc91fc75fc;
    inBuf[8789] = 256'h61fc55fc5ffc79fc96fcb4fccbfcd6fcdffce0fcd7fccffccffcd7fceefc0efd;
    inBuf[8790] = 256'h2bfd3ffd45fd41fd42fd4cfd5efd7bfd98fda9fdb1fdacfd9bfd8dfd94fdb4fd;
    inBuf[8791] = 256'hf0fd38fe71fe86fe6bfe2efef7fde5fd01fe45fe8ffebffec3fea1fe73fe56fe;
    inBuf[8792] = 256'h55fe72fea2fecffeedfef7feeafeccfeabfe96fe95feadfed6fe03ff26ff38ff;
    inBuf[8793] = 256'h3eff44ff4aff4fff4cff3aff21ff0fff15ff3dff82ffd0ff1100340033001b00;
    inBuf[8794] = 256'hf8ffd5ffc2ffc5ffdafffcff22004300610081009f00bd00d900eb00e900d600;
    inBuf[8795] = 256'hbd00ac00a900b800d500f3000701110116011d012e0143015801690170017101;
    inBuf[8796] = 256'h75017c0185019201940187017901700170018401a501c701eb01050213022002;
    inBuf[8797] = 256'h2c0238024e02660271026c02520227020102f60115026702d10230036e037603;
    inBuf[8798] = 256'h510322030003f80210032e033f03430335032103210337036203a703e9031004;
    inBuf[8799] = 256'h1c04ff03c00383035c0357037c03b203e003fe03050400040704130421043504;
    inBuf[8800] = 256'h370422040f04fd03f6030b04300459048f04b804cf04e104e404d904d604d104;
    inBuf[8801] = 256'hc104b504a50493049704af04db041e0558057f059d05a305960590057c054f05;
    inBuf[8802] = 256'h2405fa04d804de0409054c05a305ee051a062d061806e405b10581055c055805;
    inBuf[8803] = 256'h640576059605b105c405e105f705050612061006030601060106040617061d06;
    inBuf[8804] = 256'h0d06f705cf05a4059b05ab05d10511064d0678069c06a806a2069d068a066d06;
    inBuf[8805] = 256'h5a063d061606fd05ee05ee05120647067d06b106c806bc06a6068b067b068a06;
    inBuf[8806] = 256'ha106b006b106880641060206d805d70512066906c00605071007e1069e065306;
    inBuf[8807] = 256'h18061006280646065d064f062006f505dd05e70520066c06ae06db06d706ac06;
    inBuf[8808] = 256'h760638060606f805fe050d062c06410646064c064a064506520660066e067f06;
    inBuf[8809] = 256'h7b06600644061d06f105d905c805bc05c505d405e405ff05120617061b061306;
    inBuf[8810] = 256'hfe05ed05d305af05930573055205450541054a056e059605b405ce05d105b605;
    inBuf[8811] = 256'h8c05570524050905ff040705260541054e0556054c053505270519050a050505;
    inBuf[8812] = 256'hfb04ec04e604db04ce04cb04c004b704c004ca04ce04d804d204bb04a4048604;
    inBuf[8813] = 256'h630449042d0413040b040c0416042f043f04400440043a04310429041204ea03;
    inBuf[8814] = 256'hba038303540342034303540375039403ad03c003bf03a80389035e0333031603;
    inBuf[8815] = 256'hff02ef02e102cc02be02c802e002040330034b0348032f03fd02c00288025802;
    inBuf[8816] = 256'h37022c022f023c0249025002590264026c0273027602650245021b02eb01c101;
    inBuf[8817] = 256'ha2018001640151014401470161018401a701c001bf01a5017c014a011901f000;
    inBuf[8818] = 256'hcc00b200a20099009c00aa00c300e200000111010f01f300bd007c003d001000;
    inBuf[8819] = 256'h01000d0026003e004c004c0045003c003b004200450038001800deff96ff58ff;
    inBuf[8820] = 256'h32ff2eff4fff82ffafffcbffccffaeff7bff42ff11fff5feebfeebfeeffeebfe;
    inBuf[8821] = 256'hd8fec0feaafea3feb0fec2fecdfecffec3feadfe98fe81fe62fe3bfe0bfedffd;
    inBuf[8822] = 256'hcafdd3fdf8fd2bfe57fe6efe6cfe4dfe25fe02fee2fdc9fdb8fda7fd94fd87fd;
    inBuf[8823] = 256'h7dfd7cfd8bfda2fdbdfdd6fddcfdcbfda8fd75fd3ffd14fdf3fcddfcd3fccffc;
    inBuf[8824] = 256'hd3fcdbfce0fce6fceefceefcf0fcf6fcebfccefca6fc71fc3dfc1cfc0afc0efc;
    inBuf[8825] = 256'h27fc44fc64fc8dfcacfcbcfcbcfc9efc6cfc3afc0efcf3fbeefbf1fbf3fbf4fb;
    inBuf[8826] = 256'hf1fbfbfb18fc39fc5dfc7afc78fc5bfc2dfce8fb9ffb65fb3ffb3ffb67fb96fb;
    inBuf[8827] = 256'hbffbd3fbc2fba6fb94fb85fb84fb90fb8cfb7bfb69fb4dfb34fb27fb17fb0afb;
    inBuf[8828] = 256'h08fb08fb19fb40fb66fb89fba0fb95fb7bfb5ffb39fb1afb0dfb00fbf7faf8fa;
    inBuf[8829] = 256'hf6fafafa07fb0ffb20fb41fb5cfb70fb77fb5bfb2afbf2fab8fa98fa98faa1fa;
    inBuf[8830] = 256'hb7fad5fae5faf2fa06fb16fb31fb4ffb58fb4efb2ffbeefaa8fa77fa5cfa6efa;
    inBuf[8831] = 256'ha7fae9fa29fb57fb5ffb55fb48fb34fb25fb17fbf9fad7fab1fa83fa66fa66fa;
    inBuf[8832] = 256'h71fa93facbfafffa2efb51fb5afb57fb4bfb26fbfbfacffa9ffa84fa89fa9ffa;
    inBuf[8833] = 256'hcdfa08fb33fb56fb74fb80fb88fb8dfb81fb6ffb58fb34fb12fbfdfaf2fafffa;
    inBuf[8834] = 256'h26fb52fb7cfb98fb96fb83fb6dfb5afb57fb5bfb55fb4efb3cfb14fbf3fae5fa;
    inBuf[8835] = 256'he5fa06fb43fb80fbb6fbdbfbd7fbb7fb90fb67fb50fb4efb51fb5efb71fb82fb;
    inBuf[8836] = 256'ha4fbd8fb08fc35fc5cfc6bfc6dfc67fc50fc2dfcfffbc6fb9cfb90fb9bfbc7fb;
    inBuf[8837] = 256'h09fc42fc71fc98fca5fc9efc84fc55fc22fcfbfbdffbd4fbd4fbcdfbcffbe0fb;
    inBuf[8838] = 256'hfefb36fc7ffcbbfce4fcf3fce3fcc5fca8fc8bfc79fc71fc6bfc72fc8afca7fc;
    inBuf[8839] = 256'hcefc01fd33fd67fd92fda4fd9cfd75fd32fdf2fcc4fca5fca4fcbbfcd8fcfffc;
    inBuf[8840] = 256'h30fd5efd8bfdb0fdbcfdb3fd97fd67fd37fd14fd02fd0bfd27fd41fd5afd6dfd;
    inBuf[8841] = 256'h7afd96fdc5fdfefd3cfe6cfe78fe67fe3ffe02fec7fda2fd95fda5fdccfdfbfd;
    inBuf[8842] = 256'h2afe4cfe63fe7dfe9bfeb6fec9fec6fea6fe73fe36fefefde0fddafde8fd0afe;
    inBuf[8843] = 256'h35fe62fe96fec7feedfe0eff24ff26ff1cff02ffd7feacfe8cfe85fea1fed8fe;
    inBuf[8844] = 256'h19ff5bff92ffbaffd4ffe1ffe0ffd2ffb2ff85ff55ff28ff09ff02ff0fff2eff;
    inBuf[8845] = 256'h5aff8affb5ffd9fff2ff01000800ffffe3ffb6ff7aff42ff22ff24ff4aff8eff;
    inBuf[8846] = 256'hdfff2f007200a300c000c400ae0087005900340029003700520073008f00a200;
    inBuf[8847] = 256'hb700d500f900210142015401550144011f01ed00b600830063005e007500a600;
    inBuf[8848] = 256'hde000c012b01390135012a0121011a0114010b01fd00ee00e600f00018015c01;
    inBuf[8849] = 256'haf01ff01340241022c020102d401bb01b701c301d901ed01f601fd0105021502;
    inBuf[8850] = 256'h3a026a029602af02a40271022802dc01a2018c019501b101de010e023b026802;
    inBuf[8851] = 256'h8d02a302ad02a80295028202700257024202350233024a027a02b802fa023503;
    inBuf[8852] = 256'h5c037003720368035a0341031b03f302cc02ac02a202af02d00200032d034e03;
    inBuf[8853] = 256'h6a0375036a035d034a0329030603e402c502b602c002e002160351038503ad03;
    inBuf[8854] = 256'hbf03c103c703c603bb03b0039c037b0361035203500363038303af03ea031c04;
    inBuf[8855] = 256'h3a044b04440425040304dd03b0038803620344033e034b0361038303a303bd03;
    inBuf[8856] = 256'he103060421042f042004f003b90388036803640373038a03b303e9032a047204;
    inBuf[8857] = 256'ha504b0049b046a0436041b040d040404fe03ee03dd03e50302042c045c047604;
    inBuf[8858] = 256'h72045d0434040004d703b4039903920392039803a903b803c703e40307042a04;
    inBuf[8859] = 256'h4b04550445042704f603c003a3039a03a203c103eb0318044b0478049904b104;
    inBuf[8860] = 256'hb2049d047b0449041004dc03ac038d038c039803af03d303f503120431044604;
    inBuf[8861] = 256'h4e0447042404ec03ad036a03320317031303250352038d03cd03100443045f04;
    inBuf[8862] = 256'h6c04630443041104cc037d0338030d030e033e037f03be03f1030b0418042c04;
    inBuf[8863] = 256'h390432040b04b8034903e602a3028d02a602d102010337036d03a103d703f803;
    inBuf[8864] = 256'hf203cc038a033803ee02b302880276028102b00202036103b303ea03f603de03;
    inBuf[8865] = 256'hb9038d035d032603df0290024d0221021d0246028702cf0212033a0342033003;
    inBuf[8866] = 256'h0403cc0296025e022d020d02f601e901ed01fd011f0259029902d30200030803;
    inBuf[8867] = 256'hed02c3029502700258023f021e02f801d401cd01f0012d026f02a002a8028f02;
    inBuf[8868] = 256'h6c0246022002fa01c60185014a0123011c01340158017e019b01a901b201b701;
    inBuf[8869] = 256'hb1019f0185015f0138011301f200e000e700fd00230155018301ab01cb01da01;
    inBuf[8870] = 256'hd301af016f012701ec00c900c100c700c700c100be00cb00f0001a012b011801;
    inBuf[8871] = 256'hde008b0043001700fefff7fff9fffaff070024004500620075007b0079007200;
    inBuf[8872] = 256'h610042001600e9ffd2ffdcff030031004a004500320025002b00450055004200;
    inBuf[8873] = 256'h0900baff74ff4cff41ff45ff49ff42ff3bff46ff5dff78ff90ff96ff85ff67ff;
    inBuf[8874] = 256'h3dff0affd6fea5fe84fe80fe9afecdfe10ff51ff86ffa9ffb5ffadff93ff6fff;
    inBuf[8875] = 256'h49ff24fffcfed1fea3fe74fe57fe60fe89fec5fefbfe10ff03ffe5fec3fea7fe;
    inBuf[8876] = 256'h8bfe59fe0ffebcfd75fd59fd6efda0fddafd0bfe2cfe48fe60fe6afe61fe48fe;
    inBuf[8877] = 256'h25fe08fef9fdeafddafdc9fdc3fddefd22fe6dfe9ffeaafe8efe69fe58fe5afe;
    inBuf[8878] = 256'h5cfe3ffef1fd8dfd41fd29fd46fd78fd91fd86fd66fd4afd4ffd6ffd84fd73fd;
    inBuf[8879] = 256'h3efdf9fcc5fcb8fcc6fcdafce3fce0fce5fc04fd39fd76fda4fdb4fdaefda2fd;
    inBuf[8880] = 256'h96fd8ffd8ffd8bfd7bfd60fd41fd2bfd26fd39fd67fd97fda5fd89fd4dfd07fd;
    inBuf[8881] = 256'he3fcecfc03fd0afde9fc9dfc4cfc21fc24fc4bfc78fc86fc7dfc76fc7afc8efc;
    inBuf[8882] = 256'haafcb4fcacfca3fca3fcb9fcd9fce8fce5fce3fcebfc0afd33fd45fd38fd15fd;
    inBuf[8883] = 256'hf0fcecfc09fd21fd1dfdfefccffcb3fcb7fcc3fcbffc9cfc5bfc28fc1dfc2cfc;
    inBuf[8884] = 256'h40fc3bfc0efcdbfbc6fbd8fb0ffc4dfc6dfc6efc68fc6afc87fcb0fcc8fcc4fc;
    inBuf[8885] = 256'ha6fc79fc61fc76fcaefcf7fc30fd43fd3bfd28fd18fd23fd3efd47fd2dfde9fc;
    inBuf[8886] = 256'h84fc2efc05fc07fc27fc44fc3bfc19fc00fc04fc2efc62fc72fc51fc0dfcc9fb;
    inBuf[8887] = 256'haffbc1fbdffbf4fbf0fbe1fbfafb4cfcb6fc16fd4dfd4dfd35fd29fd33fd47fd;
    inBuf[8888] = 256'h41fd0ffdccfc9cfc94fcbcfcf8fc20fd2cfd24fd18fd1cfd26fd18fde9fc97fc;
    inBuf[8889] = 256'h36fcecfbbffba1fb96fb97fba1fbc8fb0efc59fc98fcbcfcbafca8fc99fc8efc;
    inBuf[8890] = 256'h8bfc85fc71fc5bfc52fc5efc8dfce0fc44fda5fdeefd0afefefddefdbefdaefd;
    inBuf[8891] = 256'ha3fd80fd3cfde3fc93fc78fc9ffce6fc1efd21fdeefcb0fc97fcaefcddfcecfc;
    inBuf[8892] = 256'hb4fc4dfceefbc8fbf4fb52fca1fcc1fcbbfcb5fcdbfc37fd9dfdd9fdcefd8dfd;
    inBuf[8893] = 256'h53fd4cfd79fdbbfde4fddafdb8fda7fdc3fd0afe4ffe5ffe33fee0fd8afd5efd;
    inBuf[8894] = 256'h5cfd64fd62fd4afd1bfdf4fceafcf6fc0efd22fd25fd25fd27fd26fd27fd2afd;
    inBuf[8895] = 256'h27fd29fd39fd54fd7afda5fdcafdedfd15fe40fe70fe9dfeb5feb9feadfe95fe;
    inBuf[8896] = 256'h82fe7dfe81fe8dfe9afe9cfe91fe7efe67fe56fe4dfe44fe32fe10fee0fdb4fd;
    inBuf[8897] = 256'h98fd8efd94fd9cfd99fd98fda9fdd8fd1efe5efe77fe64fe39fe1afe2afe64fe;
    inBuf[8898] = 256'ha0febefeb2fe97fea3fef4fe75fff1ff2c001300cbff92ff8fffb8ffd4ffb2ff;
    inBuf[8899] = 256'h4effd7fe8efe9afee5fe31ff47ff1dffe1fed0fefbfe40ff65ff3affc4fe47fe;
    inBuf[8900] = 256'h07fe1efe71fec4fee7fedbfec7fedcfe31ffacff1c0058005a003b0024002d00;
    inBuf[8901] = 256'h4d00680064003e001000fdff18005900a000c800c10098006e005f006a007600;
    inBuf[8902] = 256'h5f001700b3ff62ff4eff7fffccff0000faffc8ff99ff9bffdbff36006c005a00;
    inBuf[8903] = 256'h1900e7fff5ff4600ac00e800e100bc00b300ed005a01b901ce0194013c010e01;
    inBuf[8904] = 256'h2f017c01ac0193013701d600bf0003016e01b2019b013201bf008c00ad00f800;
    inBuf[8905] = 256'h25010801b5006600560099000301540169014d0127012a016301b501f201fc01;
    inBuf[8906] = 256'hd601a901a201d20126026e027d0250020b02e801070253029702a0025f02f701;
    inBuf[8907] = 256'hb201ba0103024d0258021502b30173018101d0011c022102db01800158018a01;
    inBuf[8908] = 256'hf4014c025f022b02ed01ee013f02b4020603ff02b2026e026f02bc0224035a03;
    inBuf[8909] = 256'h3b03ee02b302bc020803580367032c03ca0286029502df021e031f03d3026a02;
    inBuf[8910] = 256'h36025402a502ed02eb029a023d0218024402ae0207030f03d3028a027c02d002;
    inBuf[8911] = 256'h5a03c203cf037e031203e50218038403dd03de038703270308034703c4032204;
    inBuf[8912] = 256'h1b04c3035c032d035503a303c60395031d03a8028a02cf023f038e0381032803;
    inBuf[8913] = 256'hd602cc0218039203e103d1037a031b03f90232039503de03ea03bb0384037f03;
    inBuf[8914] = 256'hb103fa0330042704ea03ae039603ab03d903ef03d503a20373036a039303c603;
    inBuf[8915] = 256'hd503b70376033e033c0364039303a8038b03550340036103a803f2030a04e303;
    inBuf[8916] = 256'ha7037d038103ba03f7030904ee03b8038c039703cb0300041a040604d503b703;
    inBuf[8917] = 256'hb703cb03df03d1039a035c033503340359037d03830371035503450356037903;
    inBuf[8918] = 256'h94039a03800351033303330350038403b103c103ba03a6039b03ac03ce03ee03;
    inBuf[8919] = 256'hfa03dd03a1036703430340035d03780379035f03380324033f03710397039403;
    inBuf[8920] = 256'h5603f402a8028b02a102ce02dd02bd028d0270028702dd023f037d0383035603;
    inBuf[8921] = 256'h1c0304030f0324032c030d03d402ac02a802ce020d033a033f032c0311030603;
    inBuf[8922] = 256'h14031a03fb02b9025e020f02f30107022f024a023602fc01cf01d2010a025e02;
    inBuf[8923] = 256'h930282023a02e601ba01d50118024f0258022e02f601e701090243026b026502;
    inBuf[8924] = 256'h40022802340257026e024f02fe01b0019701c30109021c02d2014601c500a300;
    inBuf[8925] = 256'hf3006e01af017d01f20070005300a7002b017a015301d60067005900bb004801;
    inBuf[8926] = 256'h960176011001bb00ca003d01bf01f001ab011901a4009900f100590173011701;
    inBuf[8927] = 256'h820021003800b70040015c01e40017006cff45ffa1ff19003800d3ff22ffa0fe;
    inBuf[8928] = 256'hb3fe53ff170082005500c6ff51ff54ffcbff5a008d0038009fff34ff48ffccff;
    inBuf[8929] = 256'h5f0099005f00f0ffb5ffe8ff6300bf00a7001b0070ff0cff1aff68ff92ff57ff;
    inBuf[8930] = 256'hcdfe50fe35fe83fef2fe20ffe2fe60fefefd08fe72fee8fe09ffb3fe25fec5fd;
    inBuf[8931] = 256'hd6fd4dfed9fe1cfffcfea8fe71fe90fefbfe69ff93ff65ff0affccfedafe1eff;
    inBuf[8932] = 256'h58ff51fff8fe81fe35fe3afe7cfeb3fe99fe27fe99fd40fd4ffdaefd0afe0ffe;
    inBuf[8933] = 256'hadfd1cfdbefcd5fc4cfdcdfdfcfdb8fd38fde2fcfbfc7bfd13fe64fe4bfef5fd;
    inBuf[8934] = 256'hb5fdcafd2bfe8ffeaefe74fe0dfec3fdc0fdf6fd32fe42fe1dfee6fdc2fdbbfd;
    inBuf[8935] = 256'hc0fdb2fd83fd45fd0efdedfcdffcd0fcadfc80fc5bfc4dfc5bfc7cfca1fccafc;
    inBuf[8936] = 256'hf0fc09fd14fd0dfdfbfcf4fc09fd32fd61fd7bfd6efd51fd42fd57fd99fde7fd;
    inBuf[8937] = 256'h12fe0bfee4fdb6fda2fda6fda3fd88fd4efd00fdbdfc93fc75fc5afc42fc32fc;
    inBuf[8938] = 256'h3efc62fc85fc92fc81fc5cfc45fc4bfc5ffc6cfc62fc42fc2cfc36fc60fc9bfc;
    inBuf[8939] = 256'hcffceffc07fd26fd50fd85fdb5fdd2fddcfdd4fdbefda0fd7afd51fd2ffd17fd;
    inBuf[8940] = 256'hfffce3fcc1fca2fc99fca8fcbefcc7fcaefc76fc45fc3bfc5afc81fc7efc38fc;
    inBuf[8941] = 256'hd1fb85fb87fbe0fb58fca3fcabfc8efc8dfcdbfc60fdcdfde1fd94fd27fdfdfc;
    inBuf[8942] = 256'h38fda5fdf0fdd2fd5cfdeefce3fc50fdf6fd5efe37fe9dfdf4fca1fccafc2dfd;
    inBuf[8943] = 256'h59fd0ffd61fcaefb6cfbbdfb60fcebfc07fdb1fc49fc34fc91fc29fd8cfd6bfd;
    inBuf[8944] = 256'he2fc5ffc54fce4fcbafd49fe3afeaefd28fd31fde3fdd1fe59ff14ff2dfe4dfd;
    inBuf[8945] = 256'h0dfd89fd4dfeabfe41fe55fd92fc8afc45fd32fe8ffe0dfe04fd2efc21fccdfc;
    inBuf[8946] = 256'h98fdd6fd51fd76fc05fc69fc6cfd5ffea0fe14fe48fdf1fc67fd62fe2eff3dff;
    inBuf[8947] = 256'h97feccfd87fd0ffe0dffd0ffd7ff28ff51fef5fd4efe07ff81ff42ff5efe69fd;
    inBuf[8948] = 256'hfcfc56fd27fec7febffe24fe79fd50fdd4fd9dfe03ffa7feb9fdddfcb5fc5bfd;
    inBuf[8949] = 256'h55fef4fed6fe37fec4fd0dfe0dff3200c1006c008bffd8fed9fe7bff20002900;
    inBuf[8950] = 256'h7cff99fe37feb0feb2ff7e008000c1ffddfe85fee9fe94ffd5ff4dff46fe76fd;
    inBuf[8951] = 256'h6bfd1cfef6fe53ff00ff63fe20fe8efe76ff36004c00b9ff01ffbffe2dfff6ff;
    inBuf[8952] = 256'h84007800f0ff71ff7aff1e00f5006d013c019600fcffd8ff3400ae00cf006d00;
    inBuf[8953] = 256'hc5ff48ff4bffbdff35004c00e3ff3effd0fee4fe5fffe0ff0100aaff22ffd7fe;
    inBuf[8954] = 256'h0cffa6ff40007c004c00f9ffedff570006018b018f011c0199007700de008701;
    inBuf[8955] = 256'hf301cc012d0187005000ab00440192014a019600efffc9ff3700d2000f01af00;
    inBuf[8956] = 256'heaff48ff3effcbff8100d7008e00e7ff73ffa1ff64003e019a01410189001000;
    inBuf[8957] = 256'h4d0035013602a60243025f01b200ce00a5019f0208038c028401b100a5005701;
    inBuf[8958] = 256'h2e026b02c901af00d7ffd1ff8c006201a00112011f0081ffb3ff870052017901;
    inBuf[8959] = 256'he2001200c0ff3f00420117022e029001d800b4005c0166021c030a0353029501;
    inBuf[8960] = 256'h6601e1019b02f902af02f70165016001d8015c027202f9014401cf00d8003401;
    inBuf[8961] = 256'h73013e01aa001c00f9ff5700ee0047012801c0007900a9004601f10143021a02;
    inBuf[8962] = 256'hae016901940117029c02cd02950239021c026102e4024b034503d4024502ef01;
    inBuf[8963] = 256'hfa01410267023202b1012801ea000e015b01850162010101ae00ac00f3004a01;
    inBuf[8964] = 256'h67012901c0008400a60019019d01e501d801af01bc012702c80246035a030a03;
    inBuf[8965] = 256'ha0027502a8020a03410314039a0229020f025102a602b7026102d10166016001;
    inBuf[8966] = 256'ha401d601a00100014d00fdff4100e20060015901df006a007d0039013102c602;
    inBuf[8967] = 256'h9502ca0110010e01dd01f7029b035e038302cc01dc01c002d9035504d803bd02;
    inBuf[8968] = 256'hd601ca018702530364037a021401230042003901370260027e01350077ffcbff;
    inBuf[8969] = 256'hee00f90113022d01feff7aff1f008d01c702ff022b020e01a3005b01c002de03;
    inBuf[8970] = 256'hf7031003ed017d01180246031c04f303e502be014f01d201c5024703d2029e01;
    inBuf[8971] = 256'h76001600a600910100028901730086ff71ff39003901a6012b012b0078ffacff;
    inBuf[8972] = 256'hb800ef017f0220024701bb000801150230039f0329033c029e01d201b1028f03;
    inBuf[8973] = 256'hbb030803ed0124012a01dd0192029d02d301a300caffc4ff6b0022014901b400;
    inBuf[8974] = 256'hc7ff2fff5aff260000014c01df00130083ffa3ff6a005901e401d1015701f400;
    inBuf[8975] = 256'h1301bc018802fd02da024202a9017c01d2015f02b5028602e0012501c100de00;
    inBuf[8976] = 256'h5101ab019101f80029008fff6dffaeff01000e00b6ff30ffdefe00ff91ff4300;
    inBuf[8977] = 256'hb200b3006c0028002c008900090163016a013101f800fa004101ae0108022402;
    inBuf[8978] = 256'h0402d101b701c201d601c2016e01e90060000100dcffe5ffefffd7ffa0ff68ff;
    inBuf[8979] = 256'h4eff60ff87ff9fff90ff5bff1afff7fe07ff38ff6eff93ffa7ffc1fffcff5a00;
    inBuf[8980] = 256'hc6001f0150015b0158015f01740188017e014801f400a5007d008700b000cc00;
    inBuf[8981] = 256'hb80071001800d6ffc1ffc7ffbaff73fff9fe81fe46fe5ffeaefee9fed9fe8cfe;
    inBuf[8982] = 256'h46fe54fed5fe91ff1f003600deff73ff63ffd0ff7a00f400ea00760010002700;
    inBuf[8983] = 256'hce00a0010302a901d0000c00ddff4d00de00ee003e0025ff50fe39fec7fe65ff;
    inBuf[8984] = 256'h73ffcffeeefd74fdbefd91fe40ff3aff88febffd88fd1efe1cffceffc8ff3aff;
    inBuf[8985] = 256'hcafe02ffe4ffde003f01cf00faff7bffc5ffa5006a017501bc00d1ff6cffd1ff;
    inBuf[8986] = 256'h9b00090199007aff68fe15fe9cfe66ffa1ffe9fea5fdb1fcbbfcb6fddbfe4aff;
    inBuf[8987] = 256'hb1fe95fdeefc58fd94fec4ff0b003cff13fe9ffd63fe01006e01b601cc0088ff;
    inBuf[8988] = 256'hfdfeb1ff250136020502a40002ff43fed6fe21000201ab0042ffc5fd3cfdf1fd;
    inBuf[8989] = 256'h3bff0500a4ff57fe07fd92fc23fd22feaffe60fe85fddffc06fdf1fd0bffaaff;
    inBuf[8990] = 256'h90ff0dffb8feeefe94ff3d00880068001d00010030007d00a80093005a003100;
    inBuf[8991] = 256'h310044003b00f3ff7dff0affc2fea1fe87fe51fe00febefdacfdcafdf3fdf7fd;
    inBuf[8992] = 256'hc4fd77fd50fd7ffdf6fd74febbfeb5fe89fe84fed2fe66ff05005d004a00faff;
    inBuf[8993] = 256'hb8ffbfff1d009d00ef00e90094002800e8fff1ff27004e002d00bdff2fffbcfe;
    inBuf[8994] = 256'h88fe90fe9ffe80fe2afec1fd7dfd84fdcbfd1afe3bfe1efee2fdbefdd8fd2bfe;
    inBuf[8995] = 256'h8afec5fed5fee0fe18ff8eff22008f00a4006f0034003d00a3002a0169012501;
    inBuf[8996] = 256'h7e00d4ff8effcdff3c006100fbff36ff91fe7afeedfe73ff78ffc1fea7fddcfc;
    inBuf[8997] = 256'he4fcacfd8cfecbfe39fe57fdf4fc8efde1fe110053008eff84fe35fe12ff9c00;
    inBuf[8998] = 256'hc301b10180002cffd2fed5ff8801a7025c02e6005effecfed6ff4301ed012201;
    inBuf[8999] = 256'h48ff9afd33fd32feacff5d00aeff1efed9fcc2fcd3fd21ffa2ff00ffcefd0efd;
    inBuf[9000] = 256'h64fd96fec2ff1f0093ffc2fe82fe31ff70007601aa0112014a00040074003b01;
    inBuf[9001] = 256'hbf019d01ed003300e8ff22009a00df00ae00220084ff13ffe3fedbfed3feb8fe;
    inBuf[9002] = 256'h8cfe59fe2bfe04fef3fd0dfe54feb0fef8fe08ffe9fed4fe02ff7bff0e006400;
    inBuf[9003] = 256'h4b00e4ff97ffc2ff6e004101c201a9011d0199008500e20055016801ee002f00;
    inBuf[9004] = 256'ha8ffa6ff0600570032008dffc3fe54fe77fef0fe4aff2fffa2fe04fec3fdfcfd;
    inBuf[9005] = 256'h7dfeebfe07ffe3fec8fef4fe6dff0000690086006d00560064009300ce00f900;
    inBuf[9006] = 256'h0d0112011901240126011401f300d100b200900062001a00c1ff6cff29ff00ff;
    inBuf[9007] = 256'heefee4fed8fec9feb5fea3fe9efea7fec6fef7fe23ff33ff1affe4febffedbfe;
    inBuf[9008] = 256'h45ffe0ff6b00ae009f006f006300aa002901900198013d01be0076009500fc00;
    inBuf[9009] = 256'h51013b01af00fcff8dff99fff8ff470028008effc7fe3ffe37fe93fef3fefefe;
    inBuf[9010] = 256'ha9fe3dfe19fe6efe15ffaaffd6ff8fff21fff3fe3dffe4ff9000ed00e300a100;
    inBuf[9011] = 256'h7a00a00006016f019d0179011f01c8009c009d00ac00a10068001200baff79ff;
    inBuf[9012] = 256'h5fff69ff85ffa1ffa2ff71ff12ffa5fe59fe59fea5fe0aff43ff23ffc3fe7dfe;
    inBuf[9013] = 256'ha0fe3aff05008d008a001900a8ffacff48002101a7018101d3002a001000a300;
    inBuf[9014] = 256'h7f01ff01bd01e6001500d7ff4200e1000d0176005dff69fe25fe9dfe59ffb7ff;
    inBuf[9015] = 256'h69ffb0fe1bfe1dfebafe7cffdaffa2ff11ffa0febcfe65ff3000a60095002900;
    inBuf[9016] = 256'hceffdcff5f0015019c01b6016c01fc00a9009700b600da00dc00a7004e00fdff;
    inBuf[9017] = 256'hd8ffebff1d003b001c00bdff47fffbfe01ff47ff8dff8dff31ffaffe5cfe73fe;
    inBuf[9018] = 256'hebfe73ffb2ff8fff41ff25ff7aff2500c100f000a0002800fdff5d002101d101;
    inBuf[9019] = 256'hf5018001d200670085000201630143019e00ceff52ff70fff2ff61005d00d8ff;
    inBuf[9020] = 256'h22ffaffebdfe2effa0ffb7ff5cffd3fe81fea1fe20ffacfff2ffd6ff8eff75ff;
    inBuf[9021] = 256'hc0ff5b00f0002901ec0071001c002f00a30025015c012a01c10076008600e400;
    inBuf[9022] = 256'h3f014401da003c00c5ffb1fff5ff4a005d000d0084ff0effe6fe14ff61ff8aff;
    inBuf[9023] = 256'h6eff20ffd9fed0fe12ff7dffd2ffe3ffbdff97ffaaff1400b300350159011501;
    inBuf[9024] = 256'h9e004f006200c5002a014401fa008b0056008d000501570126017600acff4eff;
    inBuf[9025] = 256'h91ff2a008900470074ff9cfe5afedbfec0ff62005100aafffcfed4fe53ff1000;
    inBuf[9026] = 256'h7000280073ffe7fe01ffc5ffb70047013501ba005d007800f70074017f010601;
    inBuf[9027] = 256'h620001001b008c00f000fa00ae0051002e005a009800a1005400cbff48ff01ff;
    inBuf[9028] = 256'hf8fe0aff0ffffdfeedfe02ff44ffa1fff7ff2b00460059006b0072005e002a00;
    inBuf[9029] = 256'hedffcdfff0ff5400c80011011201da00a700a900e600330150010d017f00f0ff;
    inBuf[9030] = 256'ha6ffbeff100048002e00caff61ff47ffa0ff3800a6009100f1ff1dff95fea1fe;
    inBuf[9031] = 256'h2bffc8ff0d00d6ff64ff26ff6bff1d00d0001401c3002200b0ffc3ff52000001;
    inBuf[9032] = 256'h540119018b0022003d00db009601eb019301ba00dbff73ff9fff0d003f00e9ff;
    inBuf[9033] = 256'h2aff7cfe5dfef3fee5ff9900a3000d004affe3fe1affbbff49005600dcff46ff;
    inBuf[9034] = 256'h0dff6aff3300f500420106018400220024007900cd00dc0098002e00ebffffff;
    inBuf[9035] = 256'h5700b400e600df00b80097008d0083005300f2ff7dff1dfff6fe08ff30ff4eff;
    inBuf[9036] = 256'h5fff70ff9bffe1ff210033000d00c0ff78ff5cff72ff9cffbcffcbffdfff1500;
    inBuf[9037] = 256'h7200de0030015201500148014d0153012c01bc00160079ff2fff55ffc1ff2700;
    inBuf[9038] = 256'h4b002600ebffd8fffaff2d003700efff6affeefebcfee4fe43ff99ffbcffb0ff;
    inBuf[9039] = 256'h9effb1fff7ff530092008e005000ffffc7ffbfffdfff0800270043006900af00;
    inBuf[9040] = 256'h1401710196016b01fe007e002100fdfffdfff3ffbdff5eff09ff02ff5efff0ff;
    inBuf[9041] = 256'h67007d001f0089ff1aff08ff46ff91ff9aff46ffd2fe98fed6fe85ff5500e600;
    inBuf[9042] = 256'h0a01dc00a0009500c60002010a01c5005000e8ffc2ffeaff43009a00cf00d700;
    inBuf[9043] = 256'hbd008e0053001200d6ffabff96ff8fff80ff5aff2dff18ff32ff7affccfff8ff;
    inBuf[9044] = 256'he6ffb0ff88ff92ffc0ffdbffb3ff4effebfee2fe61ff3b00fb0041010901a500;
    inBuf[9045] = 256'h8500e0007b01d401810192008dff19ff77ff5200fa00e3000d0017ffc3fe5fff;
    inBuf[9046] = 256'h83005d013e012400c3fefffd43fe38ff080004002cff34feeafda5feffff1701;
    inBuf[9047] = 256'h45019600b8ff6fff01000001a2016a01820096ff51ffdbffba003a01fc003e00;
    inBuf[9048] = 256'ha1ffacff600033017e010301100048ff27ffa7ff49007700f6ff0fff5dfe5afe;
    inBuf[9049] = 256'hfffed8ff520020006dffbefe92fe0dffddff7a00880015008aff5fffc5ff8600;
    inBuf[9050] = 256'h26014501e00056001c006900070178015801aa00d9ff6effa8ff4d00d900dc00;
    inBuf[9051] = 256'h480089ff29ff64fff9ff5f002f0074ffa2fe44fe97fe5bfffeff0a0087ffecfe;
    inBuf[9052] = 256'hc5fe4cff420016014801c700faff6eff7aff0700a300e0009f001e00d0ff0000;
    inBuf[9053] = 256'h97003601790136019d000f00dcff090054006f003a00d0ff76ff66ffa0fff0ff;
    inBuf[9054] = 256'h1400ecff8eff35ff0bff17ff3dff4cff32ff09ff01ff3bffb0ff3900a200ca00;
    inBuf[9055] = 256'hb6008f0082009800bf00d100ac005200efffbbffddff4b00ca0019011701d200;
    inBuf[9056] = 256'h86006a007e0092006a00edff46ffc4fea6feeefe58ff92ff84ff53ff48ff93ff;
    inBuf[9057] = 256'h16007c007e0018008eff40ff58ffb3ff08001800eeffd1ff0300850013015801;
    inBuf[9058] = 256'h2c01b2003d00170045008a00a700860044001c002f006f00ac00b80087003800;
    inBuf[9059] = 256'hebffabff75ff40ff07ffd5febafec3fef1fe3cff9cff0d007600b600b9007e00;
    inBuf[9060] = 256'h2800e7ffd2ffe2fff5ffecffc8ffb2ffd5ff4000cf0041016b014e011401ed00;
    inBuf[9061] = 256'he400d6009c00270095ff26ff10ff4effb6ff090020000400ddffceffdffffcff;
    inBuf[9062] = 256'h0000d9ff8cff3bff0aff0eff48ffa2fff8ff350054005e006a008900ab00b500;
    inBuf[9063] = 256'h90003b00dfffb9ffe3ff4b00ba00ed00d0008f006e009900fa0040011f018300;
    inBuf[9064] = 256'ha9fffffed0fe15ff83ffb9ff93ff3fff16ff5bff0400b000f500a900fbff53ff;
    inBuf[9065] = 256'h19ff5cffd5ff23000a00a6ff54ff6afffbffc700620180012f01ba007b009200;
    inBuf[9066] = 256'hd400f000ad001e0099ff6effb2ff2f0089007d001a00a6ff73ffa0fffaff2f00;
    inBuf[9067] = 256'h1100aeff47ff29ff67ffd1ff25002e00f1ffadff9dffd2ff2800660063002400;
    inBuf[9068] = 256'hd5ffb1ffd9ff38009e00da00da00b70096009200b000d400cc008d002e00d1ff;
    inBuf[9069] = 256'h9effa5ffc7ffdfffd8ffb8ffa3ffb5ffe6ff19002b000c00d1ffa1ff9bffb5ff;
    inBuf[9070] = 256'hcdffc9ffacff8dff90ffc9ff1d005f0074006000420041006600a300d300d400;
    inBuf[9071] = 256'ha7006a00370024003600570069005e002c00e5ffa6ff8aff9bffd0ff09001f00;
    inBuf[9072] = 256'h0500d0ffa9ffaeffe2ff210034000300a7ff5dff59ffa2ff0a004b004000fbff;
    inBuf[9073] = 256'hb9ffbcff12008c00e600ed00a6004a001700290069009e009c0061001400e8ff;
    inBuf[9074] = 256'hf3ff210048003a00eeff90ff5cff6dffbaff10002e000000a9ff5fff61ffbbff;
    inBuf[9075] = 256'h33007e006a00feff7fff44ff78fffcff770099005700efffc2ff05009e003601;
    inBuf[9076] = 256'h6c0113016800daffb5fffeff68008b003d00a6ff24ff11ff79ff11007b007c00;
    inBuf[9077] = 256'h1f00b2ff7fffa0fff0ff2a001b00cbff72ff4bff6effbdff01001300f8ffd7ff;
    inBuf[9078] = 256'hddff0e0054008f009e0085006600590067008100910090007f00620041002100;
    inBuf[9079] = 256'h0200e4ffcfffc4ffbeffb6ffabffa3ffb0ffd7ff06001400efffabff6eff5fff;
    inBuf[9080] = 256'h89ffc7ffe3ffc1ff74ff3bff5affd7ff6f00d300d7008d0043003f008400da00;
    inBuf[9081] = 256'hf600ad002600bbffb2ff05007200a20074000f00c3ffc4ff02003c003200d7ff;
    inBuf[9082] = 256'h62ff22ff3aff8effdaffe2ffa7ff67ff62ffa8ff0a003f001c00b7ff56ff40ff;
    inBuf[9083] = 256'h81ffeaff390049002d001e0045009f00ff002f011701d00082004f0039002a00;
    inBuf[9084] = 256'h1100e8ffbaffa2ffabffc8ffecff07000c00ffffe7ffc6ff9fff78ff56ff38ff;
    inBuf[9085] = 256'h28ff2bff40ff5eff80ff9fffb9ffdbff0d004a008500a1008d00580022001100;
    inBuf[9086] = 256'h38007b00ac00ae0080004500300053009000b2008a001d00a7ff6bff85ffd4ff;
    inBuf[9087] = 256'h11000600b5ff53ff2dff63ffcaff16001000b3ff38ffe9feedfe36ff87ffaaff;
    inBuf[9088] = 256'h96ff72ff78ffc6ff4600c30009010101c300820069008500af00b4007f002200;
    inBuf[9089] = 256'hd4ffc9ffffff510088007d003c00f3ffd2ffeaff14001200d0ff65ff02ffdbfe;
    inBuf[9090] = 256'hfbfe3aff67ff67ff49ff3aff55ff97ffe2ff100015000a0009001c0039004500;
    inBuf[9091] = 256'h38002a00340060009c00c000ac006c00390041008000c500d3008900050099ff;
    inBuf[9092] = 256'h81ffbcff11003100f8ff87ff2dff26ff6fffcbfff0ffb9ff45ffdefec2fef8fe;
    inBuf[9093] = 256'h58ffa9ffcaffc4ffb6ffc1fff4ff43009500d000e400ca00860037000e001e00;
    inBuf[9094] = 256'h57008e008d004800f2ffd9ff2200a8000701f2006300aaff3eff5affc9ff1600;
    inBuf[9095] = 256'he2ff35ff86fe57fecdfe9cff34003000abff1eff03ff80ff3c00ab007b00d4ff;
    inBuf[9096] = 256'h38ff23ffafff82001301120199001200ebff4100cf00270107017e00e6ff9dff;
    inBuf[9097] = 256'hbeff2000750080004100e9ffadffa9ffc9ffe1ffcbff86ff2ffff3fef0fe21ff;
    inBuf[9098] = 256'h5dff7fff88ff8effa6ffdeff260059005a002f00fffff2ff09002f0046003800;
    inBuf[9099] = 256'h120005002d008100db000601e60094004100190024003a003100ffffb7ff7eff;
    inBuf[9100] = 256'h72ff8fffbaffd4ffcfffb3ff98ff8cff8eff8dff80ff6fff6aff7bff9affbdff;
    inBuf[9101] = 256'hdefffaff17003f0067007c007a0067004c003a002e0022002200300045006200;
    inBuf[9102] = 256'h7e0086007d006a005900540052003c000700b9ff6eff45ff4bff6fff92ffa4ff;
    inBuf[9103] = 256'ha4ff9dffa4ffc3ffe8fffcfffdffebffd4ffc8ffc7ffc8ffd0ffe3ff0a003e00;
    inBuf[9104] = 256'h690079006f005900570077009a009e007a003500f8ffefff1a0050006a005500;
    inBuf[9105] = 256'h1900e2ffd5ffecfffbffe5ffb0ff78ff5cff6dff96ffb6ffb9ffb0ffbaffefff;
    inBuf[9106] = 256'h380066005d002400e3ffc3ffd7ff08002c002100f6ffdefffeff4f00ab00de00;
    inBuf[9107] = 256'hce009600650059006800720054000c00baff89ff8dffb4ffdcffecffe1ffd5ff;
    inBuf[9108] = 256'he8ff1300330032000700c2ff8fff8affaaffd1ffe1ffd2ffbaffbeffefff3f00;
    inBuf[9109] = 256'h8b00b000a10074004a003a00430055005900440022000900090023004a006800;
    inBuf[9110] = 256'h6b00550032001000fafff0ffe1ffc5ffa3ff88ff85ffa4ffd3fff8ff0a000e00;
    inBuf[9111] = 256'h1100220043005b004d001a00ddffbdffd1ff0a003e004b003100110017005400;
    inBuf[9112] = 256'hac00e800e000990041000b000a002e0043002100d8ff9bff98ffd5ff27005500;
    inBuf[9113] = 256'h48000e00d6ffcefff7ff25002900f5ffa8ff7bff94ffe1ff3000550041001900;
    inBuf[9114] = 256'h0e0034007a00b300b3007b003100ffff010032006a0082007000450022002100;
    inBuf[9115] = 256'h3d005b0063004a001500dbffb2ffaaffc2ffe2fff6fff5ffe6ffddffecff1700;
    inBuf[9116] = 256'h46005d0050002b000600f3fff6ff00000200fdfff9ff080036006b008b008e00;
    inBuf[9117] = 256'h7e00760085009f00a60083003d00f6ffdafff2ff220042003300ffffd0ffd0ff;
    inBuf[9118] = 256'h0a0050006a004100eeffa8ffa0ffd2ff0c001d00f2ffb0ff99ffcaff2a008300;
    inBuf[9119] = 256'h9a0069002100030029007700af00a4005c000700e6ff11006600aa00b0007700;
    inBuf[9120] = 256'h2600f6ff020038006a0069002e00dbff9eff95ffc1ff0800390039001700edff;
    inBuf[9121] = 256'hd5ffe5ff120037003c001c00e6ffbaffbaffe8ff29005b0064004c0031003100;
    inBuf[9122] = 256'h54008700ab00aa007e0047002a0031004c00600053002800fefff2ff0b003900;
    inBuf[9123] = 256'h53003f000b00d7ffc1ffd8ff080025001700e8ffbaffb1ffd4ff0c003b004300;
    inBuf[9124] = 256'h2500ffffedfffeff2a005600630051003300240033005a008100900080005b00;
    inBuf[9125] = 256'h37002200260037003d002d001200fdfff6ff02001a002e002c001f0013000800;
    inBuf[9126] = 256'hfffff8ffebffdbffd1ffcfffd8ffe9fff4fff8fffbff03001600330048004d00;
    inBuf[9127] = 256'h490041003b003d0046004a00450038002e0030003d00490049003f0032002600;
    inBuf[9128] = 256'h2400250021001300faffe2ffddffecfffeff0700fdffe4ffcfffd1ffe6ff0400;
    inBuf[9129] = 256'h19001400f6ffd2ffc0ffd2fffdff2c004900440023000300feff1c004e007200;
    inBuf[9130] = 256'h6b003b000100deffe7ff150049005e0047001a00f4fff0ff1500440055003900;
    inBuf[9131] = 256'h0300d0ffb8ffc6ffe7fffaffeeffcdffb0ffaeffcbfff4ff14001c000b00f3ff;
    inBuf[9132] = 256'hebfff2ff00000c000f000c000700020006001500250035004000400033001d00;
    inBuf[9133] = 256'h0900050010001d001d000500dfffcdffd9ffffff300048002d00f2ffc3ffbeff;
    inBuf[9134] = 256'hdfff0a001800f2ffa8ff6fff6fffaaff0300430042001000ddffcaffe6ff1c00;
    inBuf[9135] = 256'h41003a000300bcff95ffa0ffccff0600300039002c001c00160024003b004600;
    inBuf[9136] = 256'h41002500ecffafff89ff85ffa6ffd8fffbfffeffe8ffceffcdfff2ff22003200;
    inBuf[9137] = 256'h1600dbff9bff7cff93ffc4ffe4ffdeffbbff9fffb0ffeaff2c0050003f00feff;
    inBuf[9138] = 256'hbbffa8ffccffffff17000100c8ff9bffa5ffe5ff340062004e000800c4ffabff;
    inBuf[9139] = 256'hc6fff8ff0f00f3ffb4ff78ff68ff93ffd8ff0e001800f5ffc9ffb5ffbfffd7ff;
    inBuf[9140] = 256'he5ffd3ffabff8aff82ff96ffbaffd6ffdfffe1ffe9fffdff1b002e002000f5ff;
    inBuf[9141] = 256'hc6ffaeffb6ffd0ffe5ffe1ffc5ffabffb2ffdeff140035002a00f6ffbcffa4ff;
    inBuf[9142] = 256'hb6ffd5ffe0ffc5ff93ff6cff72ffa2ffdbfff8ffebffc4ffa8ffb1ffd2ffe5ff;
    inBuf[9143] = 256'hd4ffa4ff74ff6aff97ffdaff04000000d9ffb4ffb9ffefff2e0049002900d8ff;
    inBuf[9144] = 256'h8aff74ff9cffe4ff19001000d6ff9aff88ffb2ff01003e003900efff8dff4fff;
    inBuf[9145] = 256'h53ff8affccffe7ffc2ff7cff50ff61ffa9ff000028000400b7ff79ff74ffabff;
    inBuf[9146] = 256'hf1ff0700dcff92ff63ff79ffccff220041001200beff89ff98ffe0ff2a003900;
    inBuf[9147] = 256'h0000acff75ff7bffb9fffcff1100f2ffb7ff87ff7aff8fffb5ffd1ffceffb4ff;
    inBuf[9148] = 256'h96ff80ff7dff90ffacffc7ffd9ffd2ffb0ff8dff84ff9effcdfff9ff0100deff;
    inBuf[9149] = 256'haaff92ffa8ffe0ff17002100f5ffb9ff96ffa5ffdbff06000300d7ffa2ff8bff;
    inBuf[9150] = 256'ha6ffd6fff2ffe7ffbbff8fff86ffa5ffcdffd9ffc0ff97ff7cff85ffb1ffdcff;
    inBuf[9151] = 256'he3ffc5ff9eff8bff9affbfffdeffe3ffccffb0ffaaffbbffd6ffecffefffe4ff;
    inBuf[9152] = 256'hdeffe3ffebfff2fff0ffdeffc9ffc3ffcaffd0ffd0ffc6ffb6ffacffb0ffbcff;
    inBuf[9153] = 256'hcdffdaffd4ffbcffa4ff97ff9dffb3ffccffd7ffcdffb6ffa1ffa0ffbaffe1ff;
    inBuf[9154] = 256'hfeff0000e5ffbeffa7ffafffd4fffbff0700f7ffd8ffbfffc3ffe2ff03000f00;
    inBuf[9155] = 256'h0400e7ffcaffbeffc7ffd7ffe2ffdfffd1ffc3ffc0ffcbffd9ffe0ffdaffc9ff;
    inBuf[9156] = 256'hbbffb7ffb8ffbbffc1ffc4ffc2ffc2ffc8ffd6ffe5ffeffff4ffefffe3ffe0ff;
    inBuf[9157] = 256'hecfff7fffcfff8ffe8ffdaffd7ffddffefff03000800fffff0ffdeffd1ffd2ff;
    inBuf[9158] = 256'hddffe6ffe9ffe5ffdeffd7ffd3ffd5ffdfffeffffafffbfff2ffdfffcbffc5ff;
    inBuf[9159] = 256'hceffdfffeefff2ffedffe3ffddffe6fffeff110016000e00faffe7ffe1ffe2ff;
    inBuf[9160] = 256'he8fff3fffafffbfffeff03000400000002000c00170019000e00f6ffd8ffc8ff;
    inBuf[9161] = 256'hcfffeaff070012000500efffe3fff2ff14002f0031001b00f6ffdfffecff0900;
    inBuf[9162] = 256'h190017000400eefff4ff1600380042002b00ffffe1ffebff100030002a00ffff;
    inBuf[9163] = 256'hccffbbffdfff2400590057002500ecffdafffcff38005f0051001400d9ffcaff;
    inBuf[9164] = 256'hecff2500490041001e00030006002c0058005f003d001100f8ff030028004100;
    inBuf[9165] = 256'h37001300eeffebff12004500630056002400f7fff2ff10003b0054003f000d00;
    inBuf[9166] = 256'he6ffe0ffffff31005300550042002a0021002f00440051005100440035003100;
    inBuf[9167] = 256'h3100300034003a003e0044004d004c0040003100260020002600320035002900;
    inBuf[9168] = 256'h19000e000c0019003200470050004c00400032002d0032003e00490049004000;
    inBuf[9169] = 256'h32002b00330048005c00680068005e0059005f00660067005c00450032003200;
    inBuf[9170] = 256'h410055005e004e0030001f0029004a0070007a005d002900fdfff8ff23005900;
    inBuf[9171] = 256'h6e0054002400000007003e008300a800990066002f00220049008300a7009d00;
    inBuf[9172] = 256'h6a0038002a0046007d00a700a100780053004600560075007f00670040002000;
    inBuf[9173] = 256'h1b003b0061006b0054002f001a002c005a008000840061002c000f0023005500;
    inBuf[9174] = 256'h8200890067003f0032004c008300b300b900990071005c0064007f0097009800;
    inBuf[9175] = 256'h7d0061005b0069007a00850078005f005300550060006d006600460029002100;
    inBuf[9176] = 256'h2f004e0069006d005a003c002e003e0061008500960086006000430041006000;
    inBuf[9177] = 256'h9000b100b00092006b00570067008f00b200b4009400660049004d006a008700;
    inBuf[9178] = 256'h8d00760052003e0048005f006b00600043002c002e0044005d0061004b003100;
    inBuf[9179] = 256'h2a0044007200930091006e0046003c005d008c00aa00a2007b00560056007900;
    inBuf[9180] = 256'ha600bc00aa007c005800590074008d008c006b0042003100450069007c006900;
    inBuf[9181] = 256'h3b001700190040006e007c0058001c00f5fffeff36007c009e0086004c002000;
    inBuf[9182] = 256'h24005a009a00ba00a4006800330029004f008a00af00a500750042002f004400;
    inBuf[9183] = 256'h6e0089007e0055002900110016003100430039001c000500010012002d003c00;
    inBuf[9184] = 256'h2d000c00f6fff9ff16003e004d0037000f00f4fffcff2c0061007b006c003c00;
    inBuf[9185] = 256'h11000c002d005c007d0075004a001900010011003c005d005e003c000900edff;
    inBuf[9186] = 256'hf9ff170030002d000a00e5ffd6ffdffffbff150016000200ebffe3fff4ff1300;
    inBuf[9187] = 256'h24001b000000e7ffe7ff0100240038002e001000f5fff3ff0c002c003a003000;
    inBuf[9188] = 256'h1500f5ffe6fff0ff08001b001a000800f3ffe5ffe7fff5ff0700150018000b00;
    inBuf[9189] = 256'hf7ffebffebfff7ff0e002700300026001400050009001f0039004b004d003e00;
    inBuf[9190] = 256'h2a002100280038004c00570051004000300025001d001f002b0032002c002000;
    inBuf[9191] = 256'h11000100fbff060019002700230011000000f9ff01001800290028001d000f00;
    inBuf[9192] = 256'h0f002500410051005400430034003f0058006c0071005e003e0031003c005600;
    inBuf[9193] = 256'h7000730057002f0016001c003a005300550037000500deffd9ffedff08001300;
    inBuf[9194] = 256'h0200e3ffc8ffbcffc8ffe0fff3fff7ffebffd6ffc9ffc7ffd2ffe8fffbff0100;
    inBuf[9195] = 256'h0000fdfff5fff2fffcff0d001d0026002900230016000c000e0016001e002900;
    inBuf[9196] = 256'h2e0028001e0016000e000d001900220021001a000c00fbfff7fffbfffdfffdff;
    inBuf[9197] = 256'hf9ffeeffe5ffe2ffdfffdaffcfffc3ffbdffbcffbdffbaffacff94ff7bff72ff;
    inBuf[9198] = 256'h7fff92ff96ff87ff69ff4cff43ff53ff6dff7cff73ff59ff42ff3fff54ff75ff;
    inBuf[9199] = 256'h8dff92ff88ff7dff80ff95ffb0ffc4ffcdffd0ffd5ffe0fff3ff060010001500;
    inBuf[9200] = 256'h1f0029003600430044003e00380035003d004800430037002b001b0010001100;
    inBuf[9201] = 256'h12000d000100eeffdbffccffc0ffbcffbdffb8ffb2ffaaffa0ff97ff90ff8aff;
    inBuf[9202] = 256'h8aff91ff99ff9dff95ff83ff75ff74ff7dff8eff9eff9eff8dff76ff69ff6bff;
    inBuf[9203] = 256'h76ff7fff7eff6eff4eff2eff1fff21ff2cff2eff1dff00ffe2fec9fec0fec5fe;
    inBuf[9204] = 256'hc2feb4fea3fe8dfe7afe76fe77fe75fe74fe72fe72fe79fe82fe8dfe93fe8cfe;
    inBuf[9205] = 256'h88fe92fea5febdfed4fedafed6fed5fed9feeafe07ff21ff2fff2dff1eff15ff;
    inBuf[9206] = 256'h19ff27ff3cff4aff47ff3fff34ff28ff29ff32ff34ff32ff2aff19ff06fff9fe;
    inBuf[9207] = 256'hf2feeefeebfee5fedcfecffec5febffeb9feb5feb4feb1feaefeaefea9fe9efe;
    inBuf[9208] = 256'h95fe8ffe90fe9ffeb7fec4fec1feb6feaffeb8fed4fefafe18ff21ff19ff15ff;
    inBuf[9209] = 256'h1fff3fff70ff9affabffb1ffbaffcbffefff2000440054005d00650079009800;
    inBuf[9210] = 256'hb700c800c700c200cb00df00f200fe00f700df00cb00c400ca00d100c900ad00;
    inBuf[9211] = 256'h8a00690054004d00470039001b00f3ffcfffb8ffaaffa0ff93ff80ff6cff57ff;
    inBuf[9212] = 256'h42ff36ff33ff31ff31ff32ff34ff30ff29ff24ff21ff26ff35ff43ff4aff4cff;
    inBuf[9213] = 256'h47ff40ff47ff57ff65ff6bff66ff59ff4aff3aff33ff36ff32ff27ff1aff00ff;
    inBuf[9214] = 256'he1fed0fec4feb7feaafe92fe71fe50fe2ffe19fe08feedfdcffdb0fd8dfd75fd;
    inBuf[9215] = 256'h66fd4dfd34fd1afdf5fcd9fccafcb8fca5fc8cfc64fc3afc1ffc14fc18fc17fc;
    inBuf[9216] = 256'h00fcdbfbb3fb91fb8cfb9efbadfbacfb96fb71fb54fb50fb66fb8afba4fbabfb;
    inBuf[9217] = 256'ha7fba3fbaffbd7fb0afc39fc5efc75fc8afcb0fce5fc22fd64fd99fdbefde8fd;
    inBuf[9218] = 256'h1cfe5cfeaafef1fe23ff4bff73ffa1ffdfff23005b0081009500a700cb00fb00;
    inBuf[9219] = 256'h2c0154016701670163016b018201a101b701b701a30188017f018a019901a101;
    inBuf[9220] = 256'h97017e0168015b015c0168016b015f01540149014001480156015d0164016901;
    inBuf[9221] = 256'h72018901a301ba01d501eb0100022602520277029d02c102de0207033a036a03;
    inBuf[9222] = 256'ha103d80304042d0456048104b704eb0416053e055a0568058005a005bb05d705;
    inBuf[9223] = 256'hec05ef05ed05ee05f205fd050206f605e505cb05b005a905a705960584056f05;
    inBuf[9224] = 256'h55054a054b054f055c055e0555055e0576059605ca05fb0518063a0663069806;
    inBuf[9225] = 256'hee0649079707e7072b086508ba081d097b09d909230a570a900acc0a080b500b;
    inBuf[9226] = 256'h8a0ba80bc00bc80bc60bd30bdb0bce0bb70b8b0b4d0b110bd10a8d0a4c0afe09;
    inBuf[9227] = 256'ha5094c09ed0893084208ea0794074007e4068f064406fb05b80576053205f604;
    inBuf[9228] = 256'hc40498047e046b044a042e041004ed03de03d703c803b80391035a0332030503;
    inBuf[9229] = 256'hcd02a20264020902b0014d01dd007900050077ffe9fe4afea0fd07fd61fca5fb;
    inBuf[9230] = 256'heefa31fa6df9bff812f85ef7b4f601f648f5adf421f498f31ef3a5f228f2bff1;
    inBuf[9231] = 256'h69f129f1fff0d5f0aef095f07df074f089f0a2f0bff0e0f0f0f00bf13af163f1;
    inBuf[9232] = 256'h99f1d2f1eaf106f22cf235f250f27df27ff27af275f242f220f217f2e4f1b6f1;
    inBuf[9233] = 256'h8cf12bf1d3f097f03cf0f5efc0ef54efeeeea2ee35eee2edb8ed6bed1eede7ec;
    inBuf[9234] = 256'h98ec5fec51ec3bec32ec3dec2fec2bec4bec6feca6ecf6ec34ed6aedb4edfced;
    inBuf[9235] = 256'h4eeebfee30ef94eff9ef54f0aff01af18af1fef172f2cbf21cf377f3bff319f4;
    inBuf[9236] = 256'h79f4b7f4f5f42ef554f581f5c2f5e8f509f63af646f64df67cf698f6aff6d9f6;
    inBuf[9237] = 256'hdaf6d3f6f2f6fcf60ef73af735f724f72df713f707f71ff70af7e7f6d1f68af6;
    inBuf[9238] = 256'h47f621f6d6f584f52ff5a4f417f496f3f7f258f2aff1d9f000f022ef33ee52ed;
    inBuf[9239] = 256'h66ec65eb68ea5ae956e878e794e6c2e50be53fe494e321e3abe26ce26ae25ae2;
    inBuf[9240] = 256'h80e2e8e24ce305e413e51de67ae726e9c2eab3ecfdee3df1cff3acf66ef974fc;
    inBuf[9241] = 256'hbaffdd024106e0094f0de610a1141e18bb1b711fdd225226c729e22cf52ff932;
    inBuf[9242] = 256'ha0353538a43aa63c8c3e46409f41e642fb43a8443c45954593458f455745cd44;
    inBuf[9243] = 256'h40447643674274415140f43ec23d643cd53a8339183894365e350f34ab329e31;
    inBuf[9244] = 256'h8530622fa92eea2d1f2db92c472cce2bbc2ba32b7d2bb32bdd2bf72b5e2cb22c;
    inBuf[9245] = 256'hf32c792dea2d3b2ebc2e242f6a2fc82f013014302f301830d62f892f022f542e;
    inBuf[9246] = 256'h972d962c692b252a9f28f9263f2543232e21011f8f1c0f1a8117b414df11050f;
    inBuf[9247] = 256'hf20be708e505af028fff95fc7ef984f6c4f3faf056eefbebafe996e7d4e52ae4;
    inBuf[9248] = 256'hb0e292e197e0cbdf5fdf27df18df66dff4dface0b7e105e374e428e623e82fea;
    inBuf[9249] = 256'h5fecc6ee34f1abf33af6b8f826fb9efdf8ff2a025a0463062d08e709760bb50c;
    inBuf[9250] = 256'hdb0dd50e6c0fd90f2210fe0fa30f2b0f510e420d230ca90aff085b0774057303;
    inBuf[9251] = 256'h8e0177ff51fd5afb46f934f75ef578f39df102f061eed9ec95eb4dea2be93fe8;
    inBuf[9252] = 256'h59e79ae614e6a1e54ee535e51be516e53ee560e599e5f3e52ee666e6a7e6c0e6;
    inBuf[9253] = 256'hd3e6efe6e3e6c9e6a9e65ee60ce6bce552e5ebe483e4fbe375e3fae270e2ede1;
    inBuf[9254] = 256'h71e1dde04ce0c7df38dfb9de5adef3dd99dd69dd44dd43dd7fddcadd34decdde;
    inBuf[9255] = 256'h5fdf08e0e6e0b0e17ee26be32ee4f1e4d6e58ee64ee736e8e7e8a3e991ea46eb;
    inBuf[9256] = 256'h0fec06edaeed5cee29ef99ef16f0b0f0daf011f166f142f134f157f107f1d5f0;
    inBuf[9257] = 256'hddf075f028f00ff07eeffbeea5eed2edf8ec39ecf1ea8ce938e866e66fe484e2;
    inBuf[9258] = 256'h21e087ddf4da07d8ecd4e1d19ece27cbacc710c455c0a9bc06b950b59bb106ae;
    inBuf[9259] = 256'h74aafea6eba314a16a9e439c7d9a01994a983c989398c499b49bfd9d22a128a5;
    inBuf[9260] = 256'h87a9a5ae93b4afba5dc1dcc884d0a7d893e18ceac1f39cfd6e075311ad1bb925;
    inBuf[9261] = 256'h702f3b396a42fa4a6353025bbb610068586db771907582787e7add7b597ceb7b;
    inBuf[9262] = 256'hdc7a0a79747633733c6faa6a7a65c05fb55934535b4c7e45603e35377730d129;
    inBuf[9263] = 256'h6c23bf1d5d186d13670fd20bd408d8064b0545042d0477043f05e106e508600b;
    inBuf[9264] = 256'h8c0efc11cb151b1a8b1e3c232728f52cc7316c36ab3ab23e2c42fb445f47e348;
    inBuf[9265] = 256'h7d499649a948c04664440541a83ce7374132ba2bfa247f1d3915c90cb803f5f9;
    inBuf[9266] = 256'h51f0ade6efdcb4d3cccaebc18db9adb1f8a9cea25b9c4296c790488c63882f85;
    inBuf[9267] = 256'h2283c881fb80538171820c84cd86608a4c8e44931699339f52a654ae7db662bf;
    inBuf[9268] = 256'h03c9a1d2bcdc6ae7d0f138fcd006d110771a1724072d5c35733dbd44474b8a51;
    inBuf[9269] = 256'h2157fc5b7e604b6436679d694d6b1b6c5c6ce86b856a7768c66559626f5e2b5a;
    inBuf[9270] = 256'h805585505d4b1c46d940bf3be7363332b62d9829ab250322e51e101c7b196e17;
    inBuf[9271] = 256'h9e1510143013b8129d123f134b14a815b2171d1ad21c1a208623eb26782acf2d;
    inBuf[9272] = 256'he930f6338e36b338823aa03b373c763c073c283bf239f9378f35d5325b2f7f2b;
    inBuf[9273] = 256'h5e277222161d73171011550a81031afc8ef439edb0e556de94d709d1ffcaedc5;
    inBuf[9274] = 256'h75c1b9bd1abb2eb9eab7bdb74db869b97abb3abe5bc156c519ca52cf63d544dc;
    inBuf[9275] = 256'h7de356ebebf3c4fc0606bc0f4b19a422e02b8f34b13c6d44524b41516c56995a;
    inBuf[9276] = 256'hc65d49600a62e162f9625662dd60be5e1a5cb3587e54a74f064a9c43ca3c7a35;
    inBuf[9277] = 256'h862d4c25d51c1614a10b9b03cffba4f42dee24e8f0e2b9de25db66d882d611d5;
    inBuf[9278] = 256'h3dd424d485d47cd515d714d993dba8de3de261e606eb17f08df538fb16011d07;
    inBuf[9279] = 256'hf60c9812f317941c8d20f7235f26ed27d02893287927e2255a231b208e1c3918;
    inBuf[9280] = 256'h4a133a0e7d081c0289fb47f45cec50e4bfdbacd2c3c9f0c020b8b7afa7a7f59f;
    inBuf[9281] = 256'h0499d192588dd8885785ce824981b380f6800182cf836686a2897b8d05921097;
    inBuf[9282] = 256'h9a9ce0a2aea9f9b00cb98cc141ca8ad307dd49e6b2efddf830011a0956104316;
    inBuf[9283] = 256'h7a1be91fdf220c259226c1265f26aa25d1238721121f7e1b791760132d0e7808;
    inBuf[9284] = 256'had02c5fb67f426ed18e5eddc45d53ccd7bc5a8beebb7e2b11aada8a802a593a2;
    inBuf[9285] = 256'h72a0009f859e1c9e169ea79e079f9b9fa6a08da1a3a20fa453a5d0a6a7a875aa;
    inBuf[9286] = 256'h78ac94ae61b009b26ab347b4ccb4c3b4feb39cb280b0d5add8aa68a7c1a30da0;
    inBuf[9287] = 256'h209c77984d95629225909f8e4f8dbb8c0f8dbd8d358f8091e293dc96b39ada9e;
    inBuf[9288] = 256'he8a318aaadb033b802c17fca5ad5cae167ee13fbf707fe13421f2e2aec33a33c;
    inBuf[9289] = 256'hde440f4c95520f59e15e25643b69916d637124755178f47a317d7b7ef87eed7e;
    inBuf[9290] = 256'h117e887c4a7a0a7704734e6e0569a063f55dfd572252324c69465a419c3c3038;
    inBuf[9291] = 256'h6e34b5302a2d592aae27442572238121af1f8b1e981d271d931d2c1e2e1fee20;
    inBuf[9292] = 256'hea226d259128ae2be42e2a320635c5374e3a323cb73da83ec53e8a3ece3d673c;
    inBuf[9293] = 256'hc53aa338ea351b33ea2f382c6c2817240f1fca19f413660d960642ff3ef715ef;
    inBuf[9294] = 256'hcce643def6d5f6cd05c68cbec7b770b1c4ab01a7b3a2e49eef9b6b9957972696;
    inBuf[9295] = 256'h5d95d3941f95eb9517975799629ce19f6fa4d5a9b0af90b642be2ec6a5ce7fd7;
    inBuf[9296] = 256'h21e0d0e89af1f9f913020e0a6f115f18461fce25fa2b2e320238473d72423b47;
    inBuf[9297] = 256'h584b2f4f6f52b1545e5655574a57b35680555f53bf50b44d1e4a6946af42c63e;
    inBuf[9298] = 256'he63a1e375b33bb2f482ced2890252922c61e4c1bcc177d143511040e3c0bae08;
    inBuf[9299] = 256'h7906fd04e90341035703c3037d04d2054307b7086d0af00b480dbe0ef10fec10;
    inBuf[9300] = 256'he2117d12f3128513f3136214e014221557159215a015a2156c15ab148a13ff11;
    inBuf[9301] = 256'hf20fa70d0a0be7077504cd000cfd8ef95ff658f383f0e3ed77eb69e9d0e775e6;
    inBuf[9302] = 256'h20e5d1e378e228e134e090df05dfbddea3deb1de68dfd0e0a1e205e5c4e79cea;
    inBuf[9303] = 256'hf5edd2f1dbf523fa5bfe2502ce056f09e20c45106f1321169418ff1a791d1520;
    inBuf[9304] = 256'hb92231255a274d29272bcd2c2e2e292f612fed2e182ecd2c352b752932278824;
    inBuf[9305] = 256'hdb21141f651c041a8e17f0146212c40f360de70a8608f3054603690088fddcfa;
    inBuf[9306] = 256'h44f8aef531f3c8f097eeddec9aeba9ea08eaa7e972e981e9d7e942eaa8eaf6ea;
    inBuf[9307] = 256'h14eb25eb3beb48eb57eb56eb40eb51eb85ebd0eb51eccbec1fed84edcdedf3ed;
    inBuf[9308] = 256'h1feef5ed60eda1ec84eb2ceae6e859e791e5d4e3e0e1f6df66dedbdc6adb2bda;
    inBuf[9309] = 256'hcfd893d79dd6a1d5c5d4fdd3fad20ed24fd19bd03fd021d009d04dd0e5d0bbd1;
    inBuf[9310] = 256'h24d3ecd4d4d60cd964dbc2dd6be02be3d2e58de829eb88edf8ef62f296f4c6f6;
    inBuf[9311] = 256'hdcf8a1fa5cfc1afe85ffcd000002b60228038b036603ee025a021d0182ffeafd;
    inBuf[9312] = 256'hcafb73f943f795f4c5f148ef7aecc0e976e7d6e441e217e0a0dd4edb71d93cd7;
    inBuf[9313] = 256'h1dd563d363d19dcf50cecccc76cb7aca47c94ec8aec7e4c633c69dc5c4c4f7c3;
    inBuf[9314] = 256'h3fc35ec27cc179c038bfe0bd65bcdcba56b9a5b7e6b51eb431b277b0f1ae63ad;
    inBuf[9315] = 256'h19acfaaacaa903a9aba877a8c2a877a93eaa92ab91adedaf02b3ceb6d8ba6ebf;
    inBuf[9316] = 256'hbec462ca9ed096d7aede07e6f1edf0f535fe22070b10dc18fa21c92a4f33123c;
    inBuf[9317] = 256'h6344104c8953335a0e60b0659f6ad06ea4729375b07766795a7aa67a747a5079;
    inBuf[9318] = 256'h70770075d171436e4e6ab765e260aa5b1256b450404bae458240383bec355c31;
    inBuf[9319] = 256'hfe2cf128ca25c2220320331e941c611b221bf61a0d1be71bd81c2e1e4d208422;
    inBuf[9320] = 256'h08250d280e2b532ee4314835b738ff3bc73e6741a0434045a74673477c473247;
    inBuf[9321] = 256'h384687448e42e13f7a3ccb386934572f0b2a2824a61df916d60f1b083c0020f8;
    inBuf[9322] = 256'h8cefebe658de8dd5efccc9c4b9bc09b536aec7a7e6a1219ddd9819957b926590;
    inBuf[9323] = 256'hbd8e448e628ee58e9890f792c895de99c49e1aa491aac9b150b9bac1cccaf9d3;
    inBuf[9324] = 256'ha4ddade783f168fb7605260f8918e021ad2ae432f13a73424249e14ff6552a5b;
    inBuf[9325] = 256'h0460436487675d6a846c886de96d876d0c6c056a6267d763dc5f7c5b8a566751;
    inBuf[9326] = 256'h244ca9462441a83b2d36c030782b64265721691cd3175313010f330b8a072204;
    inBuf[9327] = 256'h6701eefeddfca1fbb0fa22fa5bfac6fa7efbdbfc35fea0ff6c01020387044906;
    inBuf[9328] = 256'hba07fe084b0a3a0b0e0cee0c7e0df00d460e3f0e1b0edd0d560db10cc60b690a;
    inBuf[9329] = 256'hd208f106bf046402bfffcafcb6f990f67bf39ef0efed6eeb2ae934e7a0e564e4;
    inBuf[9330] = 256'h87e3e9e25ae2fee1dee1dee136e2d8e280e372e4bfe53de73be9a8eb2eee02f1;
    inBuf[9331] = 256'h14f428f782fa0efe7a01e3043808490b460e2a11c51321163118e719671bc51c;
    inBuf[9332] = 256'h021e0e1fe71f982017218221eb211622fa21a321dc20cb1fa71e341d831bc119;
    inBuf[9333] = 256'hbf17af15d313fb113910a90e080d780b230ad10896077b063d05f803da02ba01;
    inBuf[9334] = 256'ha800b5ffa6fe85fd7afc6efb6dfa95f9bdf8e0f726f77bf6dcf56bf5fbf466f4;
    inBuf[9335] = 256'hc6f3fcf2f7f1e6f0a2ef0dee5dec84ea88e8b4e6e7e409e34ee18bdfbcdd24dc;
    inBuf[9336] = 256'h93daf0d866d7bad5e5d330d280d0d4ce50cdc9cb48caf7c8cac7e4c650c6ebc5;
    inBuf[9337] = 256'hd3c50ac681c667c79fc80dcad2cbbacdb1cffad161d4ccd684d94cdc09df17e2;
    inBuf[9338] = 256'h47e573e8f0eb7eefe1f26cf6f4f939fd8900c10387062b09a20b8f0d3e0fb710;
    inBuf[9339] = 256'h8b1105124912e7112e115710f10e510dbe0bb3097d076605d002040054fd21fa;
    inBuf[9340] = 256'hb8f67af3c6eff6eb75e8aee409e1ebddb5dabed75dd5f3d2ced031cf7fcd06cc;
    inBuf[9341] = 256'h04cbf3c918c99fc809c88dc749c7dcc67ec640c6cbc549c5c7c41dc47cc3efc2;
    inBuf[9342] = 256'h5bc2c7c11ec158c076bf5fbe2dbdc9bb08ba28b830b610b42eb287b0dcae8cad;
    inBuf[9343] = 256'h98accbab93abefab74ac78ad01afb7b018b34fb6ebb93cbe4fc394c864ce00d5;
    inBuf[9344] = 256'hcedb03e3d1ea90f288fa3003f20bfa149f1e212888313b3b90447d4d0056215d;
    inBuf[9345] = 256'h3063ee68cc6de471b675bc78077bf67c287ed07e1e7fa17e767d9f7bde789275;
    inBuf[9346] = 256'hbb713b6d74682e63695db957d451c94b1f464740593a0635ca2fe02af5264e23;
    inBuf[9347] = 256'h0920cd1de61b7f1a1e1aea19f319a61a501b3e1ce81dad1fc2216b242427372a;
    inBuf[9348] = 256'hd72d8a316d355c39e53c3a403743a045bb472e49ce49f9496749194880462a44;
    inBuf[9349] = 256'h03417d3d3b394c34392f9e295c23e31ce315480e9806a6fe39f6b1edf9e4d9db;
    inBuf[9350] = 256'hd3d216ca58c1f8b83cb1c4a9e1a20d9dce974093e18f1f8df38afd89b189de89;
    inBuf[9351] = 256'h228bfa8c218f4f923596819ad89ff3a56aacccb3fbbb7ec4b7cd8ad758e14feb;
    inBuf[9352] = 256'h7bf54dffd6084612181b4423352b92323739a73f8f459f4a664faf5317572b5a;
    inBuf[9353] = 256'hb25c2e5e225f735faf5e635d8d5bb45849555a519a4c80473b42933cd8363631;
    inBuf[9354] = 256'h872bf725b920c21b0b17a2127a0e670a7d06d90241ffd3fbccf8e4f542f348f1;
    inBuf[9355] = 256'hacef92ee4cee60eed0eee7ef2bf1a2f292f476f643f830fad6fb51fde8fe3f00;
    inBuf[9356] = 256'h6501750221039a0307043204490454041a04cb037a030903990209022101f0ff;
    inBuf[9357] = 256'h63fe78fc58faf6f74ff58cf2c0ef1cedd8ea0be9b9e7d0e643e611e625e68de6;
    inBuf[9358] = 256'h32e7cde764e802e991e968eaa8eb12edceeeddf001f38ef59bf8d3fb54ff0003;
    inBuf[9359] = 256'h8006180ae10d93114815de18fc1bcd1e6621a423a025482769282a29b929392a;
    inBuf[9360] = 256'hcb2a632bea2b492c6c2c6a2c342ca62bbe2a4c294027e3244022631f931cbc19;
    inBuf[9361] = 256'hd8163714d111a20fda0d370c850af6087007ed05a20462030802b8005fff03fe;
    inBuf[9362] = 256'hdcfcd3fbd1faf4f92bf979f817f8fef711f855f8b3f811f981f9ebf92cfa3dfa;
    inBuf[9363] = 256'hf7f949f95df835f7d0f55ff4d3f226f19bef31eed3ecb0eb9bea61e928e8d6e6;
    inBuf[9364] = 256'h49e5b0e3e4e1c8df94dd3fdbd3d895d676d475d2ccd067cf52ceb7cd69cd64cd;
    inBuf[9365] = 256'hb4cd2bced6cebccfb2d0cdd1fdd223d47ad5fad691d887dab0dce6de83e15fe4;
    inBuf[9366] = 256'h49e7a0ea21ee7ff117f5abf8e4fb22ff2d029d04d706cb08290a5e0b6e0cfd0c;
    inBuf[9367] = 256'h680dcd0dd00dc30dc30d520d9f0ccc0b5b0a7b086d06bb03980060fda5f9a5f5;
    inBuf[9368] = 256'hdbf1d7edc5e920e65ee2a3de67db1dd8e2d427d262cfbdcca2ca84c88fc615c5;
    inBuf[9369] = 256'h87c324c235c12dc060bf0abfa8be9bbe18bfa3bf96c003c261c3f0c49dc6e8c7;
    inBuf[9370] = 256'h0cc9f1c945ca57ca2ccaadc932c9aec80ec880c7dfc631c68fc5b9c4bbc392c2;
    inBuf[9371] = 256'hffc04cbf95bdb6bb19bac8b87db7a0b631b6dab5fab58ab62bb752b821ba51bc;
    inBuf[9372] = 256'h57bf49c3adc7c7ccb1d2e3d88fdfcbe6eded14f587fcd403470b5f139b1b1324;
    inBuf[9373] = 256'h222d2036063f2648b8508258cb5ff3650e6bb46f847398765f796c7be17c1f7e;
    inBuf[9374] = 256'hba7eae7e027e487cab7951762d72a96db8684763ce5d21585352ef4c7447c441;
    inBuf[9375] = 256'h523c82368630272be225f820161d87198716bb14591382129512a512d7129a13;
    inBuf[9376] = 256'h46142f15b3163c181d1a9d1c581fa1226a26282aee2d7131613410373e39c73a;
    inBuf[9377] = 256'hfb3b803c5a3cf63bfd3a7f39cd376b3561320b2ffa2a3c262c216e1b0c15750e;
    inBuf[9378] = 256'h7c071d00b0f80ef100e9d6e0aed854d01fc85bc0b1b864b1edaae8a47d9f389b;
    inBuf[9379] = 256'h8397519438929b905b8f278f778f2a9001929394af970a9c42a103a7dead8bb5;
    inBuf[9380] = 256'h99bd61c6adcff6d876e235ecc9f553ff05096b12701b6b24f02cc6346e3c8b43;
    inBuf[9381] = 256'hc549b74f1a557a597c5ddf602063ec6418661d669a656364f361d85e135b5856;
    inBuf[9382] = 256'h3751d04bf145fc3f063af833ff2d35289b22241dd317ba129d0d8808c30303ff;
    inBuf[9383] = 256'h71fa82f6d8f29bef55ed8ceb4eea17ea45ead3ea27ec96ed1cef25f115f3fdf4;
    inBuf[9384] = 256'h47f77bf9b6fb4efecb002d03a905de07dd09d90b8a0dfe0e491044111412e012;
    inBuf[9385] = 256'ha4136c14131568155315b914a1131a122310db0d5f0bd708870694040e03fa01;
    inBuf[9386] = 256'h2d01a10050000700c0ff55ff7efe65fd25fcd9fa04fabbf9cbf968fa62fb7afc;
    inBuf[9387] = 256'h09feeaffd301f303fc05bb07a409a30b9a0dd80f14121e1447166418541a3c1c;
    inBuf[9388] = 256'hd11df31ee91fc120aa21db2225246d25ab26bf27bf289b291e2a392abc29a228;
    inBuf[9389] = 256'h36278725b82307224d20921e191dc81ba51ac619ce189b175116c7140c135d11;
    inBuf[9390] = 256'h850f720d5d0b3c092007430579039f01deff2cfe8cfc48fb4ffa64f99af8d9f7;
    inBuf[9391] = 256'hf9f629f659f546f406f385f19aef94ed91eb77e984e7c6e520e4cee2cfe1e5e0;
    inBuf[9392] = 256'h17e03cdf1fdee4dc9cdb40daefd89cd734d6d0d488d374d2a2d104d198d04ad0;
    inBuf[9393] = 256'h1cd041d0b7d07ad1b0d22bd4d2d5d2d7efd9f7db17de05e098e132e3bae41fe6;
    inBuf[9394] = 256'hdce7d4e9d8eb5bee30f1fef312f71efaa1fcf9fe09017202b203ce045705ca05;
    inBuf[9395] = 256'h390633062b063406bf0528058e046f03340216019dff26fee9fc69fbeaf987f8;
    inBuf[9396] = 256'ha5f660f4e9f1ccee6beb28e8b7e470e192dec9db70d9aed71cd6e7d4fed3dad2;
    inBuf[9397] = 256'ha0d15ed0c9ce2ecdb8cb2ecae2c803c853c70ac72bc74cc78bc7fac750c8d4c8;
    inBuf[9398] = 256'haec98bca9ccbf2cc2ece84cffdd01cd2fbd294d37dd305d354d23ad121d028cf;
    inBuf[9399] = 256'h23ce75cd0fcdb2cc8dcc42cc7ecb65caa9c851c6bbc3bac0aabdf7ba54b824b6;
    inBuf[9400] = 256'ha5b449b375b24cb228b285b27fb369b4e6b51cb878bac1bd10c2a5c61ccc64d2;
    inBuf[9401] = 256'h91d823df2ae6eaecf0f38bfb4603a00be1148f1ec1282833be3c9e45424e1056;
    inBuf[9402] = 256'hc95ccc62c867b56b376f3972bc74487793796f7b3d7d897e087f067f117efe7b;
    inBuf[9403] = 256'h357982750771246cb7660c61485b38554a4f5c492343313d48373d31e62bde26;
    inBuf[9404] = 256'h0322331ecd1ab417c3151c149812f311231134100510b90fa40f9a10ba115b13;
    inBuf[9405] = 256'h0e16ec18431c3f20f923c827962bb32e9e3116349c35c9364a37f8369336b435;
    inBuf[9406] = 256'h5034ef32e1303d2e962b49289224dd206e1c69171d12020c60057dfe03f734ef;
    inBuf[9407] = 256'h4de741df4fd7a2cf52c85cc1c8bae5b492afb9aacca66da35ea02e9e6f9cf99a;
    inBuf[9408] = 256'h849a809ab19ad79b6b9d559f70a246a6b6aa5bb0aab674bd35c584cd1fd62fdf;
    inBuf[9409] = 256'h4de822f1b3f9fd01e8097111d8180220ae26482dad3377392e3f974428498b4d;
    inBuf[9410] = 256'h7f516a54f656d35865596d59b858e056ae54ed513e4e3c4ac045a940983b8e36;
    inBuf[9411] = 256'h9131dc2c4528d3236e1ff61aa7164012b40d70091005a100b5fcd3f82bf55ff2;
    inBuf[9412] = 256'hf6ef18ee4fedfdec16ed11ee3bef9df0b7f2dff40ef79bf9e3fbf9fd52008e02;
    inBuf[9413] = 256'hc50439078809bd0b200e9a1049134a166919821c6e1f0e2257243426a7279528;
    inBuf[9414] = 256'hdc28ab281a2827270c26cc244f23d7218420621f8d1ecb1dc51c561b70194817;
    inBuf[9415] = 256'h1515e012b010450e6c0b5e08300513026dff12fdecfa3cf9c3f787f6e5f582f5;
    inBuf[9416] = 256'h44f577f5c4f51ff6cdf659f79bf7d2f7cbf7c1f739f826f98ffa80fcaafe1101;
    inBuf[9417] = 256'hc803b806e609200d2410e2122415fa169618d619e81afb1bc21c6d1d211e691e;
    inBuf[9418] = 256'h6f1e681eee1d481db51cb51b6c1a0f1934171a1500136610510de009a805e400;
    inBuf[9419] = 256'h0cfc07f71cf2a6ed6ee97ce50ee2e8def2db45d996d6bcd3e1d0e5cdb7ca83c7;
    inBuf[9420] = 256'h69c474c1f8be38bd1abca5bbb0bbe7bb38bcabbc52bd56bebebf77c166c368c5;
    inBuf[9421] = 256'h80c7aec9dccb24ce67d06fd26ad44fd6fcd7d5d9e8db12deb1e0aee3a6e6c6e9;
    inBuf[9422] = 256'hb7ecf3eebef004f28cf2e3f21af3f8f2fff22df337f38af30ef454f49cf4bdf4;
    inBuf[9423] = 256'h4bf4a9f3eaf2c6f1a1f094ef5bee46ed65ec65eb7eeab0e992e858e71fe6a4e4;
    inBuf[9424] = 256'h3ae31ee214e171e064e086e0e8e07be1aee199e15ae1a5e0e1df46df77dec5dd;
    inBuf[9425] = 256'h53ddcedcacdc15dd96dd6fde7fdf18e07de0b2e043e0addf12df1fde6cdd0edd;
    inBuf[9426] = 256'h8bdc49dc33dcbadb5ddb39dbe5dadcda12dbf9daf2da02dbc7dac8da12db24db;
    inBuf[9427] = 256'h41db55dbf3da84da2bda9fd93ad90ad9c8d8bbd8dcd8dfd8e9d8cfd841d882d7;
    inBuf[9428] = 256'h8bd654d533d4ffd2aad162d0f6ce7acd1bcc8bcae1c840c75cc59ec35bc239c1;
    inBuf[9429] = 256'h9cc0a9c0bbc036c150c264c3d1c4a0c60cc895c98ecb90cd67d06bd4fad886de;
    inBuf[9430] = 256'h16e5e0eb2bf3ecfa6102cb093f113f18351f6626812dd334853c2a44da4b9a53;
    inBuf[9431] = 256'hdc5a7e618667926ca1700874ad76b0786b7ab47b8a7c247d2f7d7c7c1f7bcb78;
    inBuf[9432] = 256'h7c757371a26c4967a961bc5be1552e50824a2945f13f9c3a83355b30102b2f26;
    inBuf[9433] = 256'h45214f1c091803146e10240e770c590b4c0b560b710b480c150d130ed70f8611;
    inBuf[9434] = 256'h5913c115f017391af01c5a1fcd216b249e26c528be2a042cf32c532df52c6a2c;
    inBuf[9435] = 256'h6c2bd029f7275c25f921511e071a40157b10470ba705ecffcdf956f3c9ec2fe6;
    inBuf[9436] = 256'h78dfd6d883d24fcc49c6abc03bbbe0b519b1b6ac91a84da59ea243a0009f7e9e;
    inBuf[9437] = 256'h759eb69fc6a12ea4aba7bbabe5afe8b459bab7bfacc5fbcb4dd24ad9dde093e8;
    inBuf[9438] = 256'habf00ff94a017309b511b6194e21be28b82f0336203cd241af46354b254f0452;
    inBuf[9439] = 256'h86549b56be578c58e25833582157b955a8536951e44ec34b51487c442a40923b;
    inBuf[9440] = 256'ha4366f31052c80264121281c26179812150e9409ba052402cdfe54fc10faedf7;
    inBuf[9441] = 256'h9af670f56ef446f43cf44df430f53af65af713f9bbfa5ffcaefe60019904b108;
    inBuf[9442] = 256'h010d3d1166150d193b1c251fa621c52391250e277228e129672b042d8b2ef62f;
    inBuf[9443] = 256'h46314f32fa320a3320324430c12ded2a3628d4259a234321b71ef41b0a193816;
    inBuf[9444] = 256'h731389107a0d600a4a0774041e0204000bfe5cfcb3fa12f9bbf74af699f4fdf2;
    inBuf[9445] = 256'h60f10cf0a8ef01f0ecf08bf265f44cf680f8b0faacfc80fedfffe400f8013503;
    inBuf[9446] = 256'hcc04cc06ec08210b610d9c0fec111614e81563174618b41806190919de18c518;
    inBuf[9447] = 256'h5c18c41737171f16781473129f0f510c2109d2059e02c5ffbefca0f9aef68af3;
    inBuf[9448] = 256'h50f032edcae91de65ae24bde19da11d63dd2ddce32cc3ccae6c806c85fc7c2c6;
    inBuf[9449] = 256'h2ac6b9c57ec57cc5bcc515c66ec6f5c6bac7c1c828cadacbb3cdbacfe6d12dd4;
    inBuf[9450] = 256'h96d61cd9b2db52de08e1d7e396e635e98eeb62edddee24f01ff120f23ff333f4;
    inBuf[9451] = 256'h49f597f6cbf737f9cffaf2fbd8fc89fd9dfd9efdc1fda3fda2fdb3fd5efd1cfd;
    inBuf[9452] = 256'hfbfca0fc77fc64fcecfb68fbd9fa07fa6bf918f9e4f820f9aaf924fa95fab3fa;
    inBuf[9453] = 256'h3ffa72f956f803f7c8f5b0f4b4f3f5f271f218f2fcf120f251f26af261f2f7f1;
    inBuf[9454] = 256'h0df1d0ef40ee87ec17ebf7e92ae9dde8a1e829e891e790e64ae53ae431e344e2;
    inBuf[9455] = 256'hb2e110e18ae085e0a6e01ce100e29fe2fde222e392e2bee1f1e0dcdf20df03df;
    inBuf[9456] = 256'h31df1fe0b5e146e3f4e483e670e730e8bfe8bce880e8ede7c4e680e547e420e3;
    inBuf[9457] = 256'h5fe2d6e14de1bde0e9dfe9dedddda2dc5cdbf9d946d89ad6f5d43dd3d7d189d0;
    inBuf[9458] = 256'h12cfdecdbfcc9bcb0dcbceca87cab3ca21cbafcb25cd83cf79d26bd60fdbd8df;
    inBuf[9459] = 256'h22e5dcea86f061f659fcd9014407000dc7120e194120d727e62fac387b41404a;
    inBuf[9460] = 256'h1a532d5b4862b168cc6da971ec7477777179337b7c7c797d6c7e037f317fd57e;
    inBuf[9461] = 256'h917d7c7b8c78c57474706d6bc665e15f7a59da52844c0946a53fae396f33322d;
    inBuf[9462] = 256'h75279421051c4f17c012c70ed00b0d09df0687052e042b03a902f40184019501;
    inBuf[9463] = 256'ha20126024d03b404d406b209e20c92106114c817d81a3c1dda1e0b209a208a20;
    inBuf[9464] = 256'h25202e1fc51d441c7c1a9418c416a4141712300f950b4107760221fd4cf742f1;
    inBuf[9465] = 256'h10eba7e43aded6d73fd1aaca62c43cbe6ab845b374ae06aa6fa66ba323a119a0;
    inBuf[9466] = 256'hda9f28a046a1aaa21aa413a660a8e2aa29ae26b29fb608bc69c26dc950d111da;
    inBuf[9467] = 256'h27e385ec2bf678ff4f08ec10dc181d203527c52db933ab393d3f40445a49264e;
    inBuf[9468] = 256'h4d525456cf59525c515e835f995f0c5fbb5d6b5b7858dc547850984b5e46e040;
    inBuf[9469] = 256'h523be635af309c2bcb264422b41d3a19f5147410d80b5f078b02a4fd2ff9def4;
    inBuf[9470] = 256'h22f190eeafeca1ebb3eb3eec45ed11ef19f163f329f6e3f88ffb68fe1f01ce03;
    inBuf[9471] = 256'hb7069a09750c640f3812e7148017ef19361c601e6d2059221324872597262127;
    inBuf[9472] = 256'h2327a1268925df239a21a41e051bed168612080eb3099d05be012efeeffae3f7;
    inBuf[9473] = 256'h2af5c7f279f03fee0ceca1e922e7b5e449e228e086de49dd9edc94dcf4dcd4dd;
    inBuf[9474] = 256'h3bdf01e130e3bfe584e877eb81ee97f1bcf4dcf707fb38fe3e012c04ea063409;
    inBuf[9475] = 256'h340bee0c380e630f7f1057112a12ec124d138a139f133a1386127311aa0f5b0d;
    inBuf[9476] = 256'ha50a6407eb037700e8fc69f921f6e2f2b1efa4ec85e944e605e3b8df66dc52d9;
    inBuf[9477] = 256'h79d6e0d3c5d120d0e8ce46ce0cce08ce4cceafce23cfd6cfbad0c6d10ad35fd4;
    inBuf[9478] = 256'hced577d74ad969dbcfdd3be0b2e214e529e723e902eba0ec3feec5effcf024f2;
    inBuf[9479] = 256'h1df3b4f336f485f47af460f41cf48ef307f372f2b7f120f1a0f01bf0c1ef73ef;
    inBuf[9480] = 256'hfdee73eec4ede4ec0eec5debc7ea6cea56ea6eeacbea84eb73ec8fedcaeed6ef;
    inBuf[9481] = 256'hb2f082f12af2d9f2baf38ff46ef575f65cf74ff868f947fa06fbb1fbf1fb15fc;
    inBuf[9482] = 256'h4dfc52fc6ffcacfca4fc9afc8efc19fc78fb99fa26f97cf7b8f5bdf3f6f162f0;
    inBuf[9483] = 256'hc2ee4cedeeeb83ea47e92ee808e7eae5b8e463e31de2f4e0ebdf1edf89de0ade;
    inBuf[9484] = 256'h98dd3eddf4dcc5dccfdcfcdc47ddcddd65de10dff4dfd5e0b5e1c1e2b1e39be4;
    inBuf[9485] = 256'hafe585e63ae7fee767e8c7e868e9cae92feaa9ea88ea2deadde921e991e855e8;
    inBuf[9486] = 256'hbce72ee7b2e6bfe5f6e47be4c6e340e3bee2ade17be01edf50dd82dba4d992d7;
    inBuf[9487] = 256'haed5ecd351d212d1f5cf05cf51cea0cd2acdd3cc38cc90cbabca5ac948c877c7;
    inBuf[9488] = 256'hb5c695c6d4c617c7f3c72ac96bca44cc57ce3fd098d252d54bd830dceae005e6;
    inBuf[9489] = 256'hcbeb0cf23af888fedb04a20a091052154c1a711f5225a82b8a32353a0742ca49;
    inBuf[9490] = 256'h9b51bc58d45e15640c68d96a2a6df36e6770e6711973f1739074a87446746973;
    inBuf[9491] = 256'hd371ad6fea6c8869ec65e961815d16593954f74ec3490244ca3da9371431772a;
    inBuf[9492] = 256'hbb24621fca1a8817ad144b12d710660f230e770d710c330b270ab20848078806;
    inBuf[9493] = 256'h11064b0686074d09ce0b140f9e126e16541ae21d2521f2231e26d027d9282d29;
    inBuf[9494] = 256'hfd282128b126ec24b4222b20921dd51a091857158912730f0b0c22088f037afe;
    inBuf[9495] = 256'h06f922f308edfee6dbe0d6da56d522d05acb63c7cdc38cc00fbee6bb17ba3fb9;
    inBuf[9496] = 256'h03b952b9b2baa5bce1bed3c109c541c8ffcb13d054d44ed9eedee9e48debbaf2;
    inBuf[9497] = 256'hfdf97e014409da104818941f32260c2c6b311136293a473e3542e745b4493a4d;
    inBuf[9498] = 256'h49503553ae557857cd585859ea58c557ca55fb52974f9f4b35478f42c83d0e39;
    inBuf[9499] = 256'h5b34ad2f312bc5268e22ea1e991b9d182816ac131c11c50e2e0c6e09f4065204;
    inBuf[9500] = 256'hc601e6ff68fe89fdb8fd71febbffdc015b044307b90a290e6b11811404171319;
    inBuf[9501] = 256'hed1a761cdf1d401f6d207d216b2212238623b52386231123442206216c1f601d;
    inBuf[9502] = 256'he11a2b1861159712fc0f7e0dde0a0b08f1046a01a3fdd0f9ebf528f2c1ee99eb;
    inBuf[9503] = 256'hcfe892e6a8e415e3f8e110e15de006e0d3dfcbdf27e0cbe0dde198e3e0e5abe8;
    inBuf[9504] = 256'he6eb3eef7cf276f50ef84efa46fc21fe0900f8010c0450069208ea0a5b0d910f;
    inBuf[9505] = 256'h93114e135b14de14f6146d148f1386120a114f0f750d350bc00830063603f6ff;
    inBuf[9506] = 256'h9afc0ef9a5f5a7f2ffefbdeddaeb0dea43e87de69de4a7e2b4e0c7def6dc6edb;
    inBuf[9507] = 256'h47da8dd954d998d952da86db23dd08df07e1e1e272e4b5e5b8e6b9e7e6e841ea;
    inBuf[9508] = 256'hddeba4ed66ef37f112f3d2f496f649f8aff9f1fa07fcc1fc56fdb3fda0fd5efd;
    inBuf[9509] = 256'hf5fc4dfcbafb36fb85fad5f916f926f85af7c1f63af6edf5b6f54ef5d0f42df4;
    inBuf[9510] = 256'h4af35cf26ff172f099eff2ee68ee1fee1cee44eeb7ee8cefa3f008f2abf336f5;
    inBuf[9511] = 256'h91f6baf781f814f9b8f954fa12fb0ffcf8fcccfd96fe02ff30ff59ff45ff2dff;
    inBuf[9512] = 256'h41ff23ffe6fe99fed9fdcffca7fb13fa3ff841f6c6f309f148ee6eebdde8cee6;
    inBuf[9513] = 256'h0ae5a4e388e255e10ee0b6de23dd8cdb1edad3d8dbd750d708d70cd75dd7d0d7;
    inBuf[9514] = 256'h70d850d944da52db8adcbaddfade67e0cde138e3b4e4eee5fee613e8f8e8ebe9;
    inBuf[9515] = 256'h20eb36ec50ed80ee4eeff5ef9ef0d2f0ddf0e0f05cf0aeef04efededdcecf6eb;
    inBuf[9516] = 256'hbeea9ae99be844e707e6fbe4c7e3e5e261e2dce198e15ce1b3e0c5df6fde98dc;
    inBuf[9517] = 256'haadab8d8e4d674d548d474d30ad3d9d211d3a9d349d419d5e2d541d693d6c4d6;
    inBuf[9518] = 256'h9fd6b8d602d740d70ed847d98fda61dc74de4fe075e2cee413e7e7e94dede9f0;
    inBuf[9519] = 256'h38f52ffa57fff804ed0a8210c715b81af01edf220527402beb2f6235423b9941;
    inBuf[9520] = 256'h9948ab4f8356045d76629f66c269ca6b036def6d896ee66e296f206fc56e0d6e;
    inBuf[9521] = 256'hc96c006b936882650662f85d6d59a6544f4f9749e843e83dca37e2318d2bf924;
    inBuf[9522] = 256'ha91e381834124d0df80874050e03f40051ff71fe95fde9fca7fc2bfcc1fbc8fb;
    inBuf[9523] = 256'he5fb80fcddfd9bfff801fb043508b70b470f7a126715ec17fb19e11b801dca1e;
    inBuf[9524] = 256'hde1f6c206220eb1fcb1e161d051b6a1863153012b60e0c0b600788036aff06fb;
    inBuf[9525] = 256'h31f6c2f0d7ea9be421debdd7d3d15ecc7ec77bc316c041bd41bbb7b970b8b3b7;
    inBuf[9526] = 256'h21b797b690b6e0b66db7beb8abba06bd4ec068c400c963ce56d45edab2e048e7;
    inBuf[9527] = 256'hc8ed7df487fb83029009c810aa17281e6324df298d2ebc322136ca38343b423d;
    inBuf[9528] = 256'h063f04411443124533470c49374abc4a464aa7482146c342c63e8f3a5b366132;
    inBuf[9529] = 256'hbd2e6f2b7b28b7251923b1203a1ea51b111937164013a3103e0e4f0c2e0b680a;
    inBuf[9530] = 256'hf009f509f209f0093b0a6b0aac0a6b0b600cbc0dc20fee1127146e164518b819;
    inBuf[9531] = 256'hed1a9c1bef1b151ced1bc81bdf1b111c791cf61c2c1d1f1dae1ca61b231a0718;
    inBuf[9532] = 256'h2a15ce11180e300a84062b03050021fd53fa6cf790f4b7f1c6eee1eb0ee94de6;
    inBuf[9533] = 256'he9e30ce2b6e0fcdfc2dfcbdf03e049e06fe06be02fe0c1df66df6cdf2ee0ede1;
    inBuf[9534] = 256'h9ce40fe8ecebbaef44f35df6cdf8adfa0bfcd2fc51fdbafd07fe7bfe1fffaaff;
    inBuf[9535] = 256'h3b00cc001301320125019800b1ff8efe0ffd7efb03fa64f8b3f6eaf4c5f267f0;
    inBuf[9536] = 256'hf2ed4eebade842e60ee44be22be19ae092e0f8e085e122e2c2e240e395e3afe3;
    inBuf[9537] = 256'h68e3cde20ae255e111e188e1cae2eae4bee7ecea48ee83f13af461f6e6f7b3f8;
    inBuf[9538] = 256'h1af948f93ff948f972f99ff915fae0fac9fbebfc11fecdfe27ff12ff75feaafd;
    inBuf[9539] = 256'hdefcf9fb23fb46fa15f9a3f7fdf517f442f2b7f070ef86eeeced63ede1ec6cec;
    inBuf[9540] = 256'hf5eb9eeb86eb8ceba8ebd2ebdcebcdebcdebd9eb11eca2ec6aed6beeb1eff9f0;
    inBuf[9541] = 256'h46f2b1f304f55cf6ddf73cf97dfaa5fb56fcacfcdbfcb3fc78fc58fcf0fb53fb;
    inBuf[9542] = 256'h89fa36f9a1f714f666f4e8f2b0f154f0e3ee54ed54eb25e9eae679e409e2a6df;
    inBuf[9543] = 256'h1cdda3da56d830d675d43ad360d200d2fed129d282d2f1d255d3c5d34bd4e8d4;
    inBuf[9544] = 256'hc6d5f0d655d808da05dc2dde91e027e3ade51ee865ea45ece6ed6fefbdf00af2;
    inBuf[9545] = 256'h70f39df4bff5eaf6bef76bf8fbf8f0f885f8daf797f633f5f0f375f22cf12cf0;
    inBuf[9546] = 256'hfaeee0eddaec68ebdbe942e851e683e4f7e26de136e047df5edecedd9addabdd;
    inBuf[9547] = 256'h2bdedade70dfe1dff2dfc7dfa2df89dfc2df4ce0e0e0a7e188e24be350e475e5;
    inBuf[9548] = 256'h67e673e758e8c7e835e980e970e99de9f1e940ea1feb5bec82ede4ee3af03cf1;
    inBuf[9549] = 256'h95f279f4d1f61dfa2afe5d02cf06540b830faf13f217f81b032045248128042d;
    inBuf[9550] = 256'h11325c37033d24435a49944fc5555b5b1f600764cb669868b969336a396ae869;
    inBuf[9551] = 256'h2d693268fa668465f7631d62e45f645d455a81564152194d2f47f7403b3a7233;
    inBuf[9552] = 256'h332d12273f210b1cd216d611960d8c0906066303f100e3fe90fd5dfc81fb49fb;
    inBuf[9553] = 256'h19fb1ffb9ffb25fceafc1efe53ffbe009302a7045107af0a720e7e127516e119;
    inBuf[9554] = 256'hb41cc81e1a20ed203a210a218d20a01f3f1e8b1c601ac617f414e911b90e910b;
    inBuf[9555] = 256'h5408e104440178fd6af941f511f1a9ec02e836e322def1d815d48fcf81cb57c8;
    inBuf[9556] = 256'hdfc50bc439c327c39bc3ecc4d2c604c9e9cb4bcfccd2b6d6c9daa0deade207e7;
    inBuf[9557] = 256'h82eba1f074f689fc13030b0afb100b18451f2426a22cba32f637693c4c406943;
    inBuf[9558] = 256'he8451448c449174b4c4c3f4dec4d644e6d4eee4de54c314be14800469842d33e;
    inBuf[9559] = 256'hb13a4136b431fe2c4f2803240f20981cd91974175615b0132912c710d60ff30e;
    inBuf[9560] = 256'h160e890df10c660c4d0c5b0ca80c9f0d0e0f1c1113148417261bd61e0922b024;
    inBuf[9561] = 256'h0427e028612a962b2c2c312cca2bfc2a1b2a4a295d28632737269b24b5227720;
    inBuf[9562] = 256'haf1d901a0d170613bf0e2f0a2905e5ff67fab3f449ef71ea37e6dfe252e03ade;
    inBuf[9563] = 256'h97dc51db35da5bd9bfd82ed8b2d74fd7f9d6dbd620d7d3d70bd9ccda08ddb2df;
    inBuf[9564] = 256'hb8e212e6a6e94fed01f19bf4f0f708fbd0fd1900f2014c03fd033e042704a303;
    inBuf[9565] = 256'hf702360235012e0036ff1efe0bfdfafb98fafdf838f723f5f9f2dbf08fee26ec;
    inBuf[9566] = 256'h9fe9d1e6f5e34de1e7de01ddafdbc1da34dafdd905da75da63dbbadc79de6be0;
    inBuf[9567] = 256'h45e2fce381e5cbe611e85be99eea03ec8bed2cef14f13af36ef5c6f72efa80fc;
    inBuf[9568] = 256'hd8fe1401db0215049b04480481039c02a201bc00cdff6dfeadfcc0fab8f800f7;
    inBuf[9569] = 256'hd6f5fcf46bf40af485f3e0f221f202f189efcdedb0eb75e962e766e5aae352e2;
    inBuf[9570] = 256'h44e1c3e00ce100e2a5e3c9e5e0e7c8e977ebc4ecfeed56ef96f0d6f10ff3f3f3;
    inBuf[9571] = 256'hb0f465f5d9f53ff6a7f6d1f6f9f64df790f7e8f74ef859f81ff8baf7f8f613f6;
    inBuf[9572] = 256'h1ff5c8f316f219f0abed18eba9e84ae61ce41ee215e011de20dc2fda64d8ccd6;
    inBuf[9573] = 256'h58d536d47dd32bd35cd3f4d3c2d4cbd5ffd65fd81fda23dc2cde20e0b1e1bbe2;
    inBuf[9574] = 256'h93e377e498e559e7abe94aec44ef71f290f5d1f812fceafe65015d037704f404;
    inBuf[9575] = 256'hf00437042c030902a90078ff9bfea6fdb3fca8fb0ffa37f86af686f4f1f2c7f1;
    inBuf[9576] = 256'h97f06def35ee8becaceab3e86de622e4f8e1d9df29de20ddbfdc3edd79de1be0;
    inBuf[9577] = 256'hfee1cce34de58be672e70de877e89ee8b0e8d2e802e984e952ea29eb1dec01ed;
    inBuf[9578] = 256'h92ed19ee87eeb2eef3ee29ef1eef35ef47ef11eff1eebeee3beee6edb0ed60ed;
    inBuf[9579] = 256'h5bed79ed7aedebedfceeabf08df391f729fc4c019e068d0b4810e4142419501d;
    inBuf[9580] = 256'h872186258829cd2d2c32e8363e3cef41f5474a4e6e540c5afa5ed76295656967;
    inBuf[9581] = 256'h6968c2689b68ed67ae66e364a66221605b5d745a6157c5539d4ff64a9745d63f;
    inBuf[9582] = 256'h063aeb33c72dcc278521341b2a15000f1909d703c5fe36fa87f63af39cf0fbee;
    inBuf[9583] = 256'hc5ed26ed41ed72edd9ed98ee2aefcfefc0f0b2f106f3f2f439f718fa7afd0601;
    inBuf[9584] = 256'hd1049f08190c480fda118e139814e31491140e1444132712d310ec0e5e0c6909;
    inBuf[9585] = 256'hfc053b026ffe83fa75f666f247ee11ead9e599e137ddb3d826d48ccff4cab3c6;
    inBuf[9586] = 256'hdac27cbf09bd8cbbe4ba5abbb1bc6fbebfc06ac30ec616c986cc0bd016d4a5d8;
    inBuf[9587] = 256'h55dd91e26ae875eefcf4f1fbc40299097810fa16541da0237029c72eb233d837;
    inBuf[9588] = 256'h503b573ec0409b421344fb445c456d4527459744e7430043d3416140873e2c3c;
    inBuf[9589] = 256'h4839d335f231cc2d95299a25e021631e441b59189f1562138511ff0f060f460e;
    inBuf[9590] = 256'h970d4e0d400d7a0d680ec00f4a1134130d15ab166718001a711b1b1dc11e6d20;
    inBuf[9591] = 256'h8122b92404277a29972b362d712ef72eec2e812e712de42b092ab8274b25ea22;
    inBuf[9592] = 256'h5120a71dd41a8a171914a2100a0da5096b061303d8ffb4fc7ef97df6a1f3b1f0;
    inBuf[9593] = 256'he4ed3debb9e8b5e64ee571e43be487e421e510e63ce78fe81cead6ebaceda8ef;
    inBuf[9594] = 256'hb5f1bbf3aff573f701f96afab8fb0efd8bfe15009c0109032304e3045d057e05;
    inBuf[9595] = 256'h5705f3042104e4025b0175ff5ffd4bfb15f9bef658f4b9f1feee5fecc9e95ce7;
    inBuf[9596] = 256'h59e58fe3e2e162e0d2de3eddbddb2bdac3d8bdd716d704d785d751d870d9ccda;
    inBuf[9597] = 256'h31dcd5ddc3dfc7e1fde34ae669e878ea70ec29eed4ef6df1c9f21bf465f585f6;
    inBuf[9598] = 256'hb3f7eaf8f0f9ddfa99fbe1fbdbfb8bfbcafad0f9a5f814f745f54af305f1c1ee;
    inBuf[9599] = 256'hadecb7ea23e9f8e7f3e632e695e5c6e4f3e320e31be244e1b5e033e0f9dffddf;
    inBuf[9600] = 256'hf8df39e0c9e077e192e2fee360e5fde6c4e871ea5aec68ee2ef0d4f12ff3edf3;
    inBuf[9601] = 256'h68f4baf4caf404f57df507f6d9f6d6f7a0f848f9acf995f948f9ddf83ef8a2f7;
    inBuf[9602] = 256'hfdf603f6c7f44df375f177ef80ed95ebf1e9b3e8cce752e729e710e707e7ede6;
    inBuf[9603] = 256'h85e6f5e546e557e474e3cfe256e243e2ace247e310e4f6e4d0e5b8e69be79ce8;
    inBuf[9604] = 256'hbce903eb83ec31ee23f006f2e1f38cf5a5f674f70cf825f830f850f820f801f8;
    inBuf[9605] = 256'h1cf803f802f836f81ff8f1f7c6f72af757f66af5fdf34bf27af042eefbebe6e9;
    inBuf[9606] = 256'hd0e7fee597e462e38ce21ce2c3e187e14ee1cae01fe06cdfb5de4ade46de82de;
    inBuf[9607] = 256'h14dfe6dfc4e0d5e116e350e494e5cee6cae7bae8c7e9edea5dec0eeeb5ef35f1;
    inBuf[9608] = 256'h6af218f33df3daf2e9f181f0daee3dedceeba9eaf6e978e9f2e88de806e81fe7;
    inBuf[9609] = 256'h1de6c2e4e2e216e160dfc2dd0fdd1edd78dd9ade13e040e1c9e2a1e477e626e9;
    inBuf[9610] = 256'hbfeccff0f6f515fc8002970931118c18da1f0d27852d84334f39ad3e0444d749;
    inBuf[9611] = 256'hfc4f8c56ae5dd064776b807158769e79987b417c8b7be4796a770b7424700b6c;
    inBuf[9612] = 256'hc66789635f5feb5af9555a50fa49d5421f3b3d332f2b1623651bed13ab0c1106;
    inBuf[9613] = 256'hb9ff95f93cf45bef10eb10e8eae5a1e4c2e4aae558e73cea91ed32f14bf504f9;
    inBuf[9614] = 256'h5efcacff98029f052a09fb0c72117b16a51b2921a426ab2b723066343c374b39;
    inBuf[9615] = 256'h203ac939d138d7360a34de30dd2c39285623d31d06185c12920cec06a0015ffc;
    inBuf[9616] = 256'h21f7caf11dec13e6abdf21d9a5d25dccd1c61fc245bed2bba3ba75baafbbd0bd;
    inBuf[9617] = 256'h50c08cc313c79dcad7ce77d347d8e0dddee3efe994f084f770feaf05f80cf413;
    inBuf[9618] = 256'hd91a9221f1271c2e2234c639f13ea84393476a4a424cd44c094c6d4a1e485645;
    inBuf[9619] = 256'hd14278401f3e153ce3393f3778344131832d8a2922256a20a21bcc1672129b0e;
    inBuf[9620] = 256'h680b4e09e7070e07e90605073207f30702095c0a920c250fed11431585189d1b;
    inBuf[9621] = 256'hd91eab213d24e7263929812bf02df92fe931ce33353580369b3706380a386337;
    inBuf[9622] = 256'hba359133cc30592dd1290e26f621f11dbc193e15c510ff0bea06e201d4fceff7;
    inBuf[9623] = 256'h86f37fefe0ebbde8f7e596e39fe104e0bddeabddc3dc07dc6cdb13db1fdb9cdb;
    inBuf[9624] = 256'hbcdc90de04e11ce4ade76ceb2cefb6f2eaf5c1f838fb6dfd6aff2901b8020704;
    inBuf[9625] = 256'h15050b06e406b8079f084f09a809a809ff08b5070a06ec03880112ff63fc9bf9;
    inBuf[9626] = 256'hddf608f448f1b3ee33ecf5e9fee72fe6b9e49ae3b3e224e2dee1cae1fde164e2;
    inBuf[9627] = 256'hf2e2b3e389e480e5b7e62ae8ece90eec67eed4f048f3a8f5ecf722fa56fc6efe;
    inBuf[9628] = 256'h71005d021504a505df0686077707b10645057a03ae012000f4fe2dfe9ffd19fd;
    inBuf[9629] = 256'h75fc88fb37fa76f835f687f3a4f0baed09ebc9e80de7eee57fe5a6e549e640e7;
    inBuf[9630] = 256'h3ae8fce876e9afe9f4e99beac4eb76ed8eefb8f1ccf3bdf583f74ef93efb31fd;
    inBuf[9631] = 256'h26ff0a01ab0219047105a606dd072109310af80a510beb0ad9094a0844062804;
    inBuf[9632] = 256'h5402b6005aff39fef8fc8afbfaf913f8f1f5b6f331f17feee3eb5ee934e7abe5;
    inBuf[9633] = 256'h9be4f4e3a2e346e3cae238e271e1a2e008e09bdf84dfdddf72e03fe136e216e3;
    inBuf[9634] = 256'hede3c4e474e51ee6d3e677e737e826e91cea2ceb3aece8ec32ed0eed56ec5deb;
    inBuf[9635] = 256'h69ea7ae9dfe8aee89ae8aee8e0e8dce8c6e8b1e84ee8bbe705e7dee58de45de3;
    inBuf[9636] = 256'h43e2a4e1c9e15de268e3bde4b4e542e66de6f3e54ae5d4e47ce4a9e47ae588e6;
    inBuf[9637] = 256'hf8e7b1e930eb8eeca8ed0dee06eeb1edf1ec54ec0aece8eb42ecf7ec9aed47ee;
    inBuf[9638] = 256'hbaee93ee0bee1fedd0eb9deaa7e9efe8a9e89ce88ae86de804e840e73ce6dfe4;
    inBuf[9639] = 256'h59e3d1e13de0dcdeb8dda6dce5db68dbfedafada42db90db33dc05ddb9ddb8de;
    inBuf[9640] = 256'hebdf07e17ee239e4e6e5f7e766eadcecceef49f3fff664fb8f0018063c0cec12;
    inBuf[9641] = 256'h9c195f203027932d923343394c3ecd421c47274b2d4f8b532258dd5cb5613d66;
    inBuf[9642] = 256'h0c6aeb6c916ed56ecf6db06ba768eb64c9606d5cd8573f53b04ede49d5448e3f;
    inBuf[9643] = 256'h9c392d338d2c8225751edd176611510bf605cf0005fcfef740f401f1b5eedfec;
    inBuf[9644] = 256'ha2eb69ebbeebcdecfeeedcf165f5b2f917fe6e02be069b0a270e9811c314e317;
    inBuf[9645] = 256'h0e1b101e0c21e9237126cf28d82a5b2c782dd42d262d922bda2807259820961b;
    inBuf[9646] = 256'h1b1683109f0a4f04d9fd34f76af0e0e9a8e3acdd0cd8bcd288cd8ac8fcc3e3bf;
    inBuf[9647] = 256'h6bbce1b91cb8e2b64cb615b614b6c4b647b89bba3abefcc25bc86fcee7d43edb;
    inBuf[9648] = 256'haee131e887ee03f599fbd701fb07090ea8131819621e23236e27442b582ed430;
    inBuf[9649] = 256'hea328134bc35b1361c37e236f53521346931fb2df02984250e21c21cd7188115;
    inBuf[9650] = 256'hbf128310b40e1b0d970b120a7908e3066c052c0465033e03c2030b05f2063009;
    inBuf[9651] = 256'haa0b2f0ea3103b130116f2182d1c811fc322062623290e2cd32e2231cb32c333;
    inBuf[9652] = 256'hcc330933c431f52fdb2d9e2b032927261a23931fc21bbe174f13c60e4c0aa705;
    inBuf[9653] = 256'h12018cfcbff7ecf23bee94e960e5c7e191deeadbd7d921d800d784d682d611d7;
    inBuf[9654] = 256'h23d883d93edb4cdd92df16e2cee4afe7bdeaf7ed61f1f7f49ff859fc1100a803;
    inBuf[9655] = 256'h1e07540a150d570ff910db112412e8112f113510160fc30d590cdc0a25093807;
    inBuf[9656] = 256'h16059502beffaafc4af9c1f548f2e8eec8eb16e9b7e6abe404e39de177e0acdf;
    inBuf[9657] = 256'h16dfb4dea1dec2de2edf11e05ce11be34ee5bce751eafdec87eff5f148f462f6;
    inBuf[9658] = 256'h67f865fa3ffc0dfec2ff2b015d025403f40362048e04450493036902ba00ccfe;
    inBuf[9659] = 256'hc0fc9dfa8ef882f655f41cf2d7ef7eed3deb19e90be73ce5b0e35ee263e1bfe0;
    inBuf[9660] = 256'h5be04be094e024e108e236e380e4e1e54be7a5e813eab3eb7ced9fef28f2e9f4;
    inBuf[9661] = 256'hf2f72bfb34fe0001740341058b067207db07140849084b084b084f0802087f07;
    inBuf[9662] = 256'hc3067e05eb033802380038fe68fc84fab9f819f759f59cf3f3f112f014ee13ec;
    inBuf[9663] = 256'hdce9aae7bae5f7e38ee299e1dbe05ce027e00be022e088e014e1c0e182e21fe3;
    inBuf[9664] = 256'h84e3b7e3aae384e375e38ce3e6e392e46ee562e649e7f5e764e893e87ce84ae8;
    inBuf[9665] = 256'h08e8aae74ce7e7e665e6f0e588e51ae5d5e4b5e499e4b3e4f6e436e59ee517e6;
    inBuf[9666] = 256'h72e6eee683e706e8c4e8b5e9a5eae4eb75ed1bef15f14bf35cf57df7a8f990fb;
    inBuf[9667] = 256'h79fd5fffea0052028d034c04db04470542051505d5043f04ad034203b3023102;
    inBuf[9668] = 256'hb601dc00c3ff70fea0fc8afa49f8b4f511f37cf0d2ed42ebe8e8aae6bae43be3;
    inBuf[9669] = 256'h2be29de17fe1a0e1dfe11de256e28de2c1e20ae359e395e3e5e33ee497e43ce5;
    inBuf[9670] = 256'h18e606e74be8bce912eb97ec24ee77eff3f080f2d1f340f5a6f6a6f7a2f88bf9;
    inBuf[9671] = 256'h19facafaa4fb53fc46fd83fea6ff1501ed02e9047d07e10ac00e47136a18971d;
    inBuf[9672] = 256'hbb22c327432c54301a346a37753a793d68407443c8463f4ad84d8d512a558c58;
    inBuf[9673] = 256'h885be65d7a5f0b60935f245eaa5b4e584454794f354ad4444b3fde39d134c62f;
    inBuf[9674] = 256'hce2a1a263a214a1c93179a12750d89088503b3fe99fae3f6b3f35df168efeeed;
    inBuf[9675] = 256'h59ed5aed1beef3ef79f2b0f5c4f938fef5020608f00c9c111416051a7d1d8c20;
    inBuf[9676] = 256'hff220025a726e1270229232a1d2b0a2cbb2cce2c3e2cd62a5428e5248e20461b;
    inBuf[9677] = 256'h7215500ff008af02a8fcb5f6f8f07deb1be6fce054dc07d835d411d16ece5acc;
    inBuf[9678] = 256'h1ccb91caadcaafcb62cd8ecf65d2b6d549d967ddfae1d9e65bec6ef2c4f884ff;
    inBuf[9679] = 256'h7306210daf13fd19bf1f2b25362a8d2e5a329c351a380c3a873b5f3cbf3cae3c;
    inBuf[9680] = 256'hf43bab3ae03873369d338b30422df029962616237b1fa71ba417c6131c10b30c;
    inBuf[9681] = 256'hcb094607150577036102de0131022b03b604f4069d098c0ce40f5513bd16531a;
    inBuf[9682] = 256'hd41d2521782487273a2ade2c5c2fd03188344337d839443c1a3e363fad3f403f;
    inBuf[9683] = 256'hff3d0e3c31398d356531a22c902776223a1d1c184513760ed70981052d0110fd;
    inBuf[9684] = 256'h54f9c2f591f2e1ef56edfbeae2e8cbe6f3e4a7e3cae295e239e372e448e6e1e8;
    inBuf[9685] = 256'hf0eb64ef50f35bf74efb25ff930275050008330a1e0c040ed90f7a11ee121714;
    inBuf[9686] = 256'hda1452157e155115e914451450131a12b210130f550d950bd709150854068704;
    inBuf[9687] = 256'h920279004ffe24fc20fa7af846f7a3f6a7f633f731f89ef955fb3ffd4cff4101;
    inBuf[9688] = 256'h02039004d205ce06ae0782085b09510a540b590c5c0d3f0eef0e6a0f980f6b0f;
    inBuf[9689] = 256'hef0e270e0e0da50be709d1076705bc02e8ff0cfd3bfa80f7e9f47cf241f04aee;
    inBuf[9690] = 256'h95ec11ebbbe985e86de78ce6f3e5ace5c2e51de6afe67ee774e896e9fdea93ec;
    inBuf[9691] = 256'h5dee64f083f2c7f43af79af9defb08fecfff400179023f03ac03e303aa031b03;
    inBuf[9692] = 256'h8202b101d000190024fffcfdaafcc9fa88f814f62df31ef024ed02ea06e761e4;
    inBuf[9693] = 256'hc5e16cdf7cdda2db12dae6d8c0d7c5d60ed64ad5b2d478d465d4a7d454d515d6;
    inBuf[9694] = 256'he7d6c5d761d8d7d859d9d3d971da4adb17dccadc5add9cddafddb0dd8fdd67dd;
    inBuf[9695] = 256'h34ddcddc51dcbedbf5da1cda36d92ad833d755d672d5c2d439d4b1d373d37ed3;
    inBuf[9696] = 256'ha8d32ed4efd49dd577d674d767d8bbd978db53dd85dff8e151e4d6e680e9f8eb;
    inBuf[9697] = 256'h79eef5f016f31ff51bf7cff88efa63fc01fea1ff330152022503a90396033503;
    inBuf[9698] = 256'h9e0291015200edfe19fd25fb32f905f7eff406f3edf0ceeeb5ec4ceadfe7abe5;
    inBuf[9699] = 256'h70e374e1dddf37de9bdc33dbaed949d85bd7a5d64ad67ed6e0d673d779d8b3d9;
    inBuf[9700] = 256'h32db29dd53df80e1bae3b9e54be79ee8ace962ea02eb9eeb09ec57ec99ec9bec;
    inBuf[9701] = 256'h63ec28ecd5eb5eebfaea8eeae9e93fe98fe8b0e7eae64be681e5c3e428e45ae3;
    inBuf[9702] = 256'hb1e280e282e208e36ae44fe6e7e890eceaf004f620fca90269097a104b17ab1d;
    inBuf[9703] = 256'he923b629012f29340139793dee4151468c4ad24efc52ba56ec59525c945d935d;
    inBuf[9704] = 256'h565cd7593156b8518d4ca64646408d395032e42a8f231e1ccd14cc0db606b5ff;
    inBuf[9705] = 256'h1cf9a9f2adec99e71ce353df83dc33da6ed891d744d79ad7f8d80fdbdadda9e1;
    inBuf[9706] = 256'h32e661eb6cf1fef7e0fe0b061b0dcc130e1a9e1f62246d28b82b572e6830ec31;
    inBuf[9707] = 256'hf13275336b33d932ab31d52f562dfb29ae259420ab1a1314240de50557fecef6;
    inBuf[9708] = 256'h44efd2e7e9e09fdafed42bd020cca6c8c5c597c307c22dc14ac14bc219c4e4c6;
    inBuf[9709] = 256'h7fcaabce93d317d9e9de3ae5eeeba5f28ff98f003d07d80d67148e1a88204426;
    inBuf[9710] = 256'h342b6a2fce32e934003646368535183426326e2f3d2cc428e424f320151d1619;
    inBuf[9711] = 256'h171501118f0cea0722033efe9df966f5a8f1aeee82ec1febafea1beb51ec67ee;
    inBuf[9712] = 256'h3ff1cbf40df9cffdee025208cc0d5313f018891e1a248129892e27334737d33a;
    inBuf[9713] = 256'he03d5240fb41e142ec4213428f406a3e9b3b4c386234bc2f862ac124581e9017;
    inBuf[9714] = 256'h81101d09c1019ffaabf32bed35e78ee15ddcc0d78fd302d03ccdfcca6ac9bdc8;
    inBuf[9715] = 256'hc5c8aec9a8cb63ced2d1efd54edadadea7e371e835ed13f2cff659fbcdff1104;
    inBuf[9716] = 256'h1008f00b980feb12e1155218151a1f1b731b101b081a9318cb16b9148c123a10;
    inBuf[9717] = 256'h9c0dce0acd079204680172fe9dfb1ef9f6f6fef465f33af261f102f11ff17df1;
    inBuf[9718] = 256'h1ff205f318f478f539f74df9bafb74fe5a0153044607190ab00cf20ed2104312;
    inBuf[9719] = 256'h4713eb132114d9131913dd113310440e240cdd097c07f9045b02adfffdfc65fa;
    inBuf[9720] = 256'he5f771f514f3bbf065ee31ec1dea35e89ce64ce55fe404e434e4f3e44de608e8;
    inBuf[9721] = 256'h06ea4beca3ee0cf19cf32bf6b2f840fbaefd090067029e04af069108040a0e0b;
    inBuf[9722] = 256'hb30bc20b530b710af9081f070405a4024300edfd77fb05f999f606f483f125ef;
    inBuf[9723] = 256'hc7ec8bea73e860e682e4efe28ae17ce0cadf4bdf19df45dfb1df6fe07fe1b7e2;
    inBuf[9724] = 256'h20e4bbe564e71ce9e6ea9dec3feecfef37f18ef2e1f321f55af686f77df832f9;
    inBuf[9725] = 256'h93f979f9f2f806f8b0f620f56ef390f1b5efebed24ec92ea37e9f6e7f3e626e6;
    inBuf[9726] = 256'h6ee5f3e4b3e48ce4aee416e5aae598e6d1e725e9aaea43eccfed7fef50f129f3;
    inBuf[9727] = 256'h36f567f7a0f904fc84fe08019d031a064b08350ab90bbd0c5b0d8c0d470db20c;
    inBuf[9728] = 256'he20be90af3090e09240837073406fa04970315026500a6fef6fc4ffbd1f99bf8;
    inBuf[9729] = 256'h90f7b6f60ef671f5eff49bf458f43cf455f479f4b9f428f5a6f556f644f743f8;
    inBuf[9730] = 256'h58f96bfa39fbc4fb02fcdbfb7dfb06fb79fa07fabcf98cf98af9a3f9baf9c0f9;
    inBuf[9731] = 256'h8bf902f916f8bef61cf545f34bf16fefb7ed1cecd5eab9e99fe8bbe7dce6e1e5;
    inBuf[9732] = 256'h2de59de40be4dfe3f1e311e4bbe4d1e50de7dae800eb18ed7fef15f275f4f9f6;
    inBuf[9733] = 256'h88f9b3fbd6fd0e002402a104d5078c0b16109115871bf221be28602fb735b93b;
    inBuf[9734] = 256'h024189456849774cd44ec6505e52cf534755b5560b582259bf59c9590c597957;
    inBuf[9735] = 256'h2e551752514e264a7f4581408a3b6e364c317a2c9d27a822dc1dcd188a13950e;
    inBuf[9736] = 256'hb1091605560119fe6dfbc1f9a6f826f8a3f8a2f91ffb67fdf9ffd5024706e009;
    inBuf[9737] = 256'hb10d08127b16131bf01f8824c528b52ce92f7b329634f435bb361237bd36f435;
    inBuf[9738] = 256'he8346d33af31b52f2c2d1d2a81262122331de7173712680cac06ea0052fb13f6;
    inBuf[9739] = 256'h1ff1aeecf6e8d9e562e3aae177e0c3dfb7df26e009e18ce27ee4cde6afe9f6ec;
    inBuf[9740] = 256'h8af09ff404f996fd83029207860c6c11fd15fc19911daa203323692535277728;
    inBuf[9741] = 256'h5629be299b29142912287c267024e221d61e831bf51737147b10c50c2509d105;
    inBuf[9742] = 256'hc8020500a1fd79fb77f9bef747f620f58bf48bf421f57af67ff80ffb44fef301;
    inBuf[9743] = 256'hed05470adb0e7c134718181dbe214d269c2a792efa31fc3455371939263a653a;
    inBuf[9744] = 256'h033a0a399737ee3510340032c72f362d462a052754234a1ffa1a3b162911e50b;
    inBuf[9745] = 256'h5a06d10089fb75f6d6f1d8ed4aea5ce72be57fe37fe248e294e276e3fbe4c9e6;
    inBuf[9746] = 256'he1e851ebceed62f02ef3f0f5a5f865fbf9fd6100d10233058f07060a6c0c9c0e;
    inBuf[9747] = 256'h9510351267133f14be14d7148b14dc13be123911750f8d0d910bad09f5075306;
    inBuf[9748] = 256'he304af039002a001f1005800edffccffc2ffddff36009100f4007b01ef015202;
    inBuf[9749] = 256'hc10207032703470344032c032a0323031d03320336031f03ee027302a0017e00;
    inBuf[9750] = 256'heefe00fdcdfa4bf898f5d2f2f4ef1bed66eacae765e553e380e1ffdfdbdeebdd;
    inBuf[9751] = 256'h36ddcddc8fdc92dcf1dc7cdd35de23df08e0f1e001e211e33fe4abe517e78de8;
    inBuf[9752] = 256'h1bea76ebaeecddedc1ee7def38f0acf001f154f14ff11df1daf032f05aef69ee;
    inBuf[9753] = 256'h01ed5deb9ce979e752e55de355e18ddf18de99dc56db62da66d9b1d84ad8d2d7;
    inBuf[9754] = 256'h8fd788d76cd791d705d876d82dd927da0cdb1fdc64dd88decedf31e154e26ce3;
    inBuf[9755] = 256'h72e414e595e506e629e642e65fe633e6eee598e5e7e416e43ae318e2e8e0b9df;
    inBuf[9756] = 256'h4bded2dc65dbcdd94dd8fcd69fd570d472d361d279d1c4d011d0b6cfc3cf02d0;
    inBuf[9757] = 256'hbed0ead138d3ebd4ead6e6d825db85ddaedfe9e119e4fae5ece7e0e996eb66ed;
    inBuf[9758] = 256'h36efbef04df2c7f3dff4dcf5a0f6e3f6f5f6caf62ff67bf5b1f49ff398f29df1;
    inBuf[9759] = 256'h73f060ef5eee2fed17ec25eb1bea3ee994e8cce71be78de6dae54be502e5b3e4;
    inBuf[9760] = 256'h9ee4d5e4f5e438e5c2e53ee6f1e6f8e7e8e8ece90aebd5eb81ec25ed68ed8aed;
    inBuf[9761] = 256'ha1ed50edd5ec3aec2aebeee995e8e0e62ae585e3bbe120e0b7de44dd15dc25db;
    inBuf[9762] = 256'h3dda9cd929d9a9d846d8e9d76dd70bd7b9d672d667d692d6f4d6aad799d8c1d9;
    inBuf[9763] = 256'h20db8cdc14deb1df39e1c9e251e496e5c3e6d1e791e854e92deaebead9ebfbec;
    inBuf[9764] = 256'hf9ed0def46f050f172f2dbf334f5b2f680f83dfa11fc46fe95002d036606f609;
    inBuf[9765] = 256'he50d73124217351c7d21c426e62b0d31ef35623a823e1c421d45af47c5495d4b;
    inBuf[9766] = 256'h8c4c3c4d654d034d124ca84abd485746954358409f3c95380d340b2fd0293124;
    inBuf[9767] = 256'h421e5c185712500ca606310112fca9f7c8f385f031ee8beca4ebc1eb9aec31ee;
    inBuf[9768] = 256'haaf09ef3fbf6d9fae2fe1a03a5072f0cb9105215a419b51d9b2117253428072b;
    inBuf[9769] = 256'h532d1d2f7130123108316330002ff92c6a2a3d278823671fd31aef15ec10ce0b;
    inBuf[9770] = 256'hb106ac01b2fcd4f737f3ddeee4ea6ce763e4c6e1acdf00decddc43dc59dc1edd;
    inBuf[9771] = 256'hb6defce0dde36be763eba1ef36f4e5f884fd3002af06db0ade0e9c1204164e19;
    inBuf[9772] = 256'h551ce51e1321a7227323b0235a236d222a21901f831d391bae18d815f2120210;
    inBuf[9773] = 256'hfb0c060a1a071f043b016cfeb3fb51f958f7cdf5e4f48bf4a2f448f56af6faf7;
    inBuf[9774] = 256'h2bfae5fcffff89034b07180b180f36135c17bb1b28206a249f28982c27307533;
    inBuf[9775] = 256'h6136bd38a03ae53b5d3c2e3c4b3bb539b0375035a932f82f372d612a9527b524;
    inBuf[9776] = 256'hb921ba1e911b3918cf1430117d0df80992067d030001eefe62fd95fc46fc81fc;
    inBuf[9777] = 256'h7dfddcfe9200cb0213055a07e409550cab0e3911a513d91524182a1ad51b721d;
    inBuf[9778] = 256'hb21e791f0e202d20c91f3f1f721e691d7b1c8d1b921ab219b9188c173d16b114;
    inBuf[9779] = 256'hfe125711c70f750e790dbc0c4e0c230c1c0c4b0c9a0cdd0c240d5c0d6d0d8c0d;
    inBuf[9780] = 256'hcc0d2c0ee10edf0ff51028124c131b149514ac14371457131c127210820e6f0c;
    inBuf[9781] = 256'h340af307ce05a70378013fffcffc2dfa75f79ff4cdf12cefb4ec86eacae86ee7;
    inBuf[9782] = 256'h87e62de63ae6b5e6a2e7cbe82ceac7eb67ed13efd5f08bf242f4fef5a2f73cf9;
    inBuf[9783] = 256'hdafa76fc27fee9ffa10140039a04a0055406a506aa067806fb0556059804a903;
    inBuf[9784] = 256'hb902d201c400baffadfe5cfdfafb94faf2f85ff705f6b7f4c0f33df3e9f2f1f2;
    inBuf[9785] = 256'h5df3ddf38cf46df537f6faf6bdf74df8c6f844f9aaf90afa76facafa01fb1ffb;
    inBuf[9786] = 256'h08fbb8fa3dfa90f9aff8b0f797f665f52ff4f7f2acf14df0d5ee31ed63eb73e9;
    inBuf[9787] = 256'h63e743e525e324e15edfebddf2dc87dca2dc51dd83de07e0d2e1c3e39be560e7;
    inBuf[9788] = 256'h04e969eac6eb3aedc8eeb9f015f3adf59af8b0fba3fe820125044e0625089609;
    inBuf[9789] = 256'h7f0a1c0b680b440bec0a570a67094b08f7064b0573036e012fffeffcbafa8ff8;
    inBuf[9790] = 256'ha2f6f0f465f319f2fcf0edef04ef46ee98ed17edd5ecb2ecbbec08ed81ed3aee;
    inBuf[9791] = 256'h55efb6f05ef250f446f620f8e1f956fb8dfcacfd93fe56ff0a007700a0009600;
    inBuf[9792] = 256'h27006cff81fe4cfdf2fb76fa9bf887f649f4caf163ef3aed2ceb6de9f8e794e6;
    inBuf[9793] = 256'h76e5a6e4fbe39ae378e363e370e39ce3d8e351e419e52be699e759e94feb57ed;
    inBuf[9794] = 256'h4def1ef199f2abf372f4d7f4d7f4bbf470f4e7f370f3f6f257f2e8f18df105f1;
    inBuf[9795] = 256'h93f01ef060efa6eef8ed24ed87ec4eec4cecd0ec01ee9befb5f166f460f7b5fa;
    inBuf[9796] = 256'h9afee902b7073a0d38138d194f203c27202e0135953b8641c446204b7b4ef450;
    inBuf[9797] = 256'h9f528353b753475337527650004ed44acd46ea41643c4136ac2ff82819221e1b;
    inBuf[9798] = 256'h4e14980d1f073e01d4fbddf680f268ee8bea35e748e4f7e1abe039e0c1e08be2;
    inBuf[9799] = 256'h46e5f6e8c7ed4bf36cf931000f07d90d9214be1a54208325022ae42d4a31da33;
    inBuf[9800] = 256'h9035893683369d351534c631cc2e562b4827bc22ec1de418d213e20e140a6705;
    inBuf[9801] = 256'hcb0026fc75f7c1f229eee1e909e6bfe229e051de4add3ddd3bde3ae032e3ffe6;
    inBuf[9802] = 256'h61eb33f053f58bfac5fff904f6099b0ee712a816c2194a1c2a1e611f2c209520;
    inBuf[9803] = 256'h9f207a200120061f9b1d991bea18cb154c12740e830a7c0653023afe3ffa6af6;
    inBuf[9804] = 256'hf8f2f8ef68ed5debc0e986e8d8e7b4e72ae86fe96deb0fee59f109f5e1f8e2fc;
    inBuf[9805] = 256'hd900a8047c084e0c0810ce138b17151b7f1eba219c2435277429252b542c012d;
    inBuf[9806] = 256'h052d6f2c5d2bc429bf2788253823db208a1e331cb5191d178a140b12c20fd10d;
    inBuf[9807] = 256'h100c550a9908b506ad04d5024b01170073ff4bff51ff85ffc5ffc2ff94ff4bff;
    inBuf[9808] = 256'hb9fe13fe7ffdc6fc09fc7afbecfa7cfa5afa45fa1dfae6f954f94bf8f5f64cf5;
    inBuf[9809] = 256'h65f383f1b7ef0bee9fec6beb70eac3e971e985e912ea17eb75ecfded9fef4df1;
    inBuf[9810] = 256'hf6f2c5f4d6f60df971fbf2fd430063026a043906ef07aa09300b7d0c880d0e0e;
    inBuf[9811] = 256'h200ee20d410d720c940b750a150967072f05870291ff40fcc1f82bf567f1aeed;
    inBuf[9812] = 256'h3bea31e7eae488e3d6e2b4e2d7e2cce281e20ae269e1e8e0d6e046e156e206e4;
    inBuf[9813] = 256'h21e681e8ffea62eda0efb9f186f30df56af697f7b4f8eef93ffba1fc00fe0eff;
    inBuf[9814] = 256'ha2ff9bffc4fe3efd2ffb90f8aff5c3f2c0efeeec75ea2de85fe627e545e4ebe3;
    inBuf[9815] = 256'h11e439e46de495e437e49ee30de366e22ee2c3e2e3e3c1e54ae8d7ea59edbdef;
    inBuf[9816] = 256'h90f102f339f4f0f460f5a9f58df54cf508f588f4f5f355f355f200f142efc5ec;
    inBuf[9817] = 256'habe914e60ce20fde6eda27d773d44ad260d0d7ceb5cdc7cc3fcc25cc2bcc6ccc;
    inBuf[9818] = 256'he2cc55cd0dce35cfa8d0a1d21ed5b9d77bda4cdde1df79e233e5e2e7bbeaa5ed;
    inBuf[9819] = 256'h2bf05bf21bf42bf5ebf57af6b9f6fbf622f7dbf666f6a9f55ef4d4f2f5f080ee;
    inBuf[9820] = 256'he0eb36e985e65fe4e8e2eee19ae199e16ce120e1a2e0dddf45df0bdf24dfc8df;
    inBuf[9821] = 256'he5e03fe2ede3dbe5c8e7b5e975ebc1ecbeed9aee78efbef0a2f2fef4abf751fa;
    inBuf[9822] = 256'h71fce6fd98fe72fec4fdc6fc71fb13fad0f882f765f690f5caf43ef4f4f38ff3;
    inBuf[9823] = 256'h1cf38bf287f142f0e8ee66ed1dec3aeb91ea4bea55ea5cea8aeadfea2cebb2eb;
    inBuf[9824] = 256'h6dec18edcded78eeecee56efcfef60f037f147f276f3bef4f1f5f7f6d5f77df8;
    inBuf[9825] = 256'hf8f841f940f906f994f8e9f742f7a3f6f4f54af56af41cf396f1d1efd7ed19ec;
    inBuf[9826] = 256'ha2ea61e9b3e88fe8cfe8b9e92debc2ec75ee0cf036f138f247f368f4fef545f8;
    inBuf[9827] = 256'h0ffb67fe49025806880aee0e6113f717ec1c2522a7278a2d91337e392b3f2544;
    inBuf[9828] = 256'h0848a44ad04ba24b754a9f487a464c4428420b40d33d5a3b8d382b351031492c;
    inBuf[9829] = 256'hb9268e20441a0b14350e3b0901056d0183fec8fb0cf97df6e7f37ef1bfef90ee;
    inBuf[9830] = 256'h26eeddee58f08ff2bcf562f95bfdd0014306980a110f5a137217971b691fc822;
    inBuf[9831] = 256'hc9250b287e295e2a832a0c2a46291d289426c9248a22ce1fb71c4b19b0152512;
    inBuf[9832] = 256'hce0ec90b2809df06d404df02d900b6fe73fc32fa3ff8c9f6e1f5a2f503f6d3f6;
    inBuf[9833] = 256'h12f8c4f9bdfbeefd4b008502850469061b08b709960ba00db40fd911af13e914;
    inBuf[9834] = 256'ha415b8152c155e143e13b511fd0fe40d540bbe084106ff036a026a01b6004400;
    inBuf[9835] = 256'hb8ffdefe11fe8bfd99fda9fe9100f10280059c07f608cc093e0aab0aa60b210d;
    inBuf[9836] = 256'hec0e12114d1394154018371b3c1e3a21ae232825d325dd259f25b3252c26c026;
    inBuf[9837] = 256'h2c27e1267c254423af20571ef81cce1c971dd81ed61f11208f1f861e6e1dc21c;
    inBuf[9838] = 256'h841c981cdd1c031d191d631dd51d7c1e461fb01f881fdd1e8f1df21b711ae518;
    inBuf[9839] = 256'h60170a167b14b8121d11830f040ee60cc70b740af708f2067b041102cafff0fd;
    inBuf[9840] = 256'hecfc7afc71fccefc1bfd2bfd1efdbbfc1afc9afb4ffb8cfbcafc11ff5c028306;
    inBuf[9841] = 256'he10ada0e0012ee13c31403153015d015291709190c1baf1c891d8a1ddd1cd51b;
    inBuf[9842] = 256'hce1ae319fb18eb176e166b140f12880f140ddb0ab5088b0667044902680017ff;
    inBuf[9843] = 256'h47febdfd36fd3afc7bfa28f8a5f573f31af2bbf10af2acf23af372f399f328f4;
    inBuf[9844] = 256'h67f57df729fab2fc84fe68ff44ff59fe23fde5fbb7fa9cf97af851f752f6aff5;
    inBuf[9845] = 256'h8ef5f3f5a3f643f782f738f76cf65ff584f425f44df4f2f4d0f587f60af76df7;
    inBuf[9846] = 256'hbff75df87ef9e5fa66fcbafd76fea6fe8ffe64fea3fe97ff1f012d036d054007;
    inBuf[9847] = 256'h6608b208ee0769069804c20250016600caff59ffc7feaefd09fcd3f9fdf6c6f3;
    inBuf[9848] = 256'h6ff020ed43ea2fe8fee6c0e653e749e845e9efe9ffe976e995e8a6e703e7f2e6;
    inBuf[9849] = 256'h86e7a1e80cea86ebe4ec1dee3bef5ef099f1e5f229f443f51cf6c4f65df71df8;
    inBuf[9850] = 256'h3af99efa06fc2afd95fdf5fc78fb5cf901f707f5b4f30bf324f3c6f39ef4aef5;
    inBuf[9851] = 256'hc9f6b7f785f804f904f9c4f86af825f876f898f97bfb0bfed70049030c051106;
    inBuf[9852] = 256'h4d062806fa05b8059b057c053405e104870435040604db03950319033c020401;
    inBuf[9853] = 256'h83ffb1fda2fb6df91ef7e1f4fef2b8f13af18ef1a0f215f48cf5d5f6aff712f8;
    inBuf[9854] = 256'h3df83df826f82af824f810f832f87ef810f92bfa8cfbfcfc6afe68ffd2ffc3ff;
    inBuf[9855] = 256'h0affc5fd30fc35fa0ef8f2f5c6f3bff1fbef4beedcecc5ebdbea3feaf6e9d8e9;
    inBuf[9856] = 256'hfee95eead3ea5febdeeb22ec33ec0aecabeb46eb10eb30ebaeeb8decb3edc9ee;
    inBuf[9857] = 256'hadef67f0c9f0faf057f1c6f142f2eaf24df31df37bf235f13cef08edc6ea87e8;
    inBuf[9858] = 256'hd8e604e6f4e5e6e6dde842ebe3edc5f084f34af6aef9a4fd3e02d107e70d1d14;
    inBuf[9859] = 256'h8f1ad220a926642cda31fb36173c02419745d649654dff4f7b519a5179504c4e;
    inBuf[9860] = 256'h2e4b8b478043f93e173a9334592ecd27ff203f1a1114490ee308f20305ff36fa;
    inBuf[9861] = 256'hd4f5baf145eebaebcae9b9e8a6e850e919eb07ee9af1e8f5adfa56ff2b043609;
    inBuf[9862] = 256'h390e9e135419ce1e0f24d828ac2caf2ff0313633a3333233a6311f2fcf2bca27;
    inBuf[9863] = 256'h5023981ea21974141e0fa309310404ff39faf7f53ff2e1eee0eb3ee900e778e5;
    inBuf[9864] = 256'hc7e4d9e4c5e528e76ee89ee9a1ea6bebaaecb8ee88f15ef5eef986fef002c506;
    inBuf[9865] = 256'h9409860bb30c2e0d6b0dad0dff0d6c0ea90e550e230dcc0a5407ee02e7fdc0f8;
    inBuf[9866] = 256'hdaf379efe5eb13e9dce623e5a3e33ee204e10fe098dfc5dfaee055e263e4b1e6;
    inBuf[9867] = 256'h55e900ecb1eec2f1e5f400f861fba9feb801e504d5075a0aa30c5f0e800f4010;
    inBuf[9868] = 256'hd710721149127213851439153a155114ae12d6104e0f5e0e2c0e760ea80e940e;
    inBuf[9869] = 256'h3b0ea30d5c0ddc0dfb0ea810b1127614d6150517f217c618bb19851adf1ad01a;
    inBuf[9870] = 256'h571a8a19c9184518b917da1666150113c10f340ca6085d059802eeffe4fc5ff9;
    inBuf[9871] = 256'h31f58cf023ec5ce880e5d8e323e300e33ae37ce3ade307e4bae404e619e8edea;
    inBuf[9872] = 256'h57ee1ff208f6ebf9b4fd690105056d08a70ba80e5611d9132f162b18e519451b;
    inBuf[9873] = 256'h121c8b1ccd1cb81c8f1c391c3e1ba0194217de13db0f9f0b3f073803c4ff8cfc;
    inBuf[9874] = 256'h82f991f658f3f9efd1ecf4e9aae73ee684e55be5dae5cde616e8c4e988ebf7ec;
    inBuf[9875] = 256'heded41eefaed9feda1ed2fee61efe8f02ef2d7f2c8f21bf23cf19ef071f09ef0;
    inBuf[9876] = 256'hf9f01af189f021ef07ed6feaa1e709e5e4e249e17be07ae000e1fee12ae30ee4;
    inBuf[9877] = 256'hb0e429e577e514e651e7ffe823eb7fed79ef02f12ef2fdf2eff35df51ff733f9;
    inBuf[9878] = 256'h47fbc4fca0fde2fd86fdf7fc54fc61fb28fa7ff82df692f3f4f06aee5eecdbea;
    inBuf[9879] = 256'h9de9bde823e884e7fee687e6e0e529e576e4ade303e3a1e26fe28de211e3d4e3;
    inBuf[9880] = 256'hc2e4c6e597e614e747e753e795e769e8e1e9dcebe9ed70ef1bf0c2ef87eef8ec;
    inBuf[9881] = 256'h81eb5eead7e9c0e9b8e9bce9a0e939e9eae8d4e8d6e838e9e6e979ea1aebc1eb;
    inBuf[9882] = 256'h1cec6cecb8ecb3eca6ecc5ec0eedfeedd6ef56f261f58cf82bfb0cfd24fe7efe;
    inBuf[9883] = 256'h8afe8ffe8efe8ffe54fe94fd48fc5efae0f712f512f20bef5bec2deaa1e8dde7;
    inBuf[9884] = 256'haae7abe7b0e77fe709e79ee681e6c9e68ce79ae88ae931ea87ea86ea7feac8ea;
    inBuf[9885] = 256'h77ebb4ec94eee6f09bf3adf6ddf91cfd5f005d03fd0517084c098709c208f106;
    inBuf[9886] = 256'h8304e70157ff40fda8fb29faa1f8bff627f421f1e8ed97eaafe74ee53be39fe1;
    inBuf[9887] = 256'h63e058dfd1dee5de69df74e0c6e1fae21ce438e567e604e81bea76ecd2eecdf0;
    inBuf[9888] = 256'h36f229f3def3b0f4c2f5eaf60af8dff841f984f9d8f944faf2fa87fb80fbe9fa;
    inBuf[9889] = 256'hbaf90ef891f67cf59ef40df46cf342f2daf078ef4eee11eefceebbf035f3fff5;
    inBuf[9890] = 256'h79f8bcfa06fd7fffc9023c079a0cbe124919971f92254b2bbd303236be3b0541;
    inBuf[9891] = 256'hcd45bf497b4c234ef24e114fd94e494e134d1d4b33484844d73f363bac36a032;
    inBuf[9892] = 256'he32e1e2b4527ff22381e5d198014d40fca0b2e08f6046f02660001ffc0fe63ff;
    inBuf[9893] = 256'hda0047030506e3082c0c850f04130217e41a651ea7212424f825bd274229a22a;
    inBuf[9894] = 256'h312c742d4c2e002f342fd62e162e922c3a2a6a272c24ce20bc1dd61af717fe14;
    inBuf[9895] = 256'h8d11a80d9809a1054f020700c9fe91fe12ffcbffa0009301a2022d045b06db08;
    inBuf[9896] = 256'h600b920dfe0ebc0f2d1075100011111239133014e7140b15d314d41412158915;
    inBuf[9897] = 256'h2b1638162315f3129e0f910bb7076e04e801530038ff2ffe35fd19fcfafa48fa;
    inBuf[9898] = 256'h11fa6afa74fbd8fc65fe1c00c9018803ad052808fe0a2d0e3e11f1134e163418;
    inBuf[9899] = 256'hd419891b421de51e6b207a21de21b321eb20831fab1d661bb418d9150c137810;
    inBuf[9900] = 256'h6a0eff0c1e0cb20b850b520b060ba70a5c0a6d0a0c0b4d0c1c0e29103e124114;
    inBuf[9901] = 256'h1616e417d919c31b8e1d291f4020f22090210e2291222f236a230b231d225e20;
    inBuf[9902] = 256'hf81d4b1b3318bd141611010d97082b04b3ff60fb7bf7e4f3c0f048ee60ec26eb;
    inBuf[9903] = 256'haaeaa3ea0bebe7eb08ed98eeaef012f3c0f5a8f88cfb95fef601a505b509030e;
    inBuf[9904] = 256'h02126015f5179c198f1a321bbb1b441cc21cf11c8d1c851bfb1927185016bb14;
    inBuf[9905] = 256'h63131312b110140f140de50aac0856060404c80177ff42fd72fbf6f9e0f845f8;
    inBuf[9906] = 256'hccf756f725f742f7e0f75ef98cfbfbfd66004c024c0393035203a602de010301;
    inBuf[9907] = 256'hd3ff3bfe38fcc8f931f7d4f4dff26ff17ff0d4ef1fef35eeffec7debd7e947e8;
    inBuf[9908] = 256'hdee69de593e4b1e303e3dfe297e358e543e805ece6ef50f3cbf52bf7f3f7d4f8;
    inBuf[9909] = 256'h4cfab3fcd3ffee027105ec063507c2061d0694057b05b405cb059105cc044103;
    inBuf[9910] = 256'h2f01bdfedafbd5f8d4f5d0f233f047eef4ec61ec66ec70ec58ec0bec5aeb9dea;
    inBuf[9911] = 256'h2beaf8e922eaafea50eb07ecececd0edb4ee94ef29f05cf046f0e4ef5befdcee;
    inBuf[9912] = 256'h61eee4ed5fedafeccdebc6ea9de975e869e779e6b2e508e55be4c0e34be3fbe2;
    inBuf[9913] = 256'h06e36ae3dee349e482e455e40ee404e459e45de50de7f0e8ccea57ec42edd7ed;
    inBuf[9914] = 256'h6aee21ef5af010f2d3f381f5d8f69cf72cf8c0f852f918fac9fae3fa69fa48f9;
    inBuf[9915] = 256'h8cf7d7f57ef48af338f33df31bf3c7f20ff2d6f08fef6fee87ed2aed48eda0ed;
    inBuf[9916] = 256'h43ee13efe1efd0f0d8f1c3f295f338f483f496f496f498f4cef44cf5e9f585f6;
    inBuf[9917] = 256'hedf6e6f679f6d1f50ff576f420f4daf38df318f34cf25af17bf0a7ef06ef92ee;
    inBuf[9918] = 256'hfced59edc9ec49ec3becd2eccfed32efb2f0c2f160f281f2f9f13df18df0d4ef;
    inBuf[9919] = 256'h77ef82efa4ef0cf0abf02af1bdf165f2daf243f391f36af3e0f2fbf1b3f063ef;
    inBuf[9920] = 256'h58eea2ed4ced1eedbbeceaeb94eae0e814e76ce523e428e344e26ae173e042df;
    inBuf[9921] = 256'h1ade0edd05dc26db56da4fd946d86dd7ced6e4d6f5d7c1d93cdc4cdf7ae2c8e5;
    inBuf[9922] = 256'h71e94fed65f1d3f544fa99fe1d03cf07ca0c54122518e11d6f237b28e12ce430;
    inBuf[9923] = 256'h8234b037983a073dd03e02406140bf3f233e663b913707330f2e02294024cc1f;
    inBuf[9924] = 256'h8b1b5417e212290e38092b044effd0fae0f6d3f3c4f1d4f035f197f29df40af7;
    inBuf[9925] = 256'h4df939fb1ffd0aff4d015704d407840b520fa012421588174419a01a121c6c1d;
    inBuf[9926] = 256'haa1e0a203621fd2179226322ac219b20401fcc1d831c601b4b1a1e199c17b415;
    inBuf[9927] = 256'h6213c710390ee90bfa09a708dd0775076c0783077a075107f3066b0621065f06;
    inBuf[9928] = 256'h49070c096b0bce0dc10fdb10d410e90f8a0ef90c7d0b260a92087d06e903d600;
    inBuf[9929] = 256'h9afdcdfaa9f837f769f6c6f5d5f476f392f164ef7eed43ecffebd0ec52ee0ef0;
    inBuf[9930] = 256'hacf1d0f28ef34bf42cf55bf6ddf742f94cfa22fbdcfbdafc9dfe0501a003fe05;
    inBuf[9931] = 256'h7807b80721074606b80507062d07800855091c097b07d6040602bdff84fe93fe;
    inBuf[9932] = 256'h74ff9300a4017602380380049e0695093e0d08114414a61632182e192b1aac1b;
    inBuf[9933] = 256'hd01d5220b6226b24fb24662405232221111f0f1de11a58188f158312680fa60c;
    inBuf[9934] = 256'h2b0abc072905fc010efebaf95af584f1ceee37ed99ecb4ecf7ec35ed97ed13ee;
    inBuf[9935] = 256'hddee2cf0b8f175f381f5bcf752fa85fd1c01db049f080f0c090fbc114214a716;
    inBuf[9936] = 256'hff181b1ba51c701d6b1d801cd01aae184316bd138311bb0f640ebb0da50dba0d;
    inBuf[9937] = 256'he10dd60d2f0d170ccd0a5a0921086e070f07fb063c078607c7072c089608e608;
    inBuf[9938] = 256'h31094c09f4082e0804076b05a9030f02a20073ff7bfe5dfde6fb1ffa03f8c7f5;
    inBuf[9939] = 256'hc1f3e9f121f049ee19ec90e90be7ebe4aee3ade3c2e477e633e85be9b2e96be9;
    inBuf[9940] = 256'h0ee946e983eadaec0af088f3e4f6ecf993fc13ff990106043d0609082209a309;
    inBuf[9941] = 256'hc2099c09820985096a093409c508db07aa063f0575039801c2ffccfd00fc75fa;
    inBuf[9942] = 256'he6f86ef70af669f4aef2f8f029ef7ded2eec2deba9eac5ea54eb3bec4aed21ee;
    inBuf[9943] = 256'h91ee93ee39eecbed9cedcded5bee15efa9efd6ef8aefdeee0dee4beda6ec0cec;
    inBuf[9944] = 256'h44eb19ea8ee8d0e62be50ce4aae3fae3e6e420e641e73ce80be995e91ceac8ea;
    inBuf[9945] = 256'h7eeb6eecb0ed10efacf08af25df428f6d8f722f91dfadafa44fba4fb1dfc8efc;
    inBuf[9946] = 256'h19fda3fde3fdfcfdeefdadfd95fdaefdb8fdb4fd47fd01fc05fa7cf7a0f417f2;
    inBuf[9947] = 256'h2bf0c6eeeced4feda2ec19ecf1eb57ec88ed5cef54f111f34cf4f1f458f5ddf5;
    inBuf[9948] = 256'haaf6c4f7f5f8def949fa37facff94cf9e1f894f84ef8e7f749f788f6c7f526f5;
    inBuf[9949] = 256'hc6f491f450f4f3f36ff3c1f225f2b2f132f192f09eef17ee41ec88ea39e9e0e8;
    inBuf[9950] = 256'hc1e98feb09eeacf0c2f20df476f406f442f385f2e0f184f149f1e4f082f041f0;
    inBuf[9951] = 256'h33f0a6f06ff116f261f2fff1def085ef6beef3ed65ee81efccf0e2f15af23ef2;
    inBuf[9952] = 256'heef1c1f114f2f0f2e4f38cf47ef47ff3fef175f033efa5eea7eebdeedaeeceee;
    inBuf[9953] = 256'h77ee41ee3fee3bee71eed8ee49ef45f0fcf13bf42af78bfacafdec00f203b506;
    inBuf[9954] = 256'h8f09ad0cd70f191353162a19b81b191e41207822db243827a4291f2c8d2e2831;
    inBuf[9955] = 256'hf833bb365239623b7a3ca23cef3b843ad838133720351233a830ac2d642aef26;
    inBuf[9956] = 256'h9923fe202a1ff41d421d581cb91a9b180d16951332120512f612f91432171419;
    inBuf[9957] = 256'hcd1a221c401db01e0820fd20a4217a219d20e01f681f871fa6201b2258234524;
    inBuf[9958] = 256'h6324d5234923cb228922b122b6225622b1219520421f1b1ef51cd51bb61a2f19;
    inBuf[9959] = 256'h4d174315ff12dc102a0fcb0de60c8f0c7b0cb50c470dde0d7b0e240f8b0fcc0f;
    inBuf[9960] = 256'h20106b10dc109411351292129912e2116c108d0e4b0cf7092208d3061106fb05;
    inBuf[9961] = 256'h1006dc0550051f044f027100bafe58fdaefc89fcaffc39fde0fd72fe1bffacff;
    inBuf[9962] = 256'h0f008b001601b401aa02c103cd04f4050e071c0882093a0b270d480f36119212;
    inBuf[9963] = 256'h601394134b13ef129e124f121d12e911a01179119411fc11bd12a5136114c914;
    inBuf[9964] = 256'hd514a4148814ce149315bf160a181c19b219b7195c19f318c3180a19c619a31a;
    inBuf[9965] = 256'h551b921b091bcc191e181a1604141d124210790ede0c3d0b9309fe0744065804;
    inBuf[9966] = 256'h5f023a000afe17fc5efa04f945f8f2f7f5f740f85ff814f867f752f631f59af4;
    inBuf[9967] = 256'hcbf4f7f519f8b0fa4efda8ff7701c302c303940459052106d8067607ef074908;
    inBuf[9968] = 256'ha20808098e09370abf0af20aa00a8b09de07f8052004c8022d02040213021702;
    inBuf[9969] = 256'ha601da00070045ffd3fecbfeccfe9dfe37fe79fd96fce4fb5ffbf3fa7ffaacf9;
    inBuf[9970] = 256'h62f8cff624f5b6f3d8f28af2b8f245f3f4f39cf427f570f560f5edf402f4bbf2;
    inBuf[9971] = 256'h52f1f7eff4ee86eeabee4fef40f021f1c5f11df223f20ff209f2f5f1c5f156f1;
    inBuf[9972] = 256'h75f05fef7fee1feeaaee33f032f22bf493f5d5f507f594f3cdf160f0c2efd9ef;
    inBuf[9973] = 256'hacf01ff2bdf37df556f7e4f819fad8fac5fa13fa2af93ef8d6f733f8e2f885f9;
    inBuf[9974] = 256'h95f976f84ef6a3f3e9f0e4ee00eeefed6cee0fef51ef4bef43ef48efa5ef4cf0;
    inBuf[9975] = 256'haff098f0f2efa1ee29ed17ec7ceb6beba5eb79eba4ea25e9f9e6a6e4aae214e1;
    inBuf[9976] = 256'h11e0a2df79dfaadf55e05de1e5e2d7e4ade623e8e2e88de86de7f2e56be47fe3;
    inBuf[9977] = 256'h6ce3dae3a1e45fe59ae593e598e5c7e595e6f3e746e94aea9aeadae989e824e7;
    inBuf[9978] = 256'hf0e581e5d0e545e6b3e6c8e637e681e516e512e5c5e5fce619e8f4e86be96ee9;
    inBuf[9979] = 256'h90e939ea67eb2fed3feff6f01ff2a0f274f20ff2c2f1a1f1cff11cf232f209f2;
    inBuf[9980] = 256'h9cf1f6f071f032f01df02cf019f098efc5eebdeda7ecddeb64eb03ebb1ea47ea;
    inBuf[9981] = 256'hb3e95ee9a6e9afeaacec58ef0ff267f4fff5a4f6c4f6dff648f761f814fae8fb;
    inBuf[9982] = 256'h91fdbdfe36ff46ff20ffc7fe65fedbfdebfcc7fb98fa7bf9ccf87cf82ef8bff7;
    inBuf[9983] = 256'he2f65df58df3c4f129f01bef9fee6aee74eeaceef6ee92efacf02df20ff415f6;
    inBuf[9984] = 256'hd2f715f9cef9fef9e7f9c9f9bbf9bef9b3f96af9caf8d3f7b4f6b6f510f5ecf4;
    inBuf[9985] = 256'h56f519f6f8f6bcf729f82cf8d6f728f73bf62af5f2f3a0f25df13ff076ef3cef;
    inBuf[9986] = 256'ha5efc2f08ef2cdf445f7b8f9e2fbb3fd3fff9f000f02ae0361051707a708cf09;
    inBuf[9987] = 256'h990a290b8e0b030cab0c620d150e9f0ec00e870e220eb70d9e0d090ed40ecf0f;
    inBuf[9988] = 256'ha910f7109810980f140e530c7d0a9d08c706f80453033202d1015e02f3033106;
    inBuf[9989] = 256'h9e08d00a490cef0c130df00ce90c5e0d240ef70eb00fee0fa30f320fd00ec60e;
    inBuf[9990] = 256'h660f7910a511bb125a135e13041365129911cd10db0fab0e660d2b0c3f0b030b;
    inBuf[9991] = 256'h870bb00c4c0ef80f7811bb12b51385144b15f31584160817561777177f174417;
    inBuf[9992] = 256'hda166816dd155e151915e114ac148b143d14c4135713cd122f12b8114111ca10;
    inBuf[9993] = 256'h811027108a0fac0e400d430b1b09ef060a05db03460322036c03d2033304c204;
    inBuf[9994] = 256'h7b0583062908530ae70ccf0f80129414e9154816ec156e1516153215f8150817;
    inBuf[9995] = 256'h0c18ee187a19bd19ff19291a111aa1199918fe1628154f13a0112a10ae0e050d;
    inBuf[9996] = 256'h430b99096b08f9072208a6082d096d098f09e309870a910bc50c9b0ddb0d820d;
    inBuf[9997] = 256'h9d0c7f0b570a030996073406fc045f04b104bd0533079b084a090509e5070f06;
    inBuf[9998] = 256'hf2030302700067fff1febffe8afe1cfe49fd53fcaafb9ffb5cfc91fd80fe82fe;
    inBuf[9999] = 256'h3bfdd2fa21f826f68ef599f6cff84ffb70fde1febeff86008b01bd02c3031a04;
    inBuf[10000] = 256'h82033a02d900150062009e014703ab0426058204e902b50066fe58fcbbfaacf9;
    inBuf[10001] = 256'h14f9c7f8c4f80af9a6f9cbfa7cfc71fe4b0099010f02d2014101be0087008100;
    inBuf[10002] = 256'h5100c5fffefe68fe8cfeb2ffa501b803240574059a04fa023701b9ff8dfe98fd;
    inBuf[10003] = 256'ha4fc97fbaefa48fa9dfabbfb5afdf4fe1b00a200970052002e003d0053002100;
    inBuf[10004] = 256'h44ffa2fd91fba3f976f89df839fae3fcfcffc5028a041605ae04cc031103ef02;
    inBuf[10005] = 256'h4903be03e30361035d026c011601a101ed026204510556056f04f3024901a3ff;
    inBuf[10006] = 256'hf9fd17fcd7f95ef713f567f3b5f20cf31cf466f56ef6cff66ff675f528f4e0f2;
    inBuf[10007] = 256'he7f15cf14df1c3f1bef247f45ff6d9f85bfb7afdd7fe44ffdefef9fdf4fc0bfc;
    inBuf[10008] = 256'h4efbacfaf9f922f93cf866f7bdf665f651f64ef634f6d9f524f544f475f3e4f2;
    inBuf[10009] = 256'hc7f20df375f3f1f384f43df56ef639f84ffa46fc87fd8afd4bfc1efa93f76cf5;
    inBuf[10010] = 256'h26f4def387f4caf53ef7b5f810fa4ffb9cfce9fd0bffe0ff2000b2ffe0feeafd;
    inBuf[10011] = 256'h13fdaafc9dfcaefcccfce4fcf6fc2dfd88fddcfdf7fd99fdb0fc61fbe2f97af8;
    inBuf[10012] = 256'h64f7aef64df633f63ff659f679f6a1f6d8f62ff7b7f765f81ef9bff923fa27fa;
    inBuf[10013] = 256'hcaf927f970f8e5f7cbf752f876f9ecfa50fc31fd45fdb0fce3fb57fb7afb4efc;
    inBuf[10014] = 256'h58fd14fe22fe69fd68fcdbfb43fcd9fd5100ed02f204d6056d0505040f02e7ff;
    inBuf[10015] = 256'hd2fdbcfb61f9bbf6ebf34ef190ef39ef68f0dbf2ddf593f85bfa0bfb0efb29fb;
    inBuf[10016] = 256'h19fc45fe6d01b1041007bf078806050437010aff04feeefd10febcfd8efcb1fa;
    inBuf[10017] = 256'hd9f8a6f763f7faf7e1f88ff9daf9e1f913faf3fa9dfce7fe880108041c06df07;
    inBuf[10018] = 256'h6909d00a380c840d790e0f0f3b0f010f960e080e4a0d740c8b0b8b0aa409f108;
    inBuf[10019] = 256'h5f080a08060860085909150b750d4e103c13d215ec1773196c1a0b1b491b0c1b;
    inBuf[10020] = 256'h661a371970174215ac12d30f3e0d3e0b360a950a140c1b0e271067117811bd10;
    inBuf[10021] = 256'h900f6b0eea0df60d400eb30e190f900f96104f12ba149917191a9b1be51bce1a;
    inBuf[10022] = 256'hbe18711645149a12c1118e11e111a81279132114a514f8145b15261640176d18;
    inBuf[10023] = 256'h4b1945191f1811166d13af10380e040cff09130825065c04f202fc01a001f901;
    inBuf[10024] = 256'hf7028c0484066408c5094e0ac6097908e70666055804d5037a03090360023f01;
    inBuf[10025] = 256'hd1ff7efe63fdcdfc19fd2efef7ff5602bd04b306f20719082f07a605cd031c02;
    inBuf[10026] = 256'h09018600640076005f0004008afffdfe8afe5afe5afea2fe6effd80013033106;
    inBuf[10027] = 256'hd809900ddd1035135f147e14ca13a012691154106b0f9a0ea10d3f0c4f0aca07;
    inBuf[10028] = 256'hd404c201f3fec8fc98fb8ffba9fcb9fe62013704e9064a09420bd60c020e9a0e;
    inBuf[10029] = 256'h740e8a0dfe0b1d0a3d088506d904f2029800cefde6fa6af8d1f643f6adf6caf7;
    inBuf[10030] = 256'h3cf9ccfa6dfc0bfe9dff2001920203047d05e70602086c08cd071c06ab030901;
    inBuf[10031] = 256'hc5fe22fdfafbe9fa83f9a5f78bf59df352f2e0f131f22ff3bbf4b4f627f9f4fb;
    inBuf[10032] = 256'hacfe0501ca02de0398044105aa058c058204390221ff15fcccf9bdf892f853f8;
    inBuf[10033] = 256'h77f7fff57ff430f4bbf598f8b8fbc8fdd5fd53fc80fa61f99df9d2fab9fb72fb;
    inBuf[10034] = 256'hdef972f74af54cf478f455f52df646f67bf5fbf3d9f132ef0aec60e8a1e477e1;
    inBuf[10035] = 256'h65dfdadec7df97e1d4e326e638e807ea7feb47ec4aecb3ebe5eab3eaa9eb99ed;
    inBuf[10036] = 256'hfbefd3f122f2eff0d4ee91ec22ebdcea3febfaebc7ec68ed31ee3eef1ff09df0;
    inBuf[10037] = 256'h7cf097ef89eed7ed83ed99edc3ed84ed2ded28ed9cedbdee21f0e8f0cff0e1ef;
    inBuf[10038] = 256'h56eee5ecccebaaea46e975e74de599e3fce26fe392e47ee541e5c8e396e179df;
    inBuf[10039] = 256'h6bdebcde05e0cde17de3b5e4ace59fe695e7a6e8afe96cead4eac2eaffe998e8;
    inBuf[10040] = 256'h9de667e4d4e284e28ce3abe5e3e7fbe8a0e833e78de5f4e4fae524e8aceaaaec;
    inBuf[10041] = 256'ha8ed41ee51ef57f17df412f802fbe2fcb6fddcfd1bfeb1fe3cff68ffcbfe37fd;
    inBuf[10042] = 256'h2cfb23f95cf734f6aef5a8f543f65af782f86bf99ef9d5f879f714f61af5f6f4;
    inBuf[10043] = 256'h79f50cf667f675f64cf65ef6cff632f713f711f60ef4a1f1afefcfee34ef80f0;
    inBuf[10044] = 256'he3f1ccf218f310f375f3e6f473f7e3fa94fe9f0188032b04920327025e0065fe;
    inBuf[10045] = 256'h6afc68fa31f8ccf538f37ff0f8ede9eb89ea3cea0feba9ecb7eea7f0dcf146f2;
    inBuf[10046] = 256'h0cf25af185f08fef3bee8aecb5ea42e9fbe84beafcec5cf05df33bf5f5f50ef6;
    inBuf[10047] = 256'h6cf6ccf71dfab6fcb4fe3eff18fec2fbfff89af618f583f4b6f486f5cff697f8;
    inBuf[10048] = 256'hbbfad2fc77fe4eff2fff7efed1fd8efdf6fdecfe0d002d013a021d03e1036204;
    inBuf[10049] = 256'h64041904f3036704d7050a081f0a470b130bd709c5080509100ba80eb212f215;
    inBuf[10050] = 256'hf817e01824197319d519ef19ca19a619231a341cf71f9024c428072b652a3627;
    inBuf[10051] = 256'h5322da1cf8171a14601120105610e511af14db17871a811cd31d171f30211124;
    inBuf[10052] = 256'hf426e228b92842267f22951e9d1b281aa4195c192319f3186019131ba81d3e20;
    inBuf[10053] = 256'h05221f2295205f1e451ce31a711a6f1a811aa71aca1a101b6f1b3f1b2f1a7618;
    inBuf[10054] = 256'h5916aa1424146314b2146e140113dd10360fc50ec00fab1132137b13a8125b11;
    inBuf[10055] = 256'hb21071112913ee14cc1508150413c610ef0eec0db10d860d280df20c210d1a0e;
    inBuf[10056] = 256'hf70ff011321358134b12b910a80f910f87100012d2124e125f10340dbf091907;
    inBuf[10057] = 256'h9e05650538063d07dc07ee0756078a065a064707b109890ddf119315a8176417;
    inBuf[10058] = 256'h2115fe11ef0ea30c110b36094b0673028cfe4cfc4efdb8016108510f4e143916;
    inBuf[10059] = 256'h841576138611a910ae10af10bf0f540dcf094306d7037d0371050109110d6a10;
    inBuf[10060] = 256'hfa118211880fc80c2a0a64087c0736075507a207480892096a0b770dff0edf0e;
    inBuf[10061] = 256'h7c0c1a089d029dfdbafa8afa8efc6cff61016401acff54fde4fb5ffc8dfe5d01;
    inBuf[10062] = 256'h7a03f6030203a201ed0094016a037f05d906d00671058303f7016e0113026703;
    inBuf[10063] = 256'h70044c049f02d6fffefc4afb96fbc9fdcc004d035404b30350027001c4012f03;
    inBuf[10064] = 256'hbc0409055403e3ffc1fb58f8a8f6d4f65af865fa40fcc7fd37ffce00af02b404;
    inBuf[10065] = 256'h67064d0702074c053a020bfe27f93ef411f033ed03ec6cecd5ed8cef12f138f2;
    inBuf[10066] = 256'h6af35cf571f891fc1701df04f206e906fe040e0229ff1dfd77fc53fd45ffb201;
    inBuf[10067] = 256'hce03c30431042a022bff0efc4df9c2f614f4c8f0c8ecf2e86be60be625e80cec;
    inBuf[10068] = 256'h82f0aff435f82dfb04feaa0089021f032202d9ff49fd3bfbcef9b4f841f7f4f4;
    inBuf[10069] = 256'h24f2a8ef47ee52ee55ef6cf0eaf0b2f03ff052f046f1e4f2a7f412f61ef746f8;
    inBuf[10070] = 256'hf3f900fcb2fdf4fd06fc35f8c2f336f09feeedeefaef6ef082ef66ed31eb04ea;
    inBuf[10071] = 256'h62ea2cecc5ee96f185f48ef765fa8ffc66fda6fc07fbcff914fa22fc03ff1201;
    inBuf[10072] = 256'h39017cff11fdc2fb6ffc8dfeb60060010b00d9fd7efc1bfda9ff9302b003ef01;
    inBuf[10073] = 256'hc2fdd7f874f5fef436f7d4fa41fe560007010401ea00f200d000e7fff5fd34fb;
    inBuf[10074] = 256'h1bf84ff542f308f2aef134f25ff3c8f4d3f5c8f57ef484f2d9f092f004f25df4;
    inBuf[10075] = 256'h43f68af6fcf4d5f2f5f1a6f3fdf780fdca0125033f0125fddcf80ef614f55ef5;
    inBuf[10076] = 256'hcef56ff559f452f312f30ff409f623f8b9f99dfafdfa64fb32fc45fd4dfee5fe;
    inBuf[10077] = 256'hd0fe3cfe6afd80fc9dfb96fa28f955f71cf56af25fef11eca8e8b0e5d0e377e3;
    inBuf[10078] = 256'hcfe479e7aceac4ed6ff0d8f280f5a8f811fc09ff9f00510089fe48fcccfaeafa;
    inBuf[10079] = 256'h50fcdcfd4ffee2fceff9def61ff56cf578f7fef9b3fb29fce9fb22fcd2fdf000;
    inBuf[10080] = 256'h89045f078d0824080207080695055f05c6047903c2015300ccff10004f009dff;
    inBuf[10081] = 256'h64fdcff9f6f504f390f1b0f1ebf28ff46ff6d1f8fdfb1100b004ef08e60b010d;
    inBuf[10082] = 256'h3e0c450afe073b06a30553060008540ace0ce10e5b1033118411ba112a12de12;
    inBuf[10083] = 256'had131f14b01348121f10ab0d860bdd0990088507af0667065507b609340dfe10;
    inBuf[10084] = 256'hd713f2148614601384128b12e9125a12b90fa00a11040efe6bfa2cfaf0fcec00;
    inBuf[10085] = 256'h4304f205ec05430575053907620a1f0e4b11471336148614b214d4145b14ba12;
    inBuf[10086] = 256'he30f3c0ccb08b9066b067b0717093f0a730a110ae2099a0a7a0c130f9f117613;
    inBuf[10087] = 256'h411415143513a7114c0f0e0c12080304df005fffdaff0b0209050408890a510c;
    inBuf[10088] = 256'h5e0db00dec0cd00a790752033fff2cfc66fabbf997f94ff9dbf8c5f889f971fb;
    inBuf[10089] = 256'h2efea100bf01340164ff5ffd69fc23fd5aff3802b8044506f00649071e08ef09;
    inBuf[10090] = 256'h8d0c460f1e1128111f0f950ba70797045503fd03e5051908e9093b0b830c550e;
    inBuf[10091] = 256'hdb108d13381596140111bd0a0503bafba9f6dcf447f6b8f954fd61fffcfe86fc;
    inBuf[10092] = 256'h84f9bcf73df8c4fad0fd6fff63fee8fa96f66ff3cbf2acf4c9f78afa26fcedfc;
    inBuf[10093] = 256'he7fd170092034c07cb09250a90082e065304b903080423040f03a30084fdb7fa;
    inBuf[10094] = 256'h02f97ef8c1f864f96ffa3efc09ff7c02b0058f07a407790623058d04d004f304;
    inBuf[10095] = 256'ha703520081fbb6f681f356f256f213f289f001ee3aec42ed15f212fa3d032e0b;
    inBuf[10096] = 256'h4f106f124f12e610c30efd0b9708ed04bf01c2ff14ff2eff57ff2dfff8fe8dff;
    inBuf[10097] = 256'h5f01db039005db04e6007cfa9ef36dee2eec8ceceaedcceebcee66ee5fefe3f2;
    inBuf[10098] = 256'hbdf871fff6049a07060751041f01d1fecbfd4bfd0ffc26f973f4edee2eeab8e7;
    inBuf[10099] = 256'h74e84cec33f28ef8a6fd3b00020088fdfef9e4f60ff53df495f3eff180eee8e9;
    inBuf[10100] = 256'he0e522e4cae57fea3df0aef45ef65ff582f333f3e1f55ffbbd0121069c060603;
    inBuf[10101] = 256'hdefce0f668f311f3d0f470f6a2f59bf15deb1ee56ee1aee144e544ea38ee5bef;
    inBuf[10102] = 256'hcced1aeb3ce9bbe9a8ec81f06bf3eff39cf16eedfee89ee51fe46ce4a4e5eee6;
    inBuf[10103] = 256'hbae7d8e7c7e74de8f8e9f8eccbf062f4c2f65ef768f6e9f4e0f3c3f380f454f5;
    inBuf[10104] = 256'h6ff5e3f464f4c2f49cf69af95dfc70fdeafbe4f7b1f200ee0aeb5eea86eb80ed;
    inBuf[10105] = 256'haceff1f18ff413f895fc6d01990518086908ea066804a401f0fee4fbe7f7f1f2;
    inBuf[10106] = 256'habed73e9e4e7b6e960ee73f40ffad6fd92ffdeffafffcaff30005300b9ff3efe;
    inBuf[10107] = 256'h33fc64fa9ef945fa5dfca0ff90039f073d0bc90dc20e000ecf0be2080706c303;
    inBuf[10108] = 256'h14029e0011ff92fdc3fc55fd75ff6d02c604fe04660299fd3ff83ef4e4f269f4;
    inBuf[10109] = 256'hedf718fcbcff1a02fb028f0235017bff25feecfd2cffb101ab04f406af07ca06;
    inBuf[10110] = 256'h0d059b035a036704fc05fb06aa0619052803f501fc01cb024b0358028dffc1fb;
    inBuf[10111] = 256'h8af857f7a2f89dfb87fe9fff1afe8ffa8bf6def3cdf364f697fae9fee2019302;
    inBuf[10112] = 256'h0c0130fe40fb86f9ccf9e7fbf0feb1012d035903150371030c05870743096208;
    inBuf[10113] = 256'h1b0413fd68f5fdefbaee8bf1baf69afbd0fdd3fc03fab2f712f8fbfb6002f208;
    inBuf[10114] = 256'h3f0de70d4f0b2d07ae0367027f03ed055808cd09730a650bb20dc71122172a1c;
    inBuf[10115] = 256'h231f1b1ff41b89166d10ff0a1207d304ab03b802580148ff15fddafb53fcbffe;
    inBuf[10116] = 256'hab02a7065509510aee0926094809c00ae90cb10e090fb30d950bfd09110a2d0c;
    inBuf[10117] = 256'h480fdc11dd12d611690f120dcb0bca0bd20c2e0e8b0f7f11b9149019a61f7225;
    inBuf[10118] = 256'h2429be292c278022631dc918d5142c113e0d3a091d06ce04d505dd087e0c810f;
    inBuf[10119] = 256'h7f11871242134e14481568153314b511ef0e4d0d8b0d8d0f55125d14e3141214;
    inBuf[10120] = 256'h53124810400eba0b6908c4049401e4ff85002303b106300a140dad0fbd128116;
    inBuf[10121] = 256'h701a421d6c1d611aea147f0ece08d5045a02ab005cff6cfe76fef8ff7602d604;
    inBuf[10122] = 256'hf3053e0577034702f902d605d109f80cd40d210cc608640537037c02dc02c203;
    inBuf[10123] = 256'hb404d4055007b30838092a083805070110fdc9faeffa32fd7900a2030906bf07;
    inBuf[10124] = 256'h5409180bbf0c9c0d070ddd0ad6072605c403fd035e05ea06bf078e078f064305;
    inBuf[10125] = 256'h1c043403630274014900edfe92fd65fc81fbedfaabfabcfa0ffb8cfb3cfc26fd;
    inBuf[10126] = 256'h49feb2ff3e018d02450328032a02a20014ffd8fd08fd7ffce8fb1bfb56fa2bfa;
    inBuf[10127] = 256'h39fbbafd29014d04bf057f04a30095fb76f70ef615f8d3fc58028f065408bd07;
    inBuf[10128] = 256'hd205f503f902db0227037603c1036a04c1058107cf089b0843062a029dfd40fa;
    inBuf[10129] = 256'h5df943fb0dff1403b105c405110354fedcf80af4e2f0bdef5bf025f268f4a9f6;
    inBuf[10130] = 256'hbef887fad0fb70fc49fc7afb75fab6f971f95ef9d6f852f7cef4eef1deefa1ef;
    inBuf[10131] = 256'h7bf103f55df98dfd0b01bb039b05a4069f065405f9020b0027fd01fbf8f9e5f9;
    inBuf[10132] = 256'h94fad0fb45fda6fe91ff87ff4cfe0dfc54f9e4f624f5edf3e0f29ef13af09cef;
    inBuf[10133] = 256'hc2f0e9f376f8d9fc15ff1afe38fabdf477efb2eb8ae978e8fbe7f0e7fbe8feeb;
    inBuf[10134] = 256'h0ef152f746fd5b01ee02920293013801d1018b023a02fcffe0fb43f7cef37ff2;
    inBuf[10135] = 256'h7df3e9f561f812fae4fa12fbdefa0afa02f89af444f041ec59ea7aeb3bef6cf4;
    inBuf[10136] = 256'h6af9ebfce7fe00009900910025ff7dfbc6f559ef32eafde7eee899ebeeed4eee;
    inBuf[10137] = 256'h88ec29ea55e983ebd7f0f1f7abfe5d033f0586043f0272ffe0fc3efbd0fa45fb;
    inBuf[10138] = 256'h13fc6bfc80fb48f986f66af40af476f5b1f771f9acf957f8bdf64af693f73efa;
    inBuf[10139] = 256'hf7fc3cfeb3fd3dfc47fb03fc6ffe39018c020701a6fcd6f67df138eed4ede7ef;
    inBuf[10140] = 256'h5df348f7e4faa9fd52ff9fff7afe47fcc6f9cdf7f4f61ff7aef7faf7c9f7a2f7;
    inBuf[10141] = 256'h82f81afb4fff0f0498077a084c06b20131fc6af715f4f9f152f028ee31eb4ee8;
    inBuf[10142] = 256'he0e627e8c2ec0af43afc4c03b007ea08c507b3052a04040400053606d1068906;
    inBuf[10143] = 256'h020687061b09cb0d78132918281ae21815156710420ce4087905c4001efa57f2;
    inBuf[10144] = 256'h72eb80e795e712eb03f052f4c5f694f721f8aff984fcd5ff1102e7015bffb7fb;
    inBuf[10145] = 256'hdbf861f897fa56fed201860301034401fcff82002e030907660af50b5a0b5d09;
    inBuf[10146] = 256'ha2079e07e309030eaa124016be17e3164b144611130f530eed0ef70f2710a90e;
    inBuf[10147] = 256'h780b800734049302b302bc0338042503b100eafd4ffcfdfcd1ffbe0391074d0a;
    inBuf[10148] = 256'hcf0bb70c830d650e500fe60f0c100210c60f220fc20d1e0b47074b037b00f3ff;
    inBuf[10149] = 256'h160211066b0ae60dfe0f28115212fb13db15ed160316c7120d0e5f0977063306;
    inBuf[10150] = 256'hfe07720a160c070c9b0af8082308ad08650a5e0ccf0d6a0e110ef40c5f0b6f09;
    inBuf[10151] = 256'h6607bd05d9040f05520602089609ce0a930b330cfb0cae0dea0d620df80b1b0a;
    inBuf[10152] = 256'h7c08590790069c05b803a200dbfc42f9ebf68af60bf8d2fa11fe1901b2030d06;
    inBuf[10153] = 256'h9408a10b0b0f4012921420154d13450fc309e0030fff7afc87fce8fe9a023d06;
    inBuf[10154] = 256'hbf08b3096909c808ab086e09b80a850bb90ad30704031ffd55f77af2b0eec8eb;
    inBuf[10155] = 256'h89e9fde7bee79ce9feedaff4b5fc81049d0a2f0e110fd60d820b1a094007f405;
    inBuf[10156] = 256'hcb044a032601a0fea3fc20fc81fd7300e80383067407dc069e05cb0410055a06;
    inBuf[10157] = 256'hdc07aa087f08ba07f606dd068f074208da0793054401aafb3df68df29cf16df3;
    inBuf[10158] = 256'h14f721fb2efe71ff17ffeffddffc83fccdfc0afd6efc94faaff797f470f219f2;
    inBuf[10159] = 256'hccf315f707fbb0fe7f016f03d80413062707bb0742077805c7020f004afe3bfe;
    inBuf[10160] = 256'hcafff801a5030d04f902ff0026ff2efe61fe97ff4c01fb023604ad0456044703;
    inBuf[10161] = 256'hca017500b5ff7fff84ff1cff8bfdc3fa49f7c8f3d2f086ee76ec34eac5e7bfe5;
    inBuf[10162] = 256'h0ee551e673e9b0edd3f1e2f4a6f67bf709f8ddf8ebf9abfa80fa01f95ef670f3;
    inBuf[10163] = 256'h2ef15cf038f110f3bbf45ff59bf4ddf272f189f16ef3aaf6fbf9d7fb91fb81f9;
    inBuf[10164] = 256'haff679f4d6f3d4f4e6f62ff9e5fad4fb29fc4bfcd4fc1afe00002102a2037303;
    inBuf[10165] = 256'hf10015fc8df5c7ee1fe94be554e398e258e279e287e346e632ebedf136f990ff;
    inBuf[10166] = 256'hea032a061c07aa07440892087907ee03ddfd52f642efd3ea52eaa6ed64f350f9;
    inBuf[10167] = 256'h64fd99fe10fd03fa32f7e4f597f62af9ccfc8a00fa0300078209790ba00c5e0c;
    inBuf[10168] = 256'h520aaa061602b4fd9afa66f905faa6fb3afd0efebffd61fc87fab7f825f7f5f5;
    inBuf[10169] = 256'h19f548f45ef34df21ff134f01ff066f161f4def804fecf027506b308f9091c0b;
    inBuf[10170] = 256'ha60c620e6d0faa0e540b780511feabf6abf0e7ecb0ebc9ec9aef7df3c5f7a8fb;
    inBuf[10171] = 256'h81fef3fff7ffe9fe41fd5efb8af9f6f7d8f6b1f6f9f7b2fa62fe100285041005;
    inBuf[10172] = 256'hd903ab0188ff0bfe0efde5fbcef995f6d8f285ef53ed9bec17ed47ee1bf0eef2;
    inBuf[10173] = 256'h12f762fce9011f06c20785066e035400aafec5fed1ff3100acfe4ffb35f7baf3;
    inBuf[10174] = 256'hd2f17cf1f9f1a4f278f3f7f4a0f73dfbb0fe8900fcff86fdd2fac9f976fb4fff;
    inBuf[10175] = 256'h85032c06570681043a02100174019002f4026501aefdbef807f4b6f04defa7ef;
    inBuf[10176] = 256'h4df1baf384f64ef9a7fb3ffd58fea4ffe601af05bd0adf0fdb13091697167616;
    inBuf[10177] = 256'h7c168f16be15c9120a0d5b05b5fd3af849f6aaf7befa9cfdedfe70fefefcc7fb;
    inBuf[10178] = 256'hbbfb51fd5600450496089b0cab0f65119b118010a70e730c0c0a6a074504b800;
    inBuf[10179] = 256'h8dfd9ffb89fb6bfd63001603b0040805a0046c04ea04d705b4063007a7072f09;
    inBuf[10180] = 256'hb70c38127818481dc01e651c4e17ca113c0ea20d670f0f12dc13fd13fe12dd11;
    inBuf[10181] = 256'h7511161201131a13c611f80e5f0b2b0825068b050d06ba06b606b505e4033102;
    inBuf[10182] = 256'he20192033007e80b08102612e711ac0f980c130abe087808cc08180927094709;
    inBuf[10183] = 256'hb709950abd0ba70cfc0cde0c890c750c1b0d720e3d103712e5130115ac150916;
    inBuf[10184] = 256'h6b165117b418251a071b7b1af817c813b20ec009f105a2039f026c0272026e02;
    inBuf[10185] = 256'h5f0246025402b30254035504e105d707340af70cd60faa123d15fb168417b116;
    inBuf[10186] = 256'h8114ac11430fd20d860dfa0dee0d460cb4088803d3fd12f943f69ff5a7f653f8;
    inBuf[10187] = 256'hc0f9adfa88fb4efddf005106d70cfc123017ac18ad173715ae12f9102110c40f;
    inBuf[10188] = 256'h4d0f3f0ec90c710b830a280a3c0a0c0ad208040653010ffb4bf48aee56eb9deb;
    inBuf[10189] = 256'h47ef52f51efc1e0285061409cf09ec087f06a60221fe24faeef75ef84dfb97ff;
    inBuf[10190] = 256'he4032d071709240af00a8e0b8d0b400a28076802d5fc9bf7bff3d3f110f251f4;
    inBuf[10191] = 256'h12f8acfc4201d104a0068506d8046102d3ff6ffd2afbb9f8e7f52af354f1edf0;
    inBuf[10192] = 256'h38f2eef4fcf74ffa74fb5afb62fa52f9a5f84df815f8baf707f721f682f5a3f5;
    inBuf[10193] = 256'hd7f644f9b7fc940003041f0613068603e2fe1cf961f3aeee37eb67e88fe55ae2;
    inBuf[10194] = 256'h34df60dd26def2e105e8b0ee4bf452f878fb45ff1505a00cf2139f18d3187d14;
    inBuf[10195] = 256'hc60d9007cf03be02ae022201a2fc85f5b2edabe70ae5e1e534e98fedebf137f6;
    inBuf[10196] = 256'h9cfaf6fef60222060a08e1082109bd082807bc032ffe51f72bf1e8ed8eee6af2;
    inBuf[10197] = 256'h4af7a1fa1dfb6df996f784f7cff94cfdcbffb8ff2cfdb8f955f713f72ef8bef8;
    inBuf[10198] = 256'h38f76cf3c1ee90eb8aebc6ee08f482f9fbfd580104044a061108ab089c076b05;
    inBuf[10199] = 256'h1f039e013e013c014600e5fdd0fa8af8bef8dffb81006304b105ee0371007cfd;
    inBuf[10200] = 256'h9ffcf2fd2c00880116014fff8bfdfcfcc3fdc8fe94fe4ffc68f865f4bef1dff0;
    inBuf[10201] = 256'h1df105f156ef16ec61e89be5e3e45be627e95eec81ef7af28ff5daf8fbfb89fe;
    inBuf[10202] = 256'h5900b80184036206240aef0d6e107510e30d7c0961048eff2efbaaf66cf158eb;
    inBuf[10203] = 256'h11e5f9df4edd88dd52e096e425e975ed94f1e2f5c1faf8ff970494072208ff05;
    inBuf[10204] = 256'hb20139fc98f6aef10ceef6eb76eb56ec23ee3ef007f243f339f46ef57bf7b5fa;
    inBuf[10205] = 256'ha4fe5302ed04dc0526059c0317021201b0007b00b7ff1efed9fb79f9f2f7e5f7;
    inBuf[10206] = 256'h3ef981fbd5fd64ff13006300f4003f022704dc056e066105fe02500094fe91fe;
    inBuf[10207] = 256'h3f00cb020305fe058105eb03df01f5ff5dfec2fca6fabcf7f9f3afef78ebe6e7;
    inBuf[10208] = 256'h61e545e4c6e405e716ebbcf04af7d6fd5f031807c208a1082907d9040f02f4fe;
    inBuf[10209] = 256'hc3fbf7f813f781f668f77bf93efc5effc0028306c90a330fe912f9149814ab11;
    inBuf[10210] = 256'h250d6d08c104df029302cc026c02f10093fe32fcd7faf9fa23fc4afd64fd09fc;
    inBuf[10211] = 256'hbef9b6f729f79ef88dfbaffebe00f4005effe4fca3fa2ff979f8f7f7d9f6b0f4;
    inBuf[10212] = 256'he7f18eef04ef6af1ecf683fe4306f60bfc0d0f0c4a07a8013afd2bfb56fb93fc;
    inBuf[10213] = 256'h5ffdadfc89fa1bf805f7b8f89afdb2040e0c84118a130f126b0e930a3108d307;
    inBuf[10214] = 256'h9508dc086f072d04290008fd0efc5efde4ff30025a034203a20286026303ee04;
    inBuf[10215] = 256'h91069a07ae07080717063305a1047f04eb04020694071b09e609450922074604;
    inBuf[10216] = 256'hf8016d0113032e065509360b4b0b500aac095e0a680cbe0ec40f7e0e550bb007;
    inBuf[10217] = 256'h220582044e052606e10551046f02980172026904fa05a705230390ffb3fcfafb;
    inBuf[10218] = 256'h9dfd7a001f03e3042106fd075e0bd20fb3131315ac12da0c8405f1fecffa82f9;
    inBuf[10219] = 256'h1dfa48fb10fc1afcbefb97fbeafbc7fc28feedff1e02de0409084f0b5a0eda10;
    inBuf[10220] = 256'ha612c5134d14451491130d12af0f770c7e081904b3ffbbfbbff836f741f79bf8;
    inBuf[10221] = 256'hb2fad8fc8afeb6ffc4004b0291046207120aaa0b780b8d0992066e0304019eff;
    inBuf[10222] = 256'hbefeb0fdedfb40f92ef6b8f3b2f2a3f3a8f62ffb3c00c904d507a8081b07a303;
    inBuf[10223] = 256'h47ff40fb91f8cff7e4f81afbaafd0200c801fd02d5035b04870465041204c903;
    inBuf[10224] = 256'hdb037d04a5050c0750081c093e09aa088307f7053204720202012b0033006301;
    inBuf[10225] = 256'he2039107180ce2102015f617cd18791725144d0f96096f0305fd88f63bf08fea;
    inBuf[10226] = 256'h4be643e4eee44ae8c0ed3cf4c2fabc00fc05c70a6f0fc3130c1749189b16df11;
    inBuf[10227] = 256'hca0abf025cfbb9f52ef2a4f0c3f035f2e1f495f8acfc37005e02cf02fd01e700;
    inBuf[10228] = 256'h8a002f0130029202b301bfffd0fd4cfdd6fef90157054c07d9062c044b006afc;
    inBuf[10229] = 256'h5bf939f7b1f576f490f364f357f46af61ff9b6fb75fd04fe8efd87fc7afbd6fa;
    inBuf[10230] = 256'hd6fa99fb0efde8feb500f70131025501f3ffd5fe94fe45ff4000570092fed3fa;
    inBuf[10231] = 256'h0ff6ccf16fef9feff8f16af51af9bafc8800eb04c209210ed210c910b70d6e08;
    inBuf[10232] = 256'h4a0291fc4bf804f6c6f576f7cefa27ff8c03ef0685081c0822066a03ba0075fe;
    inBuf[10233] = 256'hb3fc74fbc1fac9fabafb66fd4dffd7008b0146012e0070fe1efc26f9a1f522f2;
    inBuf[10234] = 256'h96efe0ee75f0e4f3dbf7dffa12fc9dfb91fa51fab5fb89fea201a303e103bd02;
    inBuf[10235] = 256'h6b0150011403310656092a0b070b610970076206c40632088509a6091708f004;
    inBuf[10236] = 256'he50002fd17fa82f85cf863f9fefa85fc95fd2efeb7fed1ffe5019c04fa06e607;
    inBuf[10237] = 256'hb306b0033200c0fd47fdabfed4005e027d02430169ffb7fd72fc50fbc8f987f7;
    inBuf[10238] = 256'hc3f41bf21ff01cef2cef50f09cf22cf6dbfa0b00af04c707ee088b088907c106;
    inBuf[10239] = 256'h6e061206e8049d02ccffbffdadfdf4ffbc034307cd08bc07df04e4016300fb00;
    inBuf[10240] = 256'hd90237049803be00ddfc02faecf9f7fcef01a9063b090109b406c4036801deff;
    inBuf[10241] = 256'h63fefefb56f81cf4c6f0c0efb3f130f6f1fb920131068209af0b110dd70d120e;
    inBuf[10242] = 256'hee0db80dc70d690ea90f25115b12f412c612df118610f20e070d7e0a1d07d702;
    inBuf[10243] = 256'h07fe7df93cf604f5f6f580f894fb1dfe88ff0c0071008b01ac037306fa083e0a;
    inBuf[10244] = 256'ha6095807f8034200c7fcbff92bf71af5bdf36ef379f4c7f6e8f952fd76000703;
    inBuf[10245] = 256'h2105fd06b6083d0a3f0b5c0b6a0a88083606360429036603eb0439077309c50a;
    inBuf[10246] = 256'h960ab2088005df01b0fe9bfcecfb68fc8afd13ff0e019303bb065a0aa90db50f;
    inBuf[10247] = 256'hf90f8e0e220cc1093f08bb07ae076c07910620057b030302b40034ff2ffdabfa;
    inBuf[10248] = 256'h29f853f671f532f5e0f4cdf3f3f12df0b9ef67f10ff59af987fdd3ffa6002001;
    inBuf[10249] = 256'h9f02e605960a570f911236134811c30dfe0907075b05cd04c404b9047304f203;
    inBuf[10250] = 256'h5803c5022102180160ffe2fcbcf974f6e8f3ccf27af3eff591f961fd84007002;
    inBuf[10251] = 256'hfe0274024101b1ffd2fd86fbcef800f6bdf3ddf20cf452f702fcfb001305aa07;
    inBuf[10252] = 256'hd7085109140ac10b2d0ea6103012ef11bb0f490cbc08380673054706c307ac08;
    inBuf[10253] = 256'h0c08a40512026cfeabfb3ffae5f9e2f9c0f9b3f96afaaefcda003f065a0bb00e;
    inBuf[10254] = 256'h6b0fbc0de20a5308c506fb05f2047402fffd3cf892f292ee43eda4eecef18ef5;
    inBuf[10255] = 256'hcdf8e5fac9fbb3fbf4fa03fa5df958f927fab2fb6ffdaffe1affdafe7ffeb9fe;
    inBuf[10256] = 256'hf2ffdb019b0370041504e202ad013701a201880247037b03550365032504a305;
    inBuf[10257] = 256'h540765084708fd061905530312025601c500d6ff65feb9fc1efbdcf923f9c1f8;
    inBuf[10258] = 256'h6df80cf878f796f668f5fdf3a2f2edf177f2aff494f87bfd7f02f806900a510d;
    inBuf[10259] = 256'h6b0f9510f60fb30c84062bfe8df5f8eeebeb5becd5ee49f13af2aaf112f141f2;
    inBuf[10260] = 256'h2cf640fc80028d060f075104e9fff6fbfdf920fa8dfb30fd2dfe63fe61feb1fe;
    inBuf[10261] = 256'h8fff0501ce026d04680542057d03e3ffdafa70f5fcf092ee90ee57f0b2f2a4f4;
    inBuf[10262] = 256'hd7f5c2f644f8d2fa12fe1501b8026802af00a7fe4ffd32fdf3fd89fe36fe0cfd;
    inBuf[10263] = 256'hd3fbbafb9dfd470175057a080709e8062a038aff9cfd0afe4c0013032005cc05;
    inBuf[10264] = 256'h38051904190353025e01a8ffd5fc05f9dff448f1f8ee4bee4fefb6f1e1f42cf8;
    inBuf[10265] = 256'h0cfb11fd29feb4fe22ffabff43008e001d00e3fe6cfd99fc38fda1ff61036007;
    inBuf[10266] = 256'h7c0af50ba40b090aef07ce05c3039f01edfe6afb62f769f31df016ee90ed58ee;
    inBuf[10267] = 256'h11f076f259f598f8fdfb2fffbe014e03de03e503f2035604200504067d065a06;
    inBuf[10268] = 256'hef05ab05cf055006a40602060804f70090fdc7fa5cf979f9b2fa5efc01fe68ff;
    inBuf[10269] = 256'ha80000028703f804d3058d05d003a60091fc6df825f569f389f35ff550f8a0fb;
    inBuf[10270] = 256'hb6fe2b01fc027404df055d07c0087709ea08d10662036dff19fc49fa39fa64fb;
    inBuf[10271] = 256'hd0fc98fd5ffd78fcadfb9dfb5ffc95fda6fe1dff0bffebfe31fffeff1501fa01;
    inBuf[10272] = 256'h3502a1018f0083ffedfe0dffe1ff0801f1012b0283012d00e2fe91fec8ff5c02;
    inBuf[10273] = 256'h64058807b507d705ec026a006afffaff18015601d8ff01fd35fa04f942fa7cfd;
    inBuf[10274] = 256'h2f01bd03620486035d0229027503ce0519084709e8082e07a904e9011eff35fc;
    inBuf[10275] = 256'h36f983f6d9f4fdf43df722fb84ff0203b60490043a03ab018100a3ff7dfe8bfc;
    inBuf[10276] = 256'he6f97ef7b2f684f800fd20034609f80d8b103c11ad104e0f210dcd092305a4ff;
    inBuf[10277] = 256'h70fabaf645f5dff577f7cbf816f968f888f76df7b0f841fb74fe8601f4038305;
    inBuf[10278] = 256'h480689066006c105bb046503c901060048feb2fc6dfbc8fa01fb05fc73fdbefe;
    inBuf[10279] = 256'h4bffd4feb4fd9efc32fcb2fcd0fdd4fe36fff9fea7fe02ff5b0031026803e402;
    inBuf[10280] = 256'h38001dfc22f8bcf597f535f72bf91afa94f934f83ff7e8f770fa0dfe6c016503;
    inBuf[10281] = 256'h9a039b0270010401bd015d034a05f00603088f08c308dd0816096d09b709cf09;
    inBuf[10282] = 256'h5e09eb0746058101e8fc2ff839f4b2f1f9f018f2c7f489f8d2fc2501ff04d307;
    inBuf[10283] = 256'h3c090e096007be040302f3ff25ffcbff8901c803f70585071b08ae073c06ea03;
    inBuf[10284] = 256'h280184fe91fccdfb4afc91fdf2feceffe1ff6cff0dff49ff3900740153025702;
    inBuf[10285] = 256'h6b01f2ff82fe82fdfffcd0fcd3fc28fd1afedaff3d029b040c060906aa048002;
    inBuf[10286] = 256'h6200ebfe02fe28fdfffb87fa41f9edf8fbf93ffc13ffbb01d2036805d2064e08;
    inBuf[10287] = 256'had096d0a0e0a52086e05eb0157fe2efbe9f8e9f78ef81afb4cff4f040c096a0c;
    inBuf[10288] = 256'hc90d500da10b630903077b047d01e0fdeaf94cf6ebf38bf36df536f90cfecf02;
    inBuf[10289] = 256'h68062d0802084b06cc0355015cffe3fd84fca7fadff742f47ff0adede7ecdaee;
    inBuf[10290] = 256'h66f37ef996ff3e04b5063907d206a9065b079e087409de088506010396ff72fd;
    inBuf[10291] = 256'h07fde8fd12ff98ff29ff24fe47fd33fd15feacff8601370383044c057705f204;
    inBuf[10292] = 256'hc00314024f00e0fe12fef0fd56fe16ff16005d01ed02a3042906fe069f06d304;
    inBuf[10293] = 256'hc90103fe42fa4cf7a2f563f561f62bf845fa5efc4efe1000bf016e031d05c906;
    inBuf[10294] = 256'h50086709ac09c70894065603d4ff12fdd5fb4dfc05fe030048015b01670003ff;
    inBuf[10295] = 256'he3fd84fd07fe55ff3a017b03c205840733087d078105df027a00f7fe55fef8fd;
    inBuf[10296] = 256'h17fd32fb83f801f6cdf488f50df861fb21fe52ffd9fe5dfdfffbb8fbbcfc71fe;
    inBuf[10297] = 256'hddff32005dff11fe5efd0efe2f0009039b053007ba07c107e4076108f8081209;
    inBuf[10298] = 256'h3b087f0647040e0224009dfe6bfdaafcb2fcd9fd1500e2028a058307ac086109;
    inBuf[10299] = 256'h140ac00acc0a74093d06690117fcbcf76bf567f524f7a7f914fc03fe7cffbd00;
    inBuf[10300] = 256'hda01a502e0025c022c01b8ff73fea6fd70fdb7fd4dfe2aff6f004602c204b707;
    inBuf[10301] = 256'hbf0a580d090f970f1b0fce0d090c260a54089b06ea041403ee007cfef9fbf0f9;
    inBuf[10302] = 256'h07f9aaf9defb20ff7202d0049a05cb04fc021401e0ffdbfff600b10287040106;
    inBuf[10303] = 256'hcc06ea068e06de05fd040d040703d4017200f8fe92fd8ffc44fcdcfc38feedff;
    inBuf[10304] = 256'h60010902c101da00f4ffacff2e000e018801f60046ff33fde6fb43fc7efeeb01;
    inBuf[10305] = 256'h48057e073808cd07f8065b06ff0563050f04e4014fff20fd01fc0ffce0fca9fd;
    inBuf[10306] = 256'hbffd09fde5fbf2fac3fa82fbe5fc56fe30ff0dffd3fdbefb60f969f75df68bf6;
    inBuf[10307] = 256'he2f7e5f9f4fb9dfdaffe4bffb7ff200073006c00e6ff11ff5ffe52fe27ff8100;
    inBuf[10308] = 256'ha101d901e90031ff8afdabfcb9fc46fd8efd0bfdeafbdafaaafacffb00fe4c00;
    inBuf[10309] = 256'hc7010402490175007800b101ad036a05da056f046f01e0fd09fbc8f94bfa21fc;
    inBuf[10310] = 256'h6efe53005b017701c80097ff31fec9fc8afb8dfac4f913f968f8e4f7e8f7dff8;
    inBuf[10311] = 256'hf8faf8fd3301db037b05210648066a069e068606a005b503330100fff2fd4afe;
    inBuf[10312] = 256'h82ff89006400bdfe06fc38f951f7ebf61df893fad0fd5e01ca04920735095709;
    inBuf[10313] = 256'hef0753052f0252ff3cfd02fc75fb38fbf7faacfa8efac0fa3cfbe8fb8dfc06fd;
    inBuf[10314] = 256'h76fd28fe3dff8f00b9012d02990131007cfe0bfd35fcd2fb6dfbc3fa02fabef9;
    inBuf[10315] = 256'hb4fa38fddd00ab049707f108b7087207b805d103af011cff10fceff869f61df5;
    inBuf[10316] = 256'h53f5e3f655f91ffcd7fe3c011a033a047004c903980260019a006f0096008300;
    inBuf[10317] = 256'hbfff41fe80fc2ffbdefaa5fb03fd33feb8fe91fe40fe8dfee9ff11022a042905;
    inBuf[10318] = 256'h6104f401d1fe32fc06fb86fb2efd1effb200c20185024b031e049a0450042403;
    inBuf[10319] = 256'h7501f7ff4cff84ff0500f7ffd3fec0fc96fa6df9ecf9f8fbd6fe97019203b704;
    inBuf[10320] = 256'h5f05e1055b06a10664067905f9032302420085fe06fdf4fb95fb1bfc84fd75ff;
    inBuf[10321] = 256'h400141023e028401c100a8008d012703b804940565054904c6026d016b0098ff;
    inBuf[10322] = 256'hadfe69fde6fba5fa30fad8fa8bfcbffeb300ce01d7010901f2ff2fff2dff0a00;
    inBuf[10323] = 256'h8c013f039a04220594040103cb008dfee9fc43fc95fc75fd50feadfe66feabfd;
    inBuf[10324] = 256'hd3fc1dfc8efb11fb97fa40fa6afa74fb6cfd0800c002ec0428067a061a064b05;
    inBuf[10325] = 256'h420406038301c5ff06fe8afc8bfb26fb47fbadfb1cfc7cfcc3fc05fd75fd2afe;
    inBuf[10326] = 256'h13ff0900b600b000c0fff7fdb5fb9df941f8e1f75df837f9def90efaf1f908fa;
    inBuf[10327] = 256'he2fac5fc75ff3c023304b20488030601e9fd07fbf5f800f829f833f9d4fad7fc;
    inBuf[10328] = 256'h11ff5c0198038505d20637078b06e404b00293001dffa2fe0bffd9ff77009100;
    inBuf[10329] = 256'h3400d5ff0f003c012f034a05b806c4063e058f0287ff0cfdcefb0efc89fdb7ff;
    inBuf[10330] = 256'hf201a603790458046e032102eb002f002300a30035014c018d0000ff29fdc5fb;
    inBuf[10331] = 256'h72fb63fc42fe8000b102b104ae06e4082a0bd90c2e0dab0b6f0853048900e7fd;
    inBuf[10332] = 256'h90fcfbfb55fb12fa57f8d7f65ff667f7b4f97ffceefe7e002b016c01e001e002;
    inBuf[10333] = 256'h6c044c061e088a095f0a810ad509520815066303950008fe01fc9dfafaf958fa;
    inBuf[10334] = 256'hfdfb09ff3703a507f90af60b170ad905a20026fc9df949f98dfa6bfc2bfeaeff;
    inBuf[10335] = 256'h48014f03b905fd0759095309f907c8056c036a01e7ffc8fee8fd39fdb7fc60fc;
    inBuf[10336] = 256'h2afc13fc3dfce5fc38fe1e000a022b03db02100164fedbfb5dfa17fa61fa34fa;
    inBuf[10337] = 256'hc8f806f6c0f24af0c6ef91f12ef58ef98efd6f002b0233030e041a0558066207;
    inBuf[10338] = 256'hc1072707820511034e00abfd84fb0ffa4ef92af98cf95cfa86fb03fdbffe8800;
    inBuf[10339] = 256'h20024403b50360036f022801d7ffbffef4fd58fdc6fc2afc8efb2afb56fb65fc;
    inBuf[10340] = 256'h83fe910113053e082f0a320a19085a04e7ffcffbdcf845f7c5f6e6f65df731f8;
    inBuf[10341] = 256'ha1f9d8fbbcfee301c3040c07c908300a680b610cbf0c060c0b0a0e079d035d00;
    inBuf[10342] = 256'hc4fde6fb8efa76f97cf8b4f745f755f7f4f710f97dfa1bfccafd4eff5c00bf00;
    inBuf[10343] = 256'h6b009effe8feeafeeaff9a013203bb039502e8ffa1fce4f977f860f8e6f819f9;
    inBuf[10344] = 256'h91f8c7f7d2f7b8f9b6fddc026f07cc093c094c067e0278ff29fe76fe88ff6300;
    inBuf[10345] = 256'h8b0047005300570184036e063609fb0a4a0b290a0508940587034202d001eb01;
    inBuf[10346] = 256'h0902a0017900dbfe65fdbefc42fdb0fe3100da004300b5fe1cfd94fcb5fd2b00;
    inBuf[10347] = 256'heb02c4040405d3031c020e015b01db02ba04e6059505c3032c01cafe5dfd1afd;
    inBuf[10348] = 256'h92fd08feeffd3bfd6dfc49fc57fd84ff1802ff034d04c7020a0048fdbffb27fc;
    inBuf[10349] = 256'h57fe60010f048d05ba052605b304f704cd056f06fb050904070126febdfc7efd;
    inBuf[10350] = 256'h0d003903a2056b06b1056b04ac03f80313052b064f061705ce022a00e0fd63fc;
    inBuf[10351] = 256'hcdfb00fce6fc8dfefe00110460075f0a880c890d580d190cf7091907b2031b00;
    inBuf[10352] = 256'hdbfc84fa8cf915fac1fbebfdf6ff76014b02aa02d002bf024d025301c9fff2fd;
    inBuf[10353] = 256'h61fca9fb0bfc5afd12ff92006f019b0159010601d600be008000d9ffa1fee4fc;
    inBuf[10354] = 256'hecfa26f9fcf7ccf7c8f8c8fa4ffdbcff6e01fd017601520023ff57fe1dfe55fe;
    inBuf[10355] = 256'hbcfe2bffb8ff9200d7017303090516062106ec049d0299ff5efc71f92cf7a3f5;
    inBuf[10356] = 256'hcef4b4f45bf5dbf66af90dfd6501d1058b09ce0b310ce30a6e0878058b02e5ff;
    inBuf[10357] = 256'h6efd09fbdcf858f71cf7a8f8fdfb7100e3041f086009a508a9067204dd023d02;
    inBuf[10358] = 256'h380217025701ebff3ffe09fddffcc3fd2aff6100dd00760093ffe1fedefea0ff;
    inBuf[10359] = 256'hd600f10169020502e90076ff08fed1fcd8fb05fb2dfa42f95ff8a4f727f706f7;
    inBuf[10360] = 256'h4ff7edf7ccf8ddf9fffa18fc31fd59fe97ffec003d024603c503a103f302f901;
    inBuf[10361] = 256'h0d01700026000600e1ff95ff2fffeffe1ffff3ff750175038c0541072a08ee07;
    inBuf[10362] = 256'h7806f903d10077fd75fa32f8d9f67ef622f7adf804fb03fe4b0146044306b006;
    inBuf[10363] = 256'h5a059f0262ffc0fc98fb2dfc1cfe9200ad02db030d048a03a502950175003fff;
    inBuf[10364] = 256'hf8fdbcfcaefbcdfa06fa53f9c7f895f806f947fa41fca7fe170130039c041d05;
    inBuf[10365] = 256'h7f04a902ccff7ffca2f91ff891f8e6fa74fe400256052d07ba07460720067a04;
    inBuf[10366] = 256'h5d02c0ffc6fcd4f976f73df67ef61cf888faf2fc92fe01ff69fe70fdeefc8afd;
    inBuf[10367] = 256'h62fff8017c042a06ac0644069c054f059a052f066606a805dc0388018cffaefe;
    inBuf[10368] = 256'h32ffac003f022e034a03f902f802e003b005bd071509f808380750041a015cfe;
    inBuf[10369] = 256'h7cfc75fb05fbf2fa39fbf5fb38fddffe8300a401f10172018200a0ff24ff0bff;
    inBuf[10370] = 256'h04ffabfeddfdddfc38fc6ffca7fd80ff3a012802120247016a00150074002b01;
    inBuf[10371] = 256'haa018b01d400f1ff7bffccffc900f101b002a402c0014c00adfe30fd04fc46fb;
    inBuf[10372] = 256'h0ffb74fb79fcf0fd87ffea00ed019f023903d70347041a04e4028c0093fdecfa;
    inBuf[10373] = 256'h82f9c4f96ffba5fd70ff50006c005600a10072014f027c026c0125ff4efcdff9;
    inBuf[10374] = 256'ha2f8ddf845fa37fc22fec7ff3801a7023704c90507079a0755073d0677044402;
    inBuf[10375] = 256'he8ffaafde4fbfefa3ffb91fc81fe51003f01e10069ff84fd06fc8cfb2efc7efd;
    inBuf[10376] = 256'hc4fe60ff18ff27fe11fd5cfc58fcf3fcc7fd6efeb6fea9fe8ffec4fe56ff0000;
    inBuf[10377] = 256'h5900100020fff9fd47fd83fdb8fe76000202b60260023f01d6ff9ffec8fd2bfd;
    inBuf[10378] = 256'h87fcc3fb11fbebfae2fb3efecd01ef05c8098f0cdd0dcd0db60ce90a8b087c05;
    inBuf[10379] = 256'h8c01e5fc32f863f456f267f223f476f64af80ff9f5f8d0f88ff99dfba1feae01;
    inBuf[10380] = 256'hc7036f04e003e4026602ed025404fd0537078707de06960515048c02040170ff;
    inBuf[10381] = 256'hccfd36fce7faf7f94ff9c4f84af812f881f8f1f95afc3bffc9015003a3032e03;
    inBuf[10382] = 256'hac02a5021b038c033d03d201a4ff80fd35fc2ffc2afd5afe08fffcfe76fefdfd;
    inBuf[10383] = 256'h02fe84fe1fff7cff91ffa2ff1900220163022303bc02000163fed1fb26fabef9;
    inBuf[10384] = 256'h57fa46fbe5fb00fce1fb20fc45fd79ff6f028a052508c509380a96092a085206;
    inBuf[10385] = 256'h7004da02c3012e01f100cc007900d1ffe5feecfd32fdf8fc54fd36fe6effbe00;
    inBuf[10386] = 256'hef01e3027f03ac036603b4029d014600e0fe86fd49fc46fb95fa56fabdfaf0fb;
    inBuf[10387] = 256'he1fd5700fe0273056c07cd089109b9094f095b08fb06740521044803f702f702;
    inBuf[10388] = 256'hd00200024b00d5fd1bfbcaf884f798f7ebf823fbbefd39004202b9039b04fb04;
    inBuf[10389] = 256'h0205d904a1047704620451042604cc034303a9022302c8018b013c019d008dff;
    inBuf[10390] = 256'h14fe65fcc5fa74f98ef820f83af8edf84efa64fc0bfff201c0042007d708c809;
    inBuf[10391] = 256'he9093509be07c205a403d901aa0006007bff79feb6fc74fa80f8d9f719f908fc;
    inBuf[10392] = 256'hadffc1024f0436043e038302c7021104ab058e0609062c049301f7febafcb7fa;
    inBuf[10393] = 256'h77f8bcf5ddf2c0f066f054f231f6e3fa12ffd4011d039d033c0484054307a708;
    inBuf[10394] = 256'hbc080407bb03c2ff32fcd8f9faf854f963faaffbfbfc32fe47ff2500a700a900;
    inBuf[10395] = 256'h250035fffdfda5fc64fb7efa48fa17fb08fdd1ffc0020205fd059d056a044403;
    inBuf[10396] = 256'hdb0252033204a604ea03ca01b8fe8afb1bf9f2f704f8d9f8def9acfa30fbb0fb;
    inBuf[10397] = 256'h8efc05fe06002e02ed03d904e1045004ac036d03ad031c044404c903ae025f01;
    inBuf[10398] = 256'h780061000e010502a0025d02250157ff93fd6cfc34fce7fc35fe9fffb0001c01;
    inBuf[10399] = 256'hd100ffff0dff68fe57fed6fe9eff480082004700e6ffc8ff3a0042019002a803;
    inBuf[10400] = 256'h34042704b6033703df029102fb01d7001cff21fd84fbd2fa2dfb4afc8bfd56fe;
    inBuf[10401] = 256'h79fe44fe46fefafe77004a02b5031e045c03c601150008ff02fff3ff7501fa02;
    inBuf[10402] = 256'h060464042e04a6031703be02a702a2027302f6012c014d00a8ff6fff86ff97ff;
    inBuf[10403] = 256'h3bff41fedafc89fbdffa25fb27fc4ffd04fef8fd58fdbcfccdfce3fde7ff7102;
    inBuf[10404] = 256'he704cc06e30720089a0787062d05d203b102e4015201cd003e00baff84ffe1ff;
    inBuf[10405] = 256'hd7000102bd027a020c01dbfebbfc77fb6dfb68fcc1fdbdfef8fe95fe15fe0cfe;
    inBuf[10406] = 256'he7feaa00f60241050207c4075807e305c6038b01c8ffddfec4fe25ff82ff78ff;
    inBuf[10407] = 256'h01ff7cfe6dfe31ffb10061028f03bd03df026801040028ffdffee3fed4fe7cfe;
    inBuf[10408] = 256'h03fec8fd13fee1feedffd100460145010501ba00830065006600990028012702;
    inBuf[10409] = 256'h6d0391041d05ca04b20355024b01fa00620121029e026502500187ff76fda0fb;
    inBuf[10410] = 256'h6bfa0ffa97fad2fb6dfd1affa200e901f002b80328041a047e036c022d011a00;
    inBuf[10411] = 256'h6eff2cff1fff11fff6fef4fe31ffa6ff0f00faff19ff86fdc5fb77fa01fa61fa;
    inBuf[10412] = 256'h29fbd2fb19fc26fc55fceefcf7fd28ff160089009f009f00c50026019c01e901;
    inBuf[10413] = 256'hef01bd016f0111018d00b9ff8afe37fd28fcc4fb31fc29fd1efe90fe58fec7fd;
    inBuf[10414] = 256'h7cfd05fe79ff71013803340438049103ca02500232022b02e10123010a00e7fe;
    inBuf[10415] = 256'h04fe7cfd4afd63fdccfd9cfedeff6801df02e703550447040704d703c603a903;
    inBuf[10416] = 256'h4b03a102d2010c015d00a0ff8efe03fd3afbacf9caf8baf842f9f3f989fa33fb;
    inBuf[10417] = 256'h6ffca7fecf013e0500085a093e09510876072a072d07ad06d2046d0140fdacf9;
    inBuf[10418] = 256'heaf760f865fa9dfcc6fd68fd02fcacfa5cfa53fb05fd7ffefdfe6afe55fd8efc;
    inBuf[10419] = 256'h99fc64fd59fec8fe62fe6cfd99fca2fcdafd1000b9023a053907ae08a7091a0a;
    inBuf[10420] = 256'hce097708f00576029bfe0afb3df85af63cf5b1f4b3f46df516f7aff9eafc4100;
    inBuf[10421] = 256'h2a035105b1067007a8075b077a06fd0410030e0152ff05fe22fd81fc05fcc2fb;
    inBuf[10422] = 256'hf8fbd7fc4dfefaff4f01d8017b0187007effbcfe44feb6fd9cfccafa9af8d2f6;
    inBuf[10423] = 256'h43f660f7eaf90dfddfffcb01ce0263031b041f0515065806640522030f00f6fc;
    inBuf[10424] = 256'h7dfae3f802f88ef764f7aff7daf840fbd6fe17032807210a5c0bbb0a9c089f05;
    inBuf[10425] = 256'h7402a0ff5bfda3fb64fa94f93ff988f981fa10fcf3fdd7ff71019f026c03f703;
    inBuf[10426] = 256'h4f046d04380492037c022901e9ff0affc6fe2fff140027011e02c10202031803;
    inBuf[10427] = 256'h5103d803a4046d05b50513057c034301f0fe0ffde6fb62fb3dfb50fbabfb8bfc;
    inBuf[10428] = 256'h2bfe86003a03ad055c071008e2071207d3052604ec0120ff06fc26f917f73cf6;
    inBuf[10429] = 256'h95f6c1f73df9a8faecfb33fdadfe69003302a50364044d048b038202a6014b01;
    inBuf[10430] = 256'h83012302cf022d03fe0235020401d5ff12fff5fe6afffeffffffeafec3fc27fa;
    inBuf[10431] = 256'h1cf89ff70cf9e1fbfefe3d010802ae0125016401c102af041406f105fe03e400;
    inBuf[10432] = 256'hdcfd0cfceafb13fd94fe79ff48ff33fee4fc1afc45fc6afd2eff0c019902a603;
    inBuf[10433] = 256'h390470046e043a04b203ae02230126ff02fd2dfb10fad6f961fa54fb39fcbffc;
    inBuf[10434] = 256'hf0fc22fdc9fd33ff5001a7038c056b061506cc041b0385014b0055ff5bfe2bfd;
    inBuf[10435] = 256'he5fbf3fad7fadefbeafd660084029603590302021f0057fe17fd6afc16fcccfb;
    inBuf[10436] = 256'h5dfbdffaa1fafafa08fc99fd42ff91003e0158013e015701dc01c502c5036e04;
    inBuf[10437] = 256'h7f0409045a03db02e4027b035004e804d104c903e6018eff40fd69fb49fae4f9;
    inBuf[10438] = 256'h08fa73faeffa5efbc6fb54fc4afdd9fe0e01b4034f06430812098e08f706e604;
    inBuf[10439] = 256'h0903d0013f01fc007d005fffacfdcafb47fa96f9d2f9b5facffbcefca8fd8efe;
    inBuf[10440] = 256'hbaff2f019b027303480316024c00a3fec1fddbfd8cfe21fffdfeeefd4efcddfa;
    inBuf[10441] = 256'h52faf8fa9cfcaffe8f00dc019202ec0227035b0366030b032302c40042ff11fe;
    inBuf[10442] = 256'h9efd16fe54ffee005f022f0321034b02fb0092ff60fe87fdf1fc76fc03fca7fb;
    inBuf[10443] = 256'h95fb09fc22fdbffe920038025e03e903fb03db03d3030d047e04eb0400057804;
    inBuf[10444] = 256'h45039601cfff60fe99fd7bfdc8fd23fe40fe14fed9fde3fd69fe5dff6b002401;
    inBuf[10445] = 256'h4101d0003500f6ff7200ad014a03af045405fc04cd033202a9008fff03ffeafe;
    inBuf[10446] = 256'h08ff24ff1cffe6fe8ffe2dfed4fd89fd45fdf6fc8afc04fc8efb71fbf9fb48fd;
    inBuf[10447] = 256'h3aff65013c0355049e045e040304e203ff0300046d030002dcff86fdb7fbfefa;
    inBuf[10448] = 256'h78fbcbfc5afe8fff1c001500d4ffbcff00008b0015014d010601540086fff4fe;
    inBuf[10449] = 256'hddfe42ffe4ff5f006100caffc1fea4fddbfca2fcf2fc83fd01fe3cfe51fea3fe;
    inBuf[10450] = 256'ha5ff9101370404073109180a7e099907e804fa0132ffb9fc98fad9f899f704f7;
    inBuf[10451] = 256'h35f71ef88cf942fb0dfddbfeb1008d024a04a70569066c06c505c104b103ca02;
    inBuf[10452] = 256'h12027301d3003400c5ffb7ff0d009000e100b300040038ffeafe8bff1401f702;
    inBuf[10453] = 256'h6004ac04ca034e021901cf0070015202900294018eff64fd38fcc4fcf7fef801;
    inBuf[10454] = 256'h9d040b061b064a055e04ef030f045d045f04d203d702e101650191013c02fa02;
    inBuf[10455] = 256'h560310033002f900cdff05ffd2fe2affd9ff8400d5009d00f7ff3dffe1fe36ff;
    inBuf[10456] = 256'h390083018002bd02260212012000d5ff50004501290287023f029301f000a100;
    inBuf[10457] = 256'ha200a600510079ff48fe2bfd94fcbffc9cfde8fe530099019c0243036b03ed02;
    inBuf[10458] = 256'hbf01020008fe42fc0afb7afa75fac4fa3dfbdefbc0fcf1fd53ffa0008801d901;
    inBuf[10459] = 256'h9c0109015e00bbff1aff64fe90fdc7fc54fc75fc36fd5dfe84ff4b008f007200;
    inBuf[10460] = 256'h3a0024002f001b008cff4efe70fc53fa85f88cf7b2f7fef836fbf3fdbc001603;
    inBuf[10461] = 256'h9c041105780411034a0188ff06feccfcbffbcdfa13fad5f94dfa7afb14fd9efe;
    inBuf[10462] = 256'haeff2e006d00e500ec0174030005de058b050104b90176ffedfd71fdd7fda0fe;
    inBuf[10463] = 256'h3fff5afff3fe5dfe00fe22fec8feb0ff7d00f1000e010e014501e301cd02aa03;
    inBuf[10464] = 256'h1104c603dd02b501c30056007900f6007e01dc010b0230027c020c03d1039404;
    inBuf[10465] = 256'h0605e4041104ab0208019effd6fedafe87ff7e005401d6011f0280023e035204;
    inBuf[10466] = 256'h5305a305cb04c8022400b2fd28fcc2fb31fcd6fc34fd3dfd5bfd1bfecdff3502;
    inBuf[10467] = 256'ha0044406b0060606e404fa03a903d703180405048c03f902b402f2028903fc03;
    inBuf[10468] = 256'hcb03c102080108ff2afdb4fbbbfa4cfa87fa91fb68fdc4ff1602c70380046004;
    inBuf[10469] = 256'hdf037f0378039d037e03c70291015c00caff36006a01b10235037a02a70070fe;
    inBuf[10470] = 256'hb8fc10fc75fc5efd18fe36fed1fd6dfda5fdbefe74001202d1024202860047fe;
    inBuf[10471] = 256'h5dfc75fbc4fb01fd94feefffc20015013b0190013d022003d703ee031f038701;
    inBuf[10472] = 256'h97ffe4fddafc89fca1fcaffc6cfceefb9cfbe1fbdffc44fe6effcaff33ff0dfe;
    inBuf[10473] = 256'h13fdeafcc2fd41ffb9009201a0013201db001201ef0126033004990431041103;
    inBuf[10474] = 256'h7e01c1ff0efe88fc4cfb79fa28fa5dfafafad1fbbafcacfdbefe07007f01e902;
    inBuf[10475] = 256'he703240485033902a00012ffbcfd91fc6ffb50fa6df925f9c5f94ffb63fd65ff;
    inBuf[10476] = 256'hc700540147011c014a01f701df027b034b031d022300dffde6fb9ffa2dfa74fa;
    inBuf[10477] = 256'h35fb35fc48fd50fe2fffc9ff0800f0ffa7ff6dff76ffd7ff760010015e013801;
    inBuf[10478] = 256'ha700d8ff0aff66fefafdb6fd83fd57fd3dfd51fdaffd62fe5bff720075013d02;
    inBuf[10479] = 256'hbd020103280345034e031b037e026301f1ff87fe9dfd8dfd63fed1ff57017802;
    inBuf[10480] = 256'hf402d7026002d1014801b300effff3fee7fd23fd00fda9fdfdfe9b000702e102;
    inBuf[10481] = 256'h0f03b7022302a20164016f01af01060250026e024602cd010a0122004dffbcfe;
    inBuf[10482] = 256'h84fe9afedbfe2cff91ff2a001401460278033c0431043e03ad01150017ff12ff;
    inBuf[10483] = 256'hf7ff570197023a0317035c026b019c001700c4ff65ffcdfe01fe43fdf3fc5bfd;
    inBuf[10484] = 256'h83fe2100b801d2023503f9026f02f501be01bf01c201900113016000aaff22ff;
    inBuf[10485] = 256'hdffee4fe2fffbeff9500a601c402a103e703600311023d0046fe80fc1bfb1bfa;
    inBuf[10486] = 256'h78f937f972f94efad1fbcafdd5ff77014f0240027401480025ff5bfe10fe44fe;
    inBuf[10487] = 256'hddfeb2ff97006301f2012b0204028101a60076fff1fd24fc37fa7cf85af72af7;
    inBuf[10488] = 256'h0cf8d0f9fbfbf8fd51ffdaffbbff49ffd9fe98fe7bfe5bfe13fea3fd2ffdeffc;
    inBuf[10489] = 256'h1afdcffd0cffb00080022b045605af050d0583035b0102ffddfc22fbd5f9e1f8;
    inBuf[10490] = 256'h40f80af877f8abf998fbe8fd1b00bd019702bc027202fe018001f6005400aaff;
    inBuf[10491] = 256'h2eff22ffacffb200df01cc022e03fc0261029601bb00c8ffaafe68fd3cfc81fb;
    inBuf[10492] = 256'h7efb32fc47fd37fe9bfe6ffe17fe2cfe1affdc00ef029d045705fe04e1037a02;
    inBuf[10493] = 256'h2101daff76feddfc4dfb60fac5fad7fc4f004e04b0078e099a092408e3058403;
    inBuf[10494] = 256'h680190ffcefd06fc60fa3af9fbf8d5f99bfbcdfdceff2501b001ae019801de01;
    inBuf[10495] = 256'haa02cd03d5044d05f904fc03c502d5018001bf0136026802f801dc0067ff1efe;
    inBuf[10496] = 256'h78fda1fd69fe58ffeeffe2ff4aff90fe3afea2fecaff5301af0268035503ab02;
    inBuf[10497] = 256'hd7013e010c01270149013e010501de001701d901f702f303310448033d018cfe;
    inBuf[10498] = 256'hf7fb2afa7bf9c9f9aafab2fbaffcb6fdfcfe95004e02b90362041404f7027c01;
    inBuf[10499] = 256'h24003dffd1feb4feb0feaffebefefcfe7dff37000801c40147027b025702d801;
    inBuf[10500] = 256'h0b010b0004ff1efe71fdf5fc8dfc25fcc6fb9ffbf3fbf2fc9afeaf00d202a504;
    inBuf[10501] = 256'he6057a065b068b05110403029cff3bfd53fb3afa0afa97fa85fb81fc63fd3afe;
    inBuf[10502] = 256'h30ff56008d018102da0267024001bdff4dfe48fdcffcd6fc39fddefdbdfed2ff;
    inBuf[10503] = 256'h0e0146023403930337032a02ae002eff1dfecdfd47fe4bff61000f0110016e00;
    inBuf[10504] = 256'h7cffa4fe25fef9fde0fd93fdfdfc56fc06fc69fc96fd50ff2201a00293030304;
    inBuf[10505] = 256'h1804ec0372038602100132ff4efde2fb53fbbbfbe4fc60fec2ffc9006c01c601;
    inBuf[10506] = 256'hf201f401c0014901a4000900bcffedff980081014f02bd02b0024502b0012201;
    inBuf[10507] = 256'ha8002e0090ffb6fea4fd7dfc74fbbcfa77fab4fa6efb92fc04fea5ff5301eb02;
    inBuf[10508] = 256'h4b045005e205fc05af051e056f04ba03fe02280228010700ecfe10fe9ffd9cfd;
    inBuf[10509] = 256'he1fd32fe65fe76fe8ffee4fe94ff89007d011a0223029001930080ffa6fe30fe;
    inBuf[10510] = 256'h20fe56feb0fe19ff91ff2200ca007101f30131022b020302ec01090251029102;
    inBuf[10511] = 256'h880211023e0153009eff4dff56ff80ff92ff76ff47ff38ff6fffdeff4f008100;
    inBuf[10512] = 256'h5900f1ff8bff61ff79ffa0ff82ffe8fee3fdcdfc1efc2efc05fd5afec3fff200;
    inBuf[10513] = 256'hdb01a902900394047805d6055f050e0435025000cbfed0fd44fdf1fcb6fc98fc;
    inBuf[10514] = 256'hb7fc23fdbdfd3cfe56fef0fd33fd7efc2dfc73fc45fd71fec1ff1d018102ee03;
    inBuf[10515] = 256'h48055706d906a506c80581042203ed01f50023004bff4efe2cfd03fcfbfa30fa;
    inBuf[10516] = 256'ha9f95ff957f9acf990fa27fc6efe1d01b603ae05a5069006c105b904f303a503;
    inBuf[10517] = 256'hb103bc0361036b02ec0034ffa8fd95fc15fc0efc4dfca2fcf8fc55fdccfd6afe;
    inBuf[10518] = 256'h29fff7ffba006301f1017102ef026f03e0032104090476036402f3006aff25fe;
    inBuf[10519] = 256'h75fd80fd36fe51ff74004d01aa018501f100110007fffcfd24fdb8fce9fcc4fd;
    inBuf[10520] = 256'h29ffd3006e02bc03a70436057a057b053405a304db03ff0233028201d4000000;
    inBuf[10521] = 256'hf4fecbfdcbfc3cfc35fc8bfcdffce5fc94fc3dfc5bfc4afd04ff1e01fc022704;
    inBuf[10522] = 256'h8504620431043f048c04c9049c04d50393022b01f5ff1dff91fe1ffea2fd1cfd;
    inBuf[10523] = 256'hbcfcbafc37fd22fe43ff4c00f7001b01ad00c4ff97fe77fdc2fcc5fc9afd15ff;
    inBuf[10524] = 256'hcc003802ef02d30213021b015000e9ffd3ffcbff89fff0fe20fe67fd12fd44fd;
    inBuf[10525] = 256'he4fda9fe41ff7fff6dff45ff49ff9dff2c00b300e6009f00faff4eff06ff69ff;
    inBuf[10526] = 256'h6f00ba01bd02f3021b02560013fee5fb47fa78f978f91ffa42fbc6fc9bfea900;
    inBuf[10527] = 256'hbc027b048905a805da046903cb017500a9ff61ff5bff3fffcefefdfdfcfc1bfc;
    inBuf[10528] = 256'h9ffba9fb23fcd8fc91fd33fec5fe6aff3a0030011b02b902d4025e0282018d00;
    inBuf[10529] = 256'hcdff6fff6fffa3ffd6ffe3ffc8ffa2ff9effdaff5600f4008301d201ca017301;
    inBuf[10530] = 256'hed006400fbffc2ffafffadffa2ff80ff4cff19ff02ff1cff6effe9ff7000e600;
    inBuf[10531] = 256'h40018a01e2015b02ef026e0397033b03610250016d0009003200a800fe00e000;
    inBuf[10532] = 256'h3c0052ff8dfe45fe92fe43ff01008300ae009c007b0070008200a200c000df00;
    inBuf[10533] = 256'h12016c01ef017e02ef021b03fd02aa024a02fa01bc017601050158007cff97fe;
    inBuf[10534] = 256'hd7fd55fd13fd03fd19fd59fdd7fd9ffea7ffc200b301440265023002dd019f01;
    inBuf[10535] = 256'h9201ab01c901c50187010c016a00bfff2dffcefeaefec7fe02ff3fff64ff68ff;
    inBuf[10536] = 256'h53ff37ff1fff05ffd2fe75fef2fd6efd25fd4bfdf0fdf7fe1e002101da014a02;
    inBuf[10537] = 256'h8c02bc02dc02d2027802b801a00061ff3afe5dfde4fccefc12fd9ffd65fe41ff;
    inBuf[10538] = 256'h010069005400c8fffafe39febefd97fd9ffda7fd9ffda5fdfbfdcffe12007101;
    inBuf[10539] = 256'h7802d6028402c301f70063000e00caff63ffcbfe25feb0fd97fdd6fd3cfe87fe;
    inBuf[10540] = 256'h8efe53fefcfdb6fd9cfdb5fdf9fd5efedffe75ff13009e0002013b015e018b01;
    inBuf[10541] = 256'hd4012d02620237028801610002ffbefddbfc75fc7dfcd0fc52fdfdfdd3fed0ff;
    inBuf[10542] = 256'hd600b30131023502cb011a015600a6ff1bffbbfe84fe76fe8ffebffef1fe10ff;
    inBuf[10543] = 256'h17ff1cff41ffa4ff47000a01bc01320257023002ce0143019900dcff24ff9bfe;
    inBuf[10544] = 256'h71fec1fe83ff7f006101dc01c90139017100cbff91ffd7ff790027018f018401;
    inBuf[10545] = 256'h14017700f1ffa0ff72ff34ffbefe1cfe93fd7efd11fe2dff59000201c600b7ff;
    inBuf[10546] = 256'h59fe68fd7bfdb7febc00dd0273042a051c05a8042e04d003630398023e016fff;
    inBuf[10547] = 256'h98fd4cfcf5fba5fc0dfea0ffd60062014701c5003000c9ffa7ffbaffd6ffd5ff;
    inBuf[10548] = 256'ha1ff4cff02ff00ff6fff4f0068016002e002c60233027b01f500cb00e400fd00;
    inBuf[10549] = 256'hd5005e00c4ff52ff42ff9aff2900ab00ed00e800b60079004000ffffa6ff33ff;
    inBuf[10550] = 256'hc0fe79fe83fee4fe84ff3700d7004d01900198015701c500eefffefe3cfee7fd;
    inBuf[10551] = 256'h13fe9bfe2dff82ff80ff53ff4affa3ff62004201e5010d02c1014601ee00df00;
    inBuf[10552] = 256'hfa00f2008800bdffdbfe4bfe51fee5feb0ff42004b00c5ffebfe0ffe6ffd1cfd;
    inBuf[10553] = 256'h09fd24fd6afde9fdabfea8ffc000c40190020f033a0311038f02b101860039ff;
    inBuf[10554] = 256'h07fe2efdcdfcdbfc34fdb4fd54fe2cff5600d0015b038904e70439049b027b00;
    inBuf[10555] = 256'h6bfedffc05fcc2fbd7fb11fc69fc01fd01fe6fff1c01ad02bd030d0498039602;
    inBuf[10556] = 256'h65015d00b2ff62ff41ff18ffc6fe57fe05fe14fea7fe9dff98002201ed000100;
    inBuf[10557] = 256'hc2fec0fd76fd05fe2dff70005c01c001c201b801e7015502bd02ba020502a700;
    inBuf[10558] = 256'hfefe91fdd0fcdbfc7dfd4dfeecfe35ff4dff80ff13000f013e024303c503a203;
    inBuf[10559] = 256'hf40207023301b3009500bc00f4000d01ec009300130084fff4fe63fec7fd1ffd;
    inBuf[10560] = 256'h78fcf6fbc7fb14fcecfc37febfff3f017d025c03e003250452047f04ad04c004;
    inBuf[10561] = 256'h8b04e203af020b0139ff9bfd88fc32fc89fc4afd19feacfee6fedcfebbfeacfe;
    inBuf[10562] = 256'hc0fee8fe06ff0bfffafef2fe18ff84ff36001101e8018f02ea02fb02e002bc02;
    inBuf[10563] = 256'hab02a8029102350271014e0002ffe3fd39fd1efd71fde3fd2afe26feeefdc6fd;
    inBuf[10564] = 256'hecfd77fe41ff00006f0072002500c7ff92ff99ffc4ffe4ffd7ffa4ff77ff82ff;
    inBuf[10565] = 256'he2ff8000220187018d013e01ce00710047004d006600730068004a002a001300;
    inBuf[10566] = 256'h0b00110027004e008100ad00b4007b00050076ff04ffd9fef5fe28ff33ffeffe;
    inBuf[10567] = 256'h76fe14fe1bfeacfe98ff7000c7007100a0ffc8fe61fe9dfe58ff3000c800fa00;
    inBuf[10568] = 256'hea00dc0009017201e7012202fa017301b200e6ff25ff72fec7fd2efdc7fcb7fc;
    inBuf[10569] = 256'h0efdb7fd84fe4afffaffad008301870291035904a0045a04bf032803da02ce02;
    inBuf[10570] = 256'hb5022302d800f1fee3fc40fb72fa86fa37fb1ffcf9fcb5fd6ffe47ff3a001f01;
    inBuf[10571] = 256'hc1010102e7019e0154012601150112010b01f100b7005100b8ff00ff57fe00fe;
    inBuf[10572] = 256'h2ffeeafef7fff5008a0194013601bf006d0046000f0079ff61fefffcdafb8ffb;
    inBuf[10573] = 256'h7bfc82fe1c018f034a051e06450625060706e80581057804a4022e0085fd29fb;
    inBuf[10574] = 256'h74f982f83bf870f800f9e2f91afba3fc6bfe4b001902a903cf0465054e058b04;
    inBuf[10575] = 256'h4203bd01530045ffa7fe5ffe42fe33fe34fe61fed1fe79ff2b00aa00ce009900;
    inBuf[10576] = 256'h3800e4ffc4ffd4fff3fffaffdeffb4ffaaffe5ff670006018501b10182011f01;
    inBuf[10577] = 256'hc800ae00d80021014c013001d0005f001a0026007100b700ab00210028ff0cfe;
    inBuf[10578] = 256'h30fde0fc32fdfefdf7fec9ff3b003c00eaff7aff22ff08ff2eff7cffc5ffe6ff;
    inBuf[10579] = 256'hd5ffa5ff7fff83ffbaff0b0047004a001400d2ffc8ff32001c014f0269030604;
    inBuf[10580] = 256'hf4034c036602a8014c0145014a010c01690089ffc6fe74feaafe31ffa2ffa6ff;
    inBuf[10581] = 256'h2dff71fed5fda4fde2fd51fe99fe85fe29fed7fdf4fdbafe1600ab01fd02ab03;
    inBuf[10582] = 256'h8f03ca02a901800086ffcefe48fedafd77fd26fd02fd2afdb1fd93feaaffbe00;
    inBuf[10583] = 256'h9101f601e2017001d90054000300e0ffcbff9dff51ff0bff0cff8dff9700f301;
    inBuf[10584] = 256'h3e0310043204af03cc02dd011c0195002c00b9ff24ff73fec5fd3dfdf6fcf2fc;
    inBuf[10585] = 256'h28fd84fdf3fd66fed3fe32ff7fffb8ffd8ffd9ffb7ff71ff13ffb7fe80fe90fe;
    inBuf[10586] = 256'hf1fe8dff3100a100af005c00d5ff5dff2eff54ffa8ffe9ffe6ffa0ff51ff49ff;
    inBuf[10587] = 256'hbeffaa00c601b7023d035803390321032e0347033003b502d201bd00caff3aff;
    inBuf[10588] = 256'h18ff31ff37ffe8fe33fe43fd62fcdafbd3fb47fc0bfdebfdbafe63ffe9ff5b00;
    inBuf[10589] = 256'hc9003a01ad0113025a026a023102a601d300d6ffdafe0afe82fd47fd4ffd8bfd;
    inBuf[10590] = 256'hf3fd81fe2effe0ff7000bc00b80080004a004c009a001d01a301000226022e02;
    inBuf[10591] = 256'h3f027402c5020e032b030b03bf0266021a02da018c010b0140002affe8fdaefc;
    inBuf[10592] = 256'hb2fb28fb2dfbbefbb7fcd8fddcfe8bffd6ffd4ffb6ffadffceff0f004c006500;
    inBuf[10593] = 256'h5200290012002800630098008b0018004dff6dfecffdb1fd17fec3fe5effa4ff;
    inBuf[10594] = 256'h90ff59ff54ffc1ffa700d601fd02d903490457042504d5037e032503c6025802;
    inBuf[10595] = 256'hd30133017c00c0ff1bffa6fe69fe56fe4bfe2bfeedfda8fd82fd9ffd06fe9bfe;
    inBuf[10596] = 256'h31ff99ffbeffa3ff65ff24fff9fee9fee7fed9fea5fe3efeb5fd36fdfefc3ffd;
    inBuf[10597] = 256'h04fe2bff68006701f001fd01b90162012d012601370136010a01bb0076007400;
    inBuf[10598] = 256'hdb00a10190025603af038603fb024f02c301750153013001e3006400cfff54ff;
    inBuf[10599] = 256'h19ff1cff3cff44ff0eff98fe02fe7efd38fd41fd88fdecfd49fe8cfebcfeeffe;
    inBuf[10600] = 256'h38ff99fffcff3b003900f0ff77fffcfea5fe84fe8bfe9bfe97fe76fe4bfe35fe;
    inBuf[10601] = 256'h55febdfe6cff4d00440134020303a9032a049804000560059c058705fa04ef03;
    inBuf[10602] = 256'h92023101150061fffdfea8fe25fe66fd9cfc21fc43fc17fd66fec6ffce004501;
    inBuf[10603] = 256'h3501d70071002f000f00f0ffabff2bff74fea6fde5fc54fc0bfc13fc67fcf0fc;
    inBuf[10604] = 256'h89fd10fe6ffeaffef1fe5cff0600df00b8015c02ab02b002930283028c029702;
    inBuf[10605] = 256'h74020402510195001e002300a60071013202a402ae026702ff019f0155011301;
    inBuf[10606] = 256'hbf005000d5ff74ff55ff88fff9ff7100af008000d8ffd7febafdc7fc2cfceffb;
    inBuf[10607] = 256'hf3fb04fcf8fbc4fb84fb6ffbbefb8bfcc4fd30ff880093013a028e02b102c202;
    inBuf[10608] = 256'hcb02bc027702e9011b0133006dff05ff20ffb7ff96006801db01bf0127016200;
    inBuf[10609] = 256'hd8ffdbff780072015e02de02d1026002e101a001b80101023002060271019700;
    inBuf[10610] = 256'hbcff1cffcdfeb2fe95fe3bfe8cfd99fc9cfbe1faa8fa0bfbedfb05fdf7fd7dfe;
    inBuf[10611] = 256'h82fe2bfec3fd98fdd3fd6dfe34ffefff7a00dc003b01bf0176024103e3031e04;
    inBuf[10612] = 256'hd90330036602c10167014d0146012401d9007f0046004e009400ef002e013601;
    inBuf[10613] = 256'h1301ed00f00029018801e40118020e02c60148019f00d5fff6fe19fe57fdc6fc;
    inBuf[10614] = 256'h6dfc3efc22fc09fceefbe1fbf7fb40fcbbfc57fdf8fd8cfe0dff85ff08009c00;
    inBuf[10615] = 256'h3701b701f601dc017701f900a400a60006019b0126026f0268022c02ed01d501;
    inBuf[10616] = 256'hf30132026c027d025402f6017c010801bd00b100ec005a01d60133024a020f02;
    inBuf[10617] = 256'h8d01e100240061ff91fea7fda3fc9afbbafa35fa32fabafab5fbeffc2efe42ff;
    inBuf[10618] = 256'h12009e00f30020012c011601db0081001700b0ff58ff14ffddfeb0fe91fe88fe;
    inBuf[10619] = 256'h9ffed4fe23ff84ffffffa300790176026c03210465043304ba0342030e033303;
    inBuf[10620] = 256'h9503f4031404d2033403540253014b004dff64fea0fd0ffdb6fc8dfc7bfc68fc;
    inBuf[10621] = 256'h46fc1afcfcfb06fc4dfccdfc71fd19feacfe20ff7bffccff15004c005a003100;
    inBuf[10622] = 256'hdcff82ff56ff7cfff1ff8700f9001301c9003f00b6ff69ff70ffbcff23007d00;
    inBuf[10623] = 256'hb600d300ee0020017801f1017602ec0239034e032c03e502930254023a024702;
    inBuf[10624] = 256'h68027b025c02ef013201360020ff12fe22fd55fca1fb03fb86fa49fa6dfa02fb;
    inBuf[10625] = 256'hf6fb17fd2bfe06ffa3ff1d0098002501ab01f701d0011e01f8ffa2fe72fdaffc;
    inBuf[10626] = 256'h81fce5fcbcfddcfe1d005e01850279031e0462044004cd033103a00247023902;
    inBuf[10627] = 256'h6502a702ce02bd026f02fa017c010f01bb0074002600c5ff4fffcefe51fee3fd;
    inBuf[10628] = 256'h87fd3efd08fde8fce7fc0afd4efda7fd00fe44fe65fe64fe4efe3dfe49fe88fe;
    inBuf[10629] = 256'hfcfe98ff3900b300db009e000b0051ffb7fe7afeb5fe59ff31000201a1010502;
    inBuf[10630] = 256'h400269029002b102bd02ac0282024f022002f601c5017b011901ae005c003e00;
    inBuf[10631] = 256'h5a009a00d400df00a40029008affe9fe64fe06fecffdb8fdbbfdd8fd0efe5afe;
    inBuf[10632] = 256'hadfeeefe06ffe8fea0fe50fe27fe4afec4fe77ff2900990096001a004dff76fe;
    inBuf[10633] = 256'he2fdc2fd1afebffe6dffe7ff12000200ecff05006b000f01c6016102cb020e03;
    inBuf[10634] = 256'h4c039e03ff0349044a04de030a03fa01ec0012007eff1fffd2fe79fe0ffea6fd;
    inBuf[10635] = 256'h5dfd4cfd7cfde1fd69fe03ffa1ff3b00bf0012011701bc000d002fff5dfeccfd;
    inBuf[10636] = 256'h94fda7fddffd0ffe20fe16fe09fe15fe44fe8cfedcfe29ff78ffdfff72003301;
    inBuf[10637] = 256'h0902cc025003800361031103b7026d023a020e02d4017f010f0192001b00b9ff;
    inBuf[10638] = 256'h73ff4cff47ff6dffc0ff3a00be002401460111019300f5ff6aff13fff8fe0aff;
    inBuf[10639] = 256'h2eff54ff7affa3ffcffff1fff4ffc4ff5cffccfe2afe90fd09fd99fc3ffcfefb;
    inBuf[10640] = 256'he7fb0cfc7dfc3dfd42fe73ffb000d201bc0257039c03940357030403b6028102;
    inBuf[10641] = 256'h670263026802670256022e02ef019b013901d20070001c00dbffaeff8eff6dff;
    inBuf[10642] = 256'h3dfff1fe8cfe22fed9fdd5fd29fec5fe7aff0e00550047000400bcff96ff95ff;
    inBuf[10643] = 256'ha0ff8fff48ffcffe41fec1fd63fd2cfd13fd12fd2efd73fdeafd8efe4cff1200;
    inBuf[10644] = 256'hd0007f011b029c02f6022103270324033603660397038d030c030102960030ff;
    inBuf[10645] = 256'h3cfe00fe74fe46ff040056002600a3ff20ffe5fe0cff78fff2ff44005b004200;
    inBuf[10646] = 256'h1600f0ffd4ffb3ff7dff2bffc7fe6cfe36fe37fe72fedafe52ffb8ffe9ffd3ff;
    inBuf[10647] = 256'h78fff9fe8cfe66fea7fe45ff0d00b9000e01fb0098002100d0ffc7ff05006a00;
    inBuf[10648] = 256'hcf001a01440159016a0180019a01ac01a9018d0158011301c4006d000d00a4ff;
    inBuf[10649] = 256'h3dffeffed7fe0eff97ff5d003001de01420256022c02df017a01f500390037ff;
    inBuf[10650] = 256'h03fed1fce9fb7dfb97fb0bfc91fceafcfefce4fcd5fc04fd8dfd63fe62ff6100;
    inBuf[10651] = 256'h4301fd0193020e037803d6032c0471048e046104cd03cb027a011d0002ff5afe;
    inBuf[10652] = 256'h1efe19fe0efedafd92fd7dfde3fde6fe5c00e20104037b034803ad0201028101;
    inBuf[10653] = 256'h3301f1008c00eeff2eff7bfe06fee1fdf7fd1afe1afedbfd62fdd4fc68fc54fc;
    inBuf[10654] = 256'hbcfc9dfdd2fe1c003e010f028702b802b50284021b026e018a009cffe2fe8ffe;
    inBuf[10655] = 256'habfe0aff66ff88ff69ff38ff40ffbaffad00e5010c03d1030b04c40326036602;
    inBuf[10656] = 256'ha801f30041008cffe0fe5efe2efe68fe06ffd9ff9f001a012901d2003a0092ff;
    inBuf[10657] = 256'h04ffa4fe6efe4ffe2efef4fd94fd13fd90fc3ffc57fcfbfc21fe8cffe100ce01;
    inBuf[10658] = 256'h2f021c02d801ac01bc01fb0137023e020202a4015b0157019601e301ed017201;
    inBuf[10659] = 256'h6a000effc4fdeefcc0fc2efd00fef1fed7ffa90070013102d70239033803d102;
    inBuf[10660] = 256'h21026001b400240097fff4fe3dfe97fd2ffd1cfd4dfd8efdaffda3fd8afd93fd;
    inBuf[10661] = 256'he2fd6dfe07ff7effbcffd3fff7ff5200f200bd018202120356034d0303038902;
    inBuf[10662] = 256'hec0137017400b1fff9fe57fed6fd8cfd8bfde0fd7bfe2fffc0ff0400fbffdaff;
    inBuf[10663] = 256'hedff66003a011d02ab02a1020802350198007e00e5008501fb01ff018901c900;
    inBuf[10664] = 256'h070071ff0affb2fe3dfe98fdd2fc17fc9ffb95fb0bfceefc0efe27fff6ff4e00;
    inBuf[10665] = 256'h2b00bdff53ff3effacff8a008d015702ae0298025f025f02cf0294034a047d04;
    inBuf[10666] = 256'he903a9022601ddff16ffbefe80fe03fe2dfd3efcaafbd7fbe0fc7ffe35008a01;
    inBuf[10667] = 256'h41026c024d0227021202f801a601f300e5ffaefea2fd09fd05fd81fd3bfee2fe;
    inBuf[10668] = 256'h3bff40ff11ffe4feeefe49ffedffaf005a01c201d601a1014201de008d005400;
    inBuf[10669] = 256'h29000000d5ffbbffcbff13008a00060150013c01ca00250095ff52ff69ffacff;
    inBuf[10670] = 256'hd6ffb1ff3fffbbfe78feaafe4eff2800ed007301c50114028d022f03c303f503;
    inBuf[10671] = 256'h85036d02e40045ffe2fde4fc44fce3fba8fb9bfbdafb81fc89fdbafec0ff5b00;
    inBuf[10672] = 256'h7e005600270019001c000000acff45ff27ff9fff9c009c01f0013801c5ff8bfe;
    inBuf[10673] = 256'h9dfe79009d03b10643088f07eb048b01cefe83fd9dfd6afe23ff5cff2ffffcfe;
    inBuf[10674] = 256'h13ff77ffe3fff7ff7dff8afe7ffde9fc46fdc2fe060137033b043503070093fb;
    inBuf[10675] = 256'h7bf777f58df684faf3ffda0483073a078004b80072fdbefbe3fb74fdcaff6a02;
    inBuf[10676] = 256'h3e052e08bd0a0e0c0d0b1207860019f951f375f166f406fb8d02ca079a08e104;
    inBuf[10677] = 256'h86fe73f82df5cdf5bef94eff9c045808070ac909fb07ed04ee0083fc90f84af6;
    inBuf[10678] = 256'hcff69cfa15017008260ed40f340ccc03eef8f8ee26e961e99deff4f96005c00e;
    inBuf[10679] = 256'hba134013b10dab04a6fa5bf219ee16ef07f52bfedc07700f0213f611ee0c6f05;
    inBuf[10680] = 256'h5ffd8df660f29bf13bf470f9ccff94053e09d809460741022dfcd1f6e7f3aaf4;
    inBuf[10681] = 256'h57f9e5002e09930f0012c80ff009b40271fc9ff858f7a4f75df8f4f8adf92efb;
    inBuf[10682] = 256'hbefdc100e802f602a100f9fcfef989f939fcf900830597074206670249fe40fc;
    inBuf[10683] = 256'h6efd20014705b8076c0705054b02fc00ad0179039c049a03300085fb7af79df5;
    inBuf[10684] = 256'h62f6daf873fbdefcb4fc8ffb9bfaeffa01fd7d007904de07e309510a8a094408;
    inBuf[10685] = 256'h1e074a0677051204b60187fe3efbd3f8f5f7acf856fa0cfc1bfd61fd41fd53fd;
    inBuf[10686] = 256'hfafd32ff9f00cb016902700205025c019400bbffdcfe12fe8bfd7afdfdfd06ff;
    inBuf[10687] = 256'h5d00b201b9024a0363032303ac0216026801a300dcff38ffe0fee2fe27ff77ff;
    inBuf[10688] = 256'ha1ffa3ffaeff130004016902d903c704c104ad03ce01aaffc2fd64fc97fb32fb;
    inBuf[10689] = 256'h00fbe9fafffa6dfb55fcaffd37ff790004019d0075ff21fe67fde2fdadff4702;
    inBuf[10690] = 256'hc8044a065306100533038f01b500b5003301a901bd016201cf004f000f000300;
    inBuf[10691] = 256'hf0ff8bffa2fe3cfda6fb69fa17fa0ffb40fd11009902f803c2033502140044fe;
    inBuf[10692] = 256'h52fd60fd42fe89ffd500ed01bd0234033503a6028c012000c6fee2fdaefd25fe;
    inBuf[10693] = 256'h0bff14000501c00133024b02ee010f01caff6ffe6dfd23fdadfdcdfe0300cb00;
    inBuf[10694] = 256'hdf004c006cffa7fe42fe44fe85fedafe31ff96ff1800a80016012a01cf003600;
    inBuf[10695] = 256'hc7fff0ffe5007a0234047d05ec05670523047502a600e0fe2ffda1fb56fa85f9;
    inBuf[10696] = 256'h61f9fff948fbfcfcc7fe5f0095015c02c102e302da02b3026702e40121012800;
    inBuf[10697] = 256'h1fff41fec2fdbefd2dfee3fea8ff4d00b700e200de00ca00cb0003017f012802;
    inBuf[10698] = 256'hbb02dd024202d600dcfedcfc73fb0efbc0fb3efd04ff9800b2014f029302a102;
    inBuf[10699] = 256'h7e0210023501f0ff7cfe44fdbcfc27fd6dfe1d0092013d02e701cc007aff94fe;
    inBuf[10700] = 256'h85fe55ffb1001a0224039b0386030c03510261013b00dffe6afd17fc2bfbd7fa;
    inBuf[10701] = 256'h25fbeffbf4fcf8fddafea0ff5f002601e0015d026f020b026601db00be002501;
    inBuf[10702] = 256'hd1014a022a0256011d0013ffbbfe49ff7d00d001b402da0247024301270034ff;
    inBuf[10703] = 256'h83fe09feaffd64fd27fd09fd26fd9efd78fe9affba007a018e01ec00dfffecfe;
    inBuf[10704] = 256'h8ffefafef4fff20067010e011300fafe57fe7dfe5bff8b00900118022202ee01;
    inBuf[10705] = 256'hcc01ee014a02a302b30252028c019d00d2ff67ff6bffb7fffdffedff50ff29fe;
    inBuf[10706] = 256'hb7fc64fb99fa98fa5ffbadfc20fe65ff5c001601c00177023003ba03d9037203;
    inBuf[10707] = 256'h9b029901c1004c0044008600d400f800d7007500ebff57ffcbfe53fef9fdcdfd;
    inBuf[10708] = 256'he7fd5cfe2aff2e002501c501dc016a01a000caff20ffb7fe7afe49fe1efe14fe;
    inBuf[10709] = 256'h58fefefeeaffd00059015901e7005400fcff13008c002901a201cb01a8015a01;
    inBuf[10710] = 256'hff009e0028008cffd2fe24fec4fde9fda4fed1ff1f013902df02fd02a302f401;
    inBuf[10711] = 256'h0b01f4ffb5fe61fd2afc52fb16fb89fb8efce1fd3cff6d0068012e02be020403;
    inBuf[10712] = 256'hec027802d0013a01f3000c015c0196017701f30036008bff29ff18ff2fff33ff;
    inBuf[10713] = 256'h01ffa2fe40fe0cfe20fe72fee3fe4dff96ffb5ffacff81ff41ff00ffddfef5fe;
    inBuf[10714] = 256'h57fff7ffb2005d01de0136027a02bd02fa020a03c0020202e700b7ffcdfe66fe;
    inBuf[10715] = 256'h89fefefe74ffa9ff89ff2fffccfe89fe77fe93fedcfe58ff0e00ee00c5014502;
    inBuf[10716] = 256'h2a025c0108008dfe51fd91fc55fc7afce0fc7ffd6bfeb0ff3701b602d0034004;
    inBuf[10717] = 256'h030457039a021802e601e501df01ab013e01a500f3ff34ff71fec0fd48fd35fd;
    inBuf[10718] = 256'h99fd54fe1aff91ff80fff2fe2dfe95fd77fde6fdbffebcffa0004d01c3011602;
    inBuf[10719] = 256'h57028502940275022202a6011d01a40052002f002c002f001c00e4ff8fff39ff;
    inBuf[10720] = 256'h08ff19ff6cffdeff34003200b4ffcafeb3fdcffc70fcbcfc99fdbefed6ffab00;
    inBuf[10721] = 256'h36019301df0118021b02bf01ff000d0047ff02ff5aff1b00de003e0113018300;
    inBuf[10722] = 256'he6ff96ffbaff3a00d6004d0182017b01580134011b010401e200af006d002700;
    inBuf[10723] = 256'he2ff9aff43ffd5fe50fec0fd42fdf0fce3fc21fda3fd53fe15ffc9ff53009b00;
    inBuf[10724] = 256'h97004f00dcff66ff1cff20ff7dff29000301e501af0248039f03b0037f031a03;
    inBuf[10725] = 256'h9b021a02a5013501b6000c002aff18fef3fce2fb09fb85fa6ffadcfadcfb68fd;
    inBuf[10726] = 256'h56ff5a01100325047404180458038d02f5019e01630112018200b7ffdefe36fe;
    inBuf[10727] = 256'heffd14fe81fe01ff66ffaaffe6ff4100c4004c018f0145015000d9fe48fd13fc;
    inBuf[10728] = 256'h92fbdafbc5fc05fe51ff7900660111027c02ab02a8028902630245022902ff01;
    inBuf[10729] = 256'hb2013f01b1001d008fff06ff7dfef4fd88fd63fdadfd74fea0fff60032021e03;
    inBuf[10730] = 256'h970394031b033f022101f2ffe6fe1cfe98fd3ffde9fc88fc35fc29fc95fc7dfd;
    inBuf[10731] = 256'hacfec4ff7800b000950077009600fe008401e501f101a9013a01e600de002f01;
    inBuf[10732] = 256'hc5017202040352033f03c202ee01e700defffafe4afeb8fd20fd68fc99fbe7fa;
    inBuf[10733] = 256'ha2fa0bfb36fcf7fdecffa701dc0276039703810367035a0347030f03a2021302;
    inBuf[10734] = 256'h88011f01d5008600020031ff30fe40fda5fc81fcc3fc35fda4fdfefd58fed1fe;
    inBuf[10735] = 256'h76ff2b00bb00fb00e30090003400f6ffddffd7ffd2ffc7ffc2ffd7ff0c005700;
    inBuf[10736] = 256'ha900f6003e018a01d7010f021002c2012a017200dbff97ffb2ff0c0068008b00;
    inBuf[10737] = 256'h64001300cfffd2ff2e00c300510194016701d300090043ffa3fe2bfec2fd47fd;
    inBuf[10738] = 256'hb2fc18fca5fb89fbddfb9efca3fdbdfebcff7f00010154019301da013e02bb02;
    inBuf[10739] = 256'h4003b8030c0432042b04f5038903d802d701880007ff8dfd5efcb5fbaefb3afc;
    inBuf[10740] = 256'h22fd1bfee1fe4eff69ff5eff63ff9cff0b008d00f2002201270123013e018201;
    inBuf[10741] = 256'hcf01f701d5016c01e5007a00480042003700f6ff6fffc2fe2dfee3fdf3fd3dfe;
    inBuf[10742] = 256'h87fea1fe80fe41fe19fe3bfec1fe9dffa6009d013e025802db01e300bbffc0fe;
    inBuf[10743] = 256'h40fe56fee7fea7ff4800a000ba00c100e3002e018401bb01c401b301ba010002;
    inBuf[10744] = 256'h7702d702c9021802df0085ff8cfe40fe97fe3cffc3ffecffc2ff7aff41ff15ff;
    inBuf[10745] = 256'hc6fe26fe3ffd69fc15fc8dfcb8fd13fffeff110058ff4cfe92fd9dfd78fed6ff;
    inBuf[10746] = 256'h4401670222038803b403b003770301035d02b4013501f600e800e100ab002a00;
    inBuf[10747] = 256'h66ff83feb4fd2ffd1afd7dfd4afe55ff59001d0186019d018e018c01ab01d201;
    inBuf[10748] = 256'hd2017c01c400d6fff5fe5dfe20fe26fe35fe23feecfdb2fdabfd01feb6fe9dff;
    inBuf[10749] = 256'h780013015a01630160017701b401ff012602fc017801ab00c2ffe8fe3bfec3fd;
    inBuf[10750] = 256'h83fd85fdcffd5efe1effdcff6600a400a00085008400b6000701500171016501;
    inBuf[10751] = 256'h4a014c018001d0010d0200028b01c800f3ff54ff23ff6aff00009e000001fa00;
    inBuf[10752] = 256'h9000f2ff5bfff0feb5fe86fe3afec7fd54fd1efd5bfd0cfeeafe92ffb8ff55ff;
    inBuf[10753] = 256'hb0fe3bfe4ffef8fef7ffe300630161010d01b4009600c80028017c019a017b01;
    inBuf[10754] = 256'h3401ef00cb00cb00dd00eb00e300c100940067003b000e00d8ff97ff5dff4bff;
    inBuf[10755] = 256'h78ffefff9d004b01bc01c6016001a700d3ff15ff83fe1efed8fdabfda3fdd4fd;
    inBuf[10756] = 256'h39feadfef7fee8fe85fe19fe0efeb2fe0400a7010303a1035f037a0261017200;
    inBuf[10757] = 256'hc6ff3bffa5fe00fe79fd5afdcdfdaffea9ff5b00930069002c002b0084002001;
    inBuf[10758] = 256'hc3013202570241020b02d601b301a3019b018f01640101015b007fff99feeffd;
    inBuf[10759] = 256'hc0fd1ffef4fef9ffd80051014e01dd00210049ff77fec3fd3ffdf6fce2fcfcfc;
    inBuf[10760] = 256'h39fd8ffd00fe96fe4cff06009900d700ac003900c5ff98ffd6ff6d0016018701;
    inBuf[10761] = 256'ha50188016e019201fa016d029d0255029b01bd002d0041000d01510290033904;
    inBuf[10762] = 256'hed0390025d00d6fd95fb1bfab0f953fabefb87fd46ff9d004f0148019f0094ff;
    inBuf[10763] = 256'h93fe0ffe4efe49ffa300c8013c02dd01e700dcff39ff35ffadff5800f7007901;
    inBuf[10764] = 256'h0002a7025503bd0385038402e7002fffe7fd57fd66fda8fd9dfd05fd04fc05fb;
    inBuf[10765] = 256'h87fae0fa0ffcd3fdd0ffb2013c035404e704ea0469049203ab020102c801f401;
    inBuf[10766] = 256'h430261021002410128001cff71fe66fe16ff6a001e02c703d704cc046c03e400;
    inBuf[10767] = 256'hc9fdeffa0cf95ff8adf865f9f1f90ffaf1f900fa99fad4fb74fd13ff74009e01;
    inBuf[10768] = 256'hc8022904b8051607c1076207fd0505042302e3006f009500ec001401ee009d00;
    inBuf[10769] = 256'h5500380048006a0084009b00be00e600ef009c00b5ff45fea0fc42fb99fad3fa;
    inBuf[10770] = 256'hc0fbf4fc03fea8fed5feb6fe87fe7ffec8fe7fff9e00fe0159034b048a040904;
    inBuf[10771] = 256'h0103d701f30080005e004600fdff77ffddfe6cfe37fe22fefbfda4fd3afd12fd;
    inBuf[10772] = 256'h83fd9dfe1d008701620284022402a001440121010101a500ffff43ffbcfea4fe;
    inBuf[10773] = 256'hf2fe60ffa1ff9fff80ff90ff1200090134023c03db03f403a20319038002f201;
    inBuf[10774] = 256'h7501f80062009effa2fe7dfd65fc96fb33fb35fb66fb7efb5ffb27fb1dfb80fb;
    inBuf[10775] = 256'h60fc85fd9dfe7fff3f001b014b02c30329050c063106b105ee04580419040104;
    inBuf[10776] = 256'hb803f502b90154002fff86fe54fe62fe6efe59fe38fe2afe3ffe6efe96fe9efe;
    inBuf[10777] = 256'h8cfe82fe99fedbfe36ff87ffb3ffb8ff9fff70ff34fff5fec6fed2fe4aff3700;
    inBuf[10778] = 256'h7301a80270038c030e03410284011801fb00f000b7002d005bff6afe86fdc0fc;
    inBuf[10779] = 256'h13fc83fb25fb1efb99fba6fc25fedaff8201db02c4033a044a041104ba035f03;
    inBuf[10780] = 256'h04039502ef01f200b2ff75fe97fd67fdfbfd14ff450028018a01790141012d01;
    inBuf[10781] = 256'h6201d5014f028c025d02bc01bf0091ff64fe57fd73fcbefb3bfbedfae2fa23fb;
    inBuf[10782] = 256'h9ffb33fcb8fc0dfd35fd63fdd5fdbbfe2400ec01c9037105a80643072d076a06;
    inBuf[10783] = 256'h100554038e011c003fff0fff65ffefff5f0086005e000400a9ff6dff64ff91ff;
    inBuf[10784] = 256'he5ff3f0075005600bbffaafe55fd0efc33fb03fb7ffb79fcacfdd8fedcffb900;
    inBuf[10785] = 256'h770112028102b502a8026b021d02d10183012801ad00180093ff4dff61ffc4ff;
    inBuf[10786] = 256'h44009c00a3006000f9ff9dff6eff6bff7fff98ffaaffa8ff84ff26ff7afe8ffd;
    inBuf[10787] = 256'ha7fc16fc24fce4fc1ffe74ff96006401f4017b021c03c5034e048f0476041d04;
    inBuf[10788] = 256'hb0033e03be02190243014b0060ffb0fe4dfe2bfe2efe3ffe56fe7bfeadfed0fe;
    inBuf[10789] = 256'hc3fe71fee2fd49fde5fcd6fc10fd5bfd6dfd14fd5bfc89fb08fb44fb77fc8afe;
    inBuf[10790] = 256'h17018803500528062b06c0055e054f058405a905660598046c0344026e01f100;
    inBuf[10791] = 256'h9800120036ff28fe42fdd3fcf5fc71fde3fdfefdbbfd4ffd0cfd2ffdbafd74fe;
    inBuf[10792] = 256'h12ff5aff31ffa8fef5fd53fdf9fc15fdb5fdbffe01003a012402a102c002b002;
    inBuf[10793] = 256'had02ea02750337040805bc0526061d067f0531042d029effe4fc7bfad8f833f8;
    inBuf[10794] = 256'h70f835f918fad1fa5efbf2fbc4fcecfd54ffc8001a024303490420059f058705;
    inBuf[10795] = 256'hb00433037701fcff25ff0fff80ff12008700d00005015801e901930220036803;
    inBuf[10796] = 256'h36037a025201dbff41fec5fc8cfba1fa08fab9f9acf9f2f99efaabfbe8fc0cfe;
    inBuf[10797] = 256'hd9fe48ff88ffeeffb700e10127032a04a8049e043b04b7033b03ca025a02f201;
    inBuf[10798] = 256'ha30180018901a201a0016c010d01a700680065008e00bb00bf007a00e1fff7fe;
    inBuf[10799] = 256'hcefd88fc5afb86fa3efa8cfa43fb13fcb9fc22fd85fd43fe9bff79016b03d004;
    inBuf[10800] = 256'h2e0578042203da0131014f01ed018802b2025502b3012401e200e100de009900;
    inBuf[10801] = 256'hf6ff10ff2cfe81fd24fd0bfd11fd14fd06fdeffce0fcf5fc4cfd06fe28ff8f00;
    inBuf[10802] = 256'h0502450303041f04b60302035402ed01d901f3010202d1015201a9001400d0ff;
    inBuf[10803] = 256'hefff48008a007000efff39ff9efe60fe84fed0fef3feb3fe1bfe6dfdfbfcf5fc;
    inBuf[10804] = 256'h4cfdb9fdfbfdeefd9bfd3afd0afd38fde7fd22ffce00b90295040a06dd060507;
    inBuf[10805] = 256'ha006ea05180538043603f5017700eafe95fdb8fc5ffc6bfcbffc43fde8fdb3fe;
    inBuf[10806] = 256'h97ff71001d017501680111018800d4fff5fedafd85fc36fb45fa00fa8efad2fb;
    inBuf[10807] = 256'h76fd21ff9c00e9012d038204df051107ce07f0077d0797066b0510047e02a800;
    inBuf[10808] = 256'h94fe75fc9afa4df9aef8aff820f9d3f9abfa9efbb3fcf1fd4dffa900ef010e03;
    inBuf[10809] = 256'heb0365046504e103eb02b8017c0062ff8ffe12fefafd6bfe6fffd30046026003;
    inBuf[10810] = 256'hcd03a0033503e202d402fe0208039102820114009ffe67fd88fce2fb42fb9efa;
    inBuf[10811] = 256'h1dfafdf961fa37fb4efc5ffd2bfeb3fe23ff94ff2200e800ce01b0027f032104;
    inBuf[10812] = 256'h6c045204dd0325034a027601c10019007eff08ffcbfee9fe84ff770071013302;
    inBuf[10813] = 256'h900282023d02ef01a2014401a900bbff9cfe93fde7fcaefcbdfcc8fc72fc91fb;
    inBuf[10814] = 256'h56fa23f96df8a4f8e5f9f0fb60feb6008c02c5037604cd0408053d057105ab05;
    inBuf[10815] = 256'he305140638062b06b905b004fc02c20066fe5dfc0dfba0faedfa9dfb49fc9bfc;
    inBuf[10816] = 256'h7dfc1bfcb4fb86fbbcfb4dfc0ffdd5fd72fecffe01ff1fff42ff93ff2300ec00;
    inBuf[10817] = 256'he201dd02a403220455044d0442045c049804db04ed04a80415045703a2021202;
    inBuf[10818] = 256'h8001a90058ff78fd43fb2ef99ff7d8f6d2f63ff7d1f755f8d1f894f9edfaf9fc;
    inBuf[10819] = 256'h95ff5202ab044806fd06d60625062c051104fe0208022f017f000300b6ff90ff;
    inBuf[10820] = 256'h9cfff0ff8b006b018d02ad037404c2048104a80372022601e1ffbdfed2fd13fd;
    inBuf[10821] = 256'h68fccdfb3afb9afadef915f961f8ebf7e8f785f8c4f97afb72fd7dff6601f902;
    inBuf[10822] = 256'h2804fa046e05a805ed0569062307f00769082708090733050b0303016dff5efe;
    inBuf[10823] = 256'hb6fd3efdd8fc86fc51fc3dfc3bfc2efc00fca8fb42fb04fb19fb81fb14fca4fc;
    inBuf[10824] = 256'h09fd35fd4afd7dfdf9fde3fe3e00d70183030d052f06c606db068606fb057805;
    inBuf[10825] = 256'h1f05ee04d0049f042f045a0318027a0094fe9ffce5fa8af9abf848f830f848f8;
    inBuf[10826] = 256'h95f805f999f952fa08fbb6fb7bfc66fd93fe300027022704d505de061f07be06;
    inBuf[10827] = 256'h01061d05300457039702e8015a01f600a7007500660060006800850087004400;
    inBuf[10828] = 256'ha5ff98fe49fd22fc7efb85fb2afc16fdd6fd18fec1fde8fcd1fbdafa49fa45fa;
    inBuf[10829] = 256'hdcfa05fc9efd77ff4a01d7020904f504b9056606f2063707ff06360600059103;
    inBuf[10830] = 256'h1b02c70080ff12fe7cfcf0fac0f944f998f990fadbfb07fdcafd36fe85feedfe;
    inBuf[10831] = 256'h9eff80003c018b014d01880080ff92fef8fdc1fddbfd2cfea4fe49ff1e000c01;
    inBuf[10832] = 256'hf401b2021e033a033b0346036b03b60303040d04ae03d8028701d9ff09fe46fc;
    inBuf[10833] = 256'hb5fa73f985f8e0f78ff79bf703f8caf8e6f937fbaafc40fefefff7012b046006;
    inBuf[10834] = 256'h370852096c098008c4069a0464026a00dcfec1fd0dfdcdfc0afdb8fdc9fe0300;
    inBuf[10835] = 256'h00018d01aa016301f0008a003200c0fff7febefd3ffcb4fa6ff9c6f8b5f818f9;
    inBuf[10836] = 256'hedf90dfb5afcfcfddcffa601350368041d058305df054106a606eb06cf062d06;
    inBuf[10837] = 256'h06058203e5015a00ebfe9bfd68fc53fb79fa05fa1afabdfacffb11fd3efe37ff;
    inBuf[10838] = 256'h0600bb0077014402f1023d03f702f601520079fee1fcdbfb95fbf9fbc6fcc0fd;
    inBuf[10839] = 256'hcafee7ff27018202d103e4048b05ba059b0560053305340556055d0507052a04;
    inBuf[10840] = 256'ha4027f0000fe7cfb3ef9a1f7e1f6f5f6c4f730f9eafaadfc62fedbffe7009001;
    inBuf[10841] = 256'hf0011e025402bf024e03d503250403044e033102ff00f9ff5bff53ffd2ffb400;
    inBuf[10842] = 256'he80146039404ba059806fe06d9063106060559034501fcfeb9fccffa8ef908f9;
    inBuf[10843] = 256'h20f999f911fa40fa38fa2ffa77fa6dfb2efd82ff01021f046e05df059a05f104;
    inBuf[10844] = 256'h4104b20356033903380349038a03e8032d042c04b103ab024f01e4ffc3fe44fe;
    inBuf[10845] = 256'h8efe8effee002c02dd02bc02c7015e0001ff0cfeb0fdddfd26fe18fe83fd71fc;
    inBuf[10846] = 256'h1efb08faabf92cfa73fb33fde8fe2f00fe00880129023d03cf04b806aa083a0a;
    inBuf[10847] = 256'h3e0bbd0bac0b050bbb0994078604ee0054fd56fa7ff8eff758f837f915fab4fa;
    inBuf[10848] = 256'h19fb76fb06fcdcfcf3fd3cff75006601f60106029d01f20024005effdbfea0fe;
    inBuf[10849] = 256'h9dfeedfeb3ff0d01150398051508fe09e10a890a2c094c07740509041c037202;
    inBuf[10850] = 256'hb701bb0078ff17fed6fccefbe2fadff9a8f866f785f66cf655f732f9abfb4cfe;
    inBuf[10851] = 256'hb700b9023a043605b105bb055905b6041e04bf039703920385034303dd028402;
    inBuf[10852] = 256'h5b0289020b039e03080437041d04be034903d60246028401920066ff11fec8fc;
    inBuf[10853] = 256'hb2fbdafa43faeaf9c9f9dcf924faabfa6cfb5cfc70fd9afec5fff2002a027903;
    inBuf[10854] = 256'hd6042c06680772082b099a09ca09b1095609b5089e0701060004c301a1ffeefd;
    inBuf[10855] = 256'hbffcfefb7afbedfa43faa0f93cf94cf9ecf904fb5dfcb4fddbfec9ff83002501;
    inBuf[10856] = 256'hc2014b02b102fd02290342037903e0036004e3043d053105ac04d503f7027302;
    inBuf[10857] = 256'ha602ac034605f30624086e08a207d8056d03b900f6fd58fbf1f8c7f60df502f4;
    inBuf[10858] = 256'hb8f335f467f526f76cf934fc65ffdc023006dd08aa0a950bb60b610bcb0adc09;
    inBuf[10859] = 256'h8008b806910455026100f0fe16fec8fde2fd58fe41ff9e004102d303ec042d05;
    inBuf[10860] = 256'h840434039a0103008dfe28fdb9fb39fac8f8baf75bf7c4f7e8f893fa7bfc70fe;
    inBuf[10861] = 256'h51001702e203b7057c071709730a750b0d0c2f0cd40bed0a70097107ff043102;
    inBuf[10862] = 256'h5cffcdfcaefa4af9bbf8cbf84af901faa9fa33fbc5fb93fcc5fd4cff0701b402;
    inBuf[10863] = 256'he60370046204ca03e9020b0238017500d0ff3bffc3fe91febefe58ff48006d01;
    inBuf[10864] = 256'hc00220048205f506500860090e0a1a0a5a09e407cd053d038800f1fdb4fbe6f9;
    inBuf[10865] = 256'h7cf869f788f6d9f59af5e8f5e5f6b1f80bfb90fdecffc4010f030904d104a205;
    inBuf[10866] = 256'h850635079507710798066705300408034302eb01ba01b901ec015b0229031d04;
    inBuf[10867] = 256'hf1045905e304a103da01adffc7fd6bfc35fb5bfa8ef92af8fef6f4f59df4b1f5;
    inBuf[10868] = 256'h11fa99fd9bfe41ffcdffbeffd6fff8ffdefff0ff0400faff0d000e0005001900;
    inBuf[10869] = 256'h15000d0017000800ffff0300f0ffe6ffe9ffdfffe9fff9fffbff07000e000a00;
    inBuf[10870] = 256'h11000e00020004000100fdff0400050002000300fcfff9fffbfffaffffff0200;
    inBuf[10871] = 256'h03000c00130014000f000000f7fff4ffebffeffffafff5fff4fff9fff3fff3ff;
    inBuf[10872] = 256'hf7fff4fff7fffbfffcff0300030004001100160015001f002100190018001100;
    inBuf[10873] = 256'h08000600fffffafff8ffeeffe6ffe3ffe1ffe5ffe6ffe4ffeaffeefff5ff0600;
    inBuf[10874] = 256'h0e000e00130014001000120011000e000c000600faffeeffe5ffe9fff6fffeff;
    inBuf[10875] = 256'h01000100ffff020009000f000f0011000f000300f7fff7fffbfffeff05000a00;
    inBuf[10876] = 256'h0b000b0008000100fcfffafffefffefff8fff7fffcffffff0300050006000c00;
    inBuf[10877] = 256'h0a00fdfff7fff6fff2fff3fff6fff6fff6fff3fff3fff6fff4fff6fff9fff4ff;
    inBuf[10878] = 256'hf2fff9ff000006000c000c000d0014001c0020001f001e001d0011000300feff;
    inBuf[10879] = 256'hf9fff4fff1ffebffe5ffe4ffe6ffeaffedfff4ff02000b000c00140016000e00;


         
    encBuf[0] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[1] = 256'h0008000800080008000800080008000800080008000800080008000800080008;    
    encBuf[2] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[3] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[4] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[5] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[6] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[7] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[8] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[9] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[10] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[11] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[12] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[13] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[14] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[15] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[16] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[17] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[18] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[19] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[20] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[21] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[22] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[23] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[24] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[25] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[26] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[27] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[28] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[29] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[30] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[31] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[32] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[33] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[34] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[35] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[36] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[37] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[38] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[39] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[40] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[41] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[42] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[43] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[44] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[45] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[46] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[47] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[48] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[49] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[50] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[51] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[52] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[53] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[54] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[55] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[56] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[57] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[58] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[59] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[60] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[61] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[62] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[63] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[64] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[65] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[66] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[67] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[68] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[69] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[70] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[71] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[72] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[73] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[74] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[75] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[76] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[77] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[78] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[79] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[80] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[81] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[82] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[83] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[84] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[85] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[86] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[87] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[88] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[89] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[90] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[91] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[92] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[93] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[94] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[95] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[96] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[97] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[98] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[99] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[100] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[101] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[102] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[103] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[104] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[105] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[106] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[107] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[108] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[109] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[110] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[111] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[112] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[113] = 256'h0008000800080008000800080008000800080009010800080008000800080008;
    encBuf[114] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[115] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[116] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[117] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[118] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[119] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[120] = 256'h0008000800080008000800080008000800080008080000080008000800080008;
    encBuf[121] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[122] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[123] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[124] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[125] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[126] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[127] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[128] = 256'h0008000800080008000800080008000800080008000800080008000800080008;
    encBuf[129] = 256'h0008000800080000080800080009010800080008080000080008080801080008;
    encBuf[130] = 256'h0008000800090108000800080008000901080008000800090108080801080008;
    encBuf[131] = 256'h0009010800080008000800080008000800080000080800000900000800080008;
    encBuf[132] = 256'h0008000800080008000808080100090000080800000009000008080000080008;
    encBuf[133] = 256'h0008000800080008080000080008000800080800000800000900000800080008;
    encBuf[134] = 256'h0008000800080008000800080008000800080008000808080100080900000008;
    encBuf[135] = 256'h0008000901080008000800090100080800080008000800080008000800080000;
    encBuf[136] = 256'h0908010808000008000800080008000800090100080800080009010008080801;
    encBuf[137] = 256'h0808000800080000090000080008000800080008000800080008000800000900;
    encBuf[138] = 256'h0008000800080008000800080008080000080008000900000008000800080008;
    encBuf[139] = 256'h0008000808000008000800080000090000080008000800000908010808080108;
    encBuf[140] = 256'h0008000800090100090000080008000800080008000800080008000800080008;
    encBuf[141] = 256'h0008000800090108000800080008000800080008000800080008000800080008;
    encBuf[142] = 256'h0008000800080008080000080008000800080008000800080008000008080008;
    encBuf[143] = 256'h0008000800000900000009080108000800080008000808080108000800080008;
    encBuf[144] = 256'h0008000008080008000800080008000800080008000901080009010800090108;
    encBuf[145] = 256'h0008000800080009010008080800000800080000090000080800000009010908;
    encBuf[146] = 256'h0108000800080008080000080008000800090000000800080008000800080808;
    encBuf[147] = 256'h0100090000080008080801000900000900000008000800080008000800080008;
    encBuf[148] = 256'h0008000901080008000800080008000009000008000800080008000800080008;
    encBuf[149] = 256'h0800000800000808000800080008000009000008000800080008000800080008;
    encBuf[150] = 256'h0008000800080808010009080008010800080008000800080008000800080008;
    encBuf[151] = 256'h0008000800080008000800080008000800080009000000080800000800080008;
    encBuf[152] = 256'h0008000800080008000800080008000800090100080800080008000800080000;
    encBuf[153] = 256'h0808000800080008000800080008000800080008000800080008000800080008;
    encBuf[154] = 256'h0008000008080800000800080008000800080008000800080008000800080008;
    encBuf[155] = 256'h0008000800080008000009000008000800080008000800080008000900000009;
    encBuf[156] = 256'h0000000800080008000901080008000008080008000800080008000009000009;
    encBuf[157] = 256'h0000000800080008000800080008000800080008000800090108080801000908;
    encBuf[158] = 256'h0108000800080008000800080000090800000008000800090000000800000900;
    encBuf[159] = 256'h0008000800080008000800080008000901080008000800080008000800080008;
    encBuf[160] = 256'h0000090000080008000800080008000800080000090000080008000009000009;
    encBuf[161] = 256'h0108000800080008080801090100090000080808000800000008000009080100;
    encBuf[162] = 256'h0908010800080008000009080108000800080008000900000008000008080009;
    encBuf[163] = 256'h0108080000080008000901000900000008080800000009000009000000080008;
    encBuf[164] = 256'h0008000800080008000901000908010800080008000800080000090000080008;
    encBuf[165] = 256'h0008000800080008000800090000000800080808010800090000000800080008;
    encBuf[166] = 256'h00080000090800080908030603090f0b02010c0a03030103020c0e0801010200;
    encBuf[167] = 256'h0809000001040401090e0c0205080f09000109020400090001080b0908000109;
    encBuf[168] = 256'h0b090101090e0d0902000c0207030801020d0e0802010a0a0901010200000009;
    encBuf[169] = 256'h0901040403090f0d01020103040a0d01030b0f0a02020100080900000808090b;
    encBuf[170] = 256'h0c0808000706090802090e00040a0b0707070108000808080000080000080808;
    encBuf[171] = 256'h09090908090801000900000a0c0a0a0a0005030008090a010202080102000407;
    encBuf[172] = 256'h0603030208090800080305030402000801000a0b090b0c0004010800090d0b0b;
    encBuf[173] = 256'h0c0d09090a0900080b0b0b0f0d090908000100000001000001080a0802020607;
    encBuf[174] = 256'h0302030401000108080002040404020108080b0c0908080000090b0c0c0b0b0a;
    encBuf[175] = 256'h0b0c0b0b0c0b0b0c0e0b0c0a0801010108090b0d090801020304020101010203;
    encBuf[176] = 256'h030203020304030200000800040702080b0f0f0c0b0a080808080a0c0c0c0b0b;
    encBuf[177] = 256'h0a09080809080909090a0a0c0c0a090104040201000a09010406030403010000;
    encBuf[178] = 256'h020404030201000909090a0c0d0d0c0b0a0a090a0c0d0c0b0c0a090909090b0a;
    encBuf[179] = 256'h0c0b0a0b0a0c0a0a0a0908080a0c0c0b0a000206040304020202020305030403;
    encBuf[180] = 256'h0301000809090908090a0c0d0b0c0b0a0a0a0b0b0b0b0c0c0d0d0c0b0c090a08;
    encBuf[181] = 256'h090a0c0b0b0b0a0a0a0b0c0b0908020404030201000808000405040503020201;
    encBuf[182] = 256'h080a0c0b0a09010202080a0f0b0b0c09080809090b0d0d0b0b0a080001080a0f;
    encBuf[183] = 256'h0c0c0b0a090102050302080a0c0c0a0902050403030108090b0a080103050303;
    encBuf[184] = 256'h0301080a0d0b0b0b0a0009090d0e0c0a0b090008080b0d0d0b0a0a0800010101;
    encBuf[185] = 256'h01080c0d0a0b0902030603030101080001010305040404020203000101020404;
    encBuf[186] = 256'h020100090b0b0b09080a0a0a0e0b0b0e0c0b0d0b09080801080a0c0c0b0a0909;
    encBuf[187] = 256'h000a0a090b080201050402030503040401030303050502030301000008090008;
    encBuf[188] = 256'h00030405030201080b0a08090103090d0d0e0b0a0a0b0a0d0b0b0a0900080000;
    encBuf[189] = 256'h0a08040406030302030304040302030102040403050201000800010100010909;
    encBuf[190] = 256'h010107040201000b0b0a0a0a090f0b0c0c090909090a0c0b0a09000203050403;
    encBuf[191] = 256'h0404030402020304030503020100000103050403030201080808090809090908;
    encBuf[192] = 256'h000101090f0c0e0c0a0909000808080b0c0b0a0a080808010800000104060405;
    encBuf[193] = 256'h04030403030303030502020302020204040304030200000a090a0a0a0a0a0909;
    encBuf[194] = 256'h080100080d0f0d0c0b0b0b080003040302080a0c0e0b0a0a0801040504030302;
    encBuf[195] = 256'h0100000001040405030402000008080800010202010009090801020503020108;
    encBuf[196] = 256'h0b0c0c0b0900020302090f0d0c0a090003060302020000090a08010207050404;
    encBuf[197] = 256'h0201000a0b0c0a08010303040200080a0b0c0a0b09080003040203040101080b;
    encBuf[198] = 256'h0c0b0d0901010404010201000202030503030504040503030301000008010403;
    encBuf[199] = 256'h03040108090b0d0b0c0a08000102010a0d0e0c0b0a0909090900080900090b0b;
    encBuf[200] = 256'h0f0b0a0908000009080808060503040108080a0a010406050303040200000a0a;
    encBuf[201] = 256'h09090104030303000908090900090d0a0c0a000000000b0f0a0c0b0a0b0b0b0d;
    encBuf[202] = 256'h0a09000002090c0c0d0c090a0900080a08090a090a0c090b0b01020204000a08;
    encBuf[203] = 256'h0a0903090e0c0d0c08010406030201090b0b0c09010203060200010909080908;
    encBuf[204] = 256'h010102040100030101050200010b0f0d0c0d0a0a0900000101090e0c0e0b0a09;
    encBuf[205] = 256'h0901010101080b0c0c0c0a090901010001090b0c0c0b08080002010101020205;
    encBuf[206] = 256'h0304040202020202030303040303040201090c0c0b0b0a08080800090c0b0d0c;
    encBuf[207] = 256'h0b0c0b0b0c0b0d0c0a0b0a09080a0c0d0d0c0a0a0900000100090b0d0b0a0a09;
    encBuf[208] = 256'h080102030201090c0d0b0901030503010a0c0c0a09000103040100090b0c0b09;
    encBuf[209] = 256'h00060505030202000a0a0a090307030302000a0c0b09000205020208090a0a09;
    encBuf[210] = 256'h09080a0c0b0d0d0b0b0e0b0b0b0a080000090f0d0c0b0a090003020100090b0c;
    encBuf[211] = 256'h0b0a090102060403030200080909010504040402020201030203040201000000;
    encBuf[212] = 256'h0101010100090a0b0f0d0c0c0a090800030101090e0c0b0c090900020201080a;
    encBuf[213] = 256'h0f0b0c0a09080103030201000a0a0a0a01030505030201010908090900000800;
    encBuf[214] = 256'h080d0c0b0d09080801010a0b0c0e09000307050202010809090a010205040302;
    encBuf[215] = 256'h01000a0b0a0803070503030200080a090a0908000800090c0c0e0c0b0b090801;
    encBuf[216] = 256'h00000b0f0c0c0a09080001080a0b0c0c09090801010304040303020008000307;
    encBuf[217] = 256'h0504020301000000000100010101030503030308090a0c0a0102050303020008;
    encBuf[218] = 256'h0a0d0e0c0c0c0a0909000008080a0b0b0b0b0b0900030605030402010008090a;
    encBuf[219] = 256'h0a09090002060304040108090c0b0a09020504040201080a0b0d0b0b09000305;
    encBuf[220] = 256'h040101000a0b0a0b08020506040302020008090a080102050303020201000202;
    encBuf[221] = 256'h04020201090a0c0a0a000101000d0f0f0d0b0c0a090900010201080a0c0c0b0b;
    encBuf[222] = 256'h0901030504020000090a09080204050402020208000002040604030201000808;
    encBuf[223] = 256'h010204040202080b0b0d0a0a09080008090a0c0d0b0c0b0908020403010a0d0d;
    encBuf[224] = 256'h0b0b080003030200090b0d09080307040303030000090800030505030301080a;
    encBuf[225] = 256'h0c0b0a0a080202040100090c0b0c090900000800090800020503030101090a0c;
    encBuf[226] = 256'h0d0b0900070604040200000a0a09010305050202010809090a0a090a09000801;
    encBuf[227] = 256'h010a0c0f0c0c0a0a09080808080a0a0a0b0a0a09080801030505040403030302;
    encBuf[228] = 256'h02020101020102030405060303030100090a090306050403020208090c0e0b0c;
    encBuf[229] = 256'h0b0a090100000a0d0e0c0a0a090000000001000202020008090a080103060200;
    encBuf[230] = 256'h080a00020504030008080803070603030200000a09090800000100090d0d0d0c;
    encBuf[231] = 256'h0b0c0a0a080800090a0c0c0a0a09080101010201000101010304040304020302;
    encBuf[232] = 256'h02010305060305030202010809090908010201090f0d0b0c0a0909090a0b0d0b;
    encBuf[233] = 256'h0c0a0a0b0a0a0a0b090909080909080003070404040203030204020303040102;
    encBuf[234] = 256'h030103040304030101090b0e0b0d0a0a0a0a090a0c0d0d0b0d0b0a0a090a090a;
    encBuf[235] = 256'h0a090a08080809090b0a01050604030302010303030503020202020505040303;
    encBuf[236] = 256'h020100000001020101080a0b0e0b0d0c0c0d0b0c0b0b0a0b0a0b0b0c0b0a0b0a;
    encBuf[237] = 256'h0909000204060304030101000908090000020304040402030200000809000204;
    encBuf[238] = 256'h07050304010100090b0b0d0c0b0b0c0a0909080809090b0a0901040603020100;
    encBuf[239] = 256'h080a090a09080a000909090b0f0e0c0c0c0a0a09000203040202010100080809;
    encBuf[240] = 256'h0a0a090802060603050302030101000000030305030401020808090b0f0b0d0b;
    encBuf[241] = 256'h0c0c0b0b0c0b0b0a0b0a0909090a0900000204030200090a0b0b080207050504;
    encBuf[242] = 256'h040303030100080a090901030504030101080a0c0d0d0b0d0b0b0c0a0a0a0909;
    encBuf[243] = 256'h0a080a090b0a0c0b0c0a0a080205060404040303030303020100080909090003;
    encBuf[244] = 256'h0505020200090c0c0c0c0a0b0b0a0a090908090b0d0c0c0a0b0a09090a0b0c0c;
    encBuf[245] = 256'h0b0b09010206040304020202020102040404050303020201080a0a0c0b0c0a0a;
    encBuf[246] = 256'h0a0a090909090b0b0d0b0b09000206030202090b0d0d0b0b0a0a090002030403;
    encBuf[247] = 256'h01080c0d0b0a0804060404030202010100000808080908080001030403030304;
    encBuf[248] = 256'h04030201080b0c0b080106040301000808010606040403020101010205030502;
    encBuf[249] = 256'h01000909090a0908080909090001040303000809080407070304030201000a0c;
    encBuf[250] = 256'h0c0c0a0a0a0909090a0b0b0b090a0a0c0f0d0c0b0a090001010100080a0b0908;
    encBuf[251] = 256'h0800090a0b090307070703020202020101020101000a0b0c0b09010307030202;
    encBuf[252] = 256'h08090b0b0b0a0a080909010407050404020108090c0b0b0b0b09090001020503;
    encBuf[253] = 256'h040402000008090808020102030101020108020b0d0c0f0e0b0d0c0a0b090801;
    encBuf[254] = 256'h04050305020101000809080908080801010305040304030201080809090b0a0c;
    encBuf[255] = 256'h0b0c0a0a000405050301010a0c0d0c0c0b0b0a0a080003040302080a0f0d0c0b;
    encBuf[256] = 256'h0d0a0a0b09090a0a090b00010407040304010000000003050603050302030302;
    encBuf[257] = 256'h020108090a0a08010506050303040100080a0c0c0d0b0b0c0a0b0a0a090b0c0c;
    encBuf[258] = 256'h0c0c0b0c0a0b0909080001030305030403020303020303050305030502030303;
    encBuf[259] = 256'h02010008090b0c0c0c0b0b0b0b0a0b0b0c0d0b0d0c0b0b0b0c0a0b0909080102;
    encBuf[260] = 256'h0203030301010800000204050504030503030303030301010100080101020303;
    encBuf[261] = 256'h0302000a0c0e0d0c0c0c0c0b0c0b0b0c090a0809000800080809090800010404;
    encBuf[262] = 256'h060305040303040202020101010001010000000a0a0b0c0c0b0c0c0c0c0c0b0c;
    encBuf[263] = 256'h0b0b0a0b0a09090801010102000000090908020406050303030100000a090800;
    encBuf[264] = 256'h020703050503040302040304040403040304020201010809080a090909090b0d;
    encBuf[265] = 256'h0d0c0d0b0d0b0b0b0c0a09090900080001000101030404050304030305020303;
    encBuf[266] = 256'h0303020202010000090a0a0c0b0b0d0b0c0b0c0c0b0c0b0b0c0a0a0a0a080800;
    encBuf[267] = 256'h00020103020203020203030303030403040203020108090c0d0c0b0c0b0a0a00;
    encBuf[268] = 256'h01040504040203030202010101020204040303030100090d0d0d0c0c0c0b0c0b;
    encBuf[269] = 256'h0b0a0b0a0a090a090a0808000103040504040403040403030304020202020101;
    encBuf[270] = 256'h01000808090a0a0c0b0c0c0b0c0c0b0b0d0a0b0a090a08090800080100000108;
    encBuf[271] = 256'h000000020505040403030402030303030503030303020201020201030101000b;
    encBuf[272] = 256'h0e0e0c0c0c0c0b0c0b0b0b0c0a0a0a0b0b0c0b0c0b0a09080001020304040304;
    encBuf[273] = 256'h0305030204020202020203030203010100080a0b0c0e0c0c0b0c0b0c0a09090a;
    encBuf[274] = 256'h09090b0a0c0b0b0c0a0b0a0b0a09080002020401020000080101050504040403;
    encBuf[275] = 256'h03050304030403030202020100000809090a0b0c0c0b0d0c0c0d0b0d0b0b0b0c;
    encBuf[276] = 256'h0a0a08090800010102030305020403030404040403040302030302010100080a;
    encBuf[277] = 256'h0b0e0b0c0b0c0a0c0a0c0a0c0b0b0b0c0b0a0909080001020402030303030204;
    encBuf[278] = 256'h030305040201020808090b0c0909010405040503020303020404050604040404;
    encBuf[279] = 256'h03030303010000090a0a0a0b0a0a0c0b0e0c0c0d0b0c0b0b0b0a0a0800000201;
    encBuf[280] = 256'h03030303050403050303050302040302030302020000080a0b0c0c0b0c0b0b0b;
    encBuf[281] = 256'h0b0c0b0b0c0c0b0b0b0b0b0a090801010204020303020201000a090c0c0a0b0b;
    encBuf[282] = 256'h0909090000080000090b0b0c0a00040707050403040203030101010008090909;
    encBuf[283] = 256'h0909090a0a0d0c0d0d0b0d0c0a0c0a0a0a090a08080000020203050204030303;
    encBuf[284] = 256'h05030304040302030303020108080b0c0c0c0b0b0b0a0b0a0a0a0a0a0b0b0c0b;
    encBuf[285] = 256'h090901030505040304030302010009090a0c0b0c0b0b0b0c0a09080801020103;
    encBuf[286] = 256'h02030405040404030403040304020101080a0d0c0d0b0c0a0b0b0b0b0c0b0b0b;
    encBuf[287] = 256'h0c0b0c0a09090801020404040203030203030402030202010108090a0a0c0c0b;
    encBuf[288] = 256'h0d0b0d0b0c0c0a0b0b0a0b0b0a0a090800010201020001010203050203010008;
    encBuf[289] = 256'h090b0a090e0b0e0d0c0a0b090001040403030402040403040402030202020101;
    encBuf[290] = 256'h010109090b0d0c0c0b0d0b0b0d0b0b0b0b0b0a090a0900000105040404040304;
    encBuf[291] = 256'h0203020202020303050203020101090a0c0d0c0c0b0d0a0b0a09090909090a0a;
    encBuf[292] = 256'h09090908010001020204060305030201080a0d0c0b0d0b0b0b0b0a0a09010204;
    encBuf[293] = 256'h0404020303020405040704040503050303040201010008090a0a0b0a0a0a0b0c;
    encBuf[294] = 256'h0d0c0d0b0d0b0b0b0a0a09080002020304020303030404030503040303040303;
    encBuf[295] = 256'h0302020200090a0c0b0d0b0c0a0a0b0a0a0a0a0b0c0b0c0a0b0a0a0908010203;
    encBuf[296] = 256'h0304030200000a0d0b0e0c0b0b0c0a0b09090801020203030303030404040504;
    encBuf[297] = 256'h04040403020303020000090b0c0c0b0b0b0b0c0b0b0c0b0d0b0c0b0c0b0b0b0a;
    encBuf[298] = 256'h0a08000203050305030402030203020302030305030503050203020100090a0c;
    encBuf[299] = 256'h0b0c0b0b0a0a09090908090b0b0e0c0c0b0a0a08000305030402020200000809;
    encBuf[300] = 256'h0a0b0c0b0a080206050403030303020302020203020102030304030501080c0e;
    encBuf[301] = 256'h0d0d0b0c0b0b0b0b0b0b0a0a0a090909090a0b0b0b0802070504040303030402;
    encBuf[302] = 256'h020202010109090a0a0b0a090a090c0d0d0b0d0b0b0b0c0a0b0a0b0909010104;
    encBuf[303] = 256'h02030100090b0b0c090a0a090a0b090801050304010a0e0c0c0a080205040503;
    encBuf[304] = 256'h020302030202010108090a090908010201090c0f0d0b0c0b0c0a0a0b0a0b0a09;
    encBuf[305] = 256'h000205040403040302030302030303030303040402020208090c0e0b0c0c0a09;
    encBuf[306] = 256'h0909080909090b09090a0808090b0b0c0c0a0a0901030404050201000b0e0d0c;
    encBuf[307] = 256'h0d0a0b0c0a090909080900000801040306050403040304050306040305030402;
    encBuf[308] = 256'h02020008080a0b0a0b0b0b0a0b0d0b0e0c0c0b0c0b0b0b0a0800020203040303;
    encBuf[309] = 256'h03030304040304030404020402020302010000090b0b0d0c0b0b0b0a0b0a0909;
    encBuf[310] = 256'h090a0a0c0b0c0b0b090901010203020100090b0c0d0e0b0d0b0c0c0a0a0a0808;
    encBuf[311] = 256'h01020305030403030303030303050404030403020200080b0c0c0b0d0a0b0b0b;
    encBuf[312] = 256'h0c0a0b0a0b0b0b0c0b0b0c0a0b09090801020405040404020303010101080800;
    encBuf[313] = 256'h000102030305030201000a0c0d0c0b0a0b080801020303030503030404020101;
    encBuf[314] = 256'h0000010104030402000a0c0d0d0c0b0c0c0b0c0b0a0908010102020203020403;
    encBuf[315] = 256'h0504030304020302040204020201090a0d0c0b0c0a0b0a0a0a0b0a0a0a09090b;
    encBuf[316] = 256'h0d0c0c0b0a0901020403030108090b0c0b0b0b0d0c0c0b0c0a0a090000000008;
    encBuf[317] = 256'h000103050504020302020203050404020300080b0d0c0c0b0b0b0b0c0b0c0b0b;
    encBuf[318] = 256'h0b0a090909090a090802060504040302030302030303020208090c0b0b0a0a08;
    encBuf[319] = 256'h080a0c0d0c0c0b0b09090908080808010305050403030201000000000000080a;
    encBuf[320] = 256'h0c0b0d0a090a08090c0c0b0e0a090002050403030303040303040301000a0d0c;
    encBuf[321] = 256'h0b0c0a090a090a0b0e0c0c0c0c0a0c0a0a0a0a09080800010202030305040504;
    encBuf[322] = 256'h040403050204030404040304030202010009090b0c0b0b0b0b0c0b0c0c0c0c0b;
    encBuf[323] = 256'h0c0b0b0b0a090801030403040303030402040303030403030303040302020200;
    encBuf[324] = 256'h090a0d0c0b0c0c0a0a0a090808000108090a0c0b0c0b0909000008080a0c0c0c;
    encBuf[325] = 256'h0c0b0c0b0c0b0c0b0a0b0a080002040504040304030303020202020303040402;
    encBuf[326] = 256'h0200080b0d0c0c0b0c0b0b0b0b0a0b0b0b0a0a0a0a0a0a0a0909000203050404;
    encBuf[327] = 256'h04040305030303020100080a0909080203060403030303020200000008000205;
    encBuf[328] = 256'h06040404020108090b0d0c0a0b0a0b0a0a0a09090908090a0c0b0d0a0a000306;
    encBuf[329] = 256'h0503040303030402030402010100090909090908090a0c0d0c0c0b0c0b0b0c0b;
    encBuf[330] = 256'h0b0b0b09000203050202010808090a0808080008090808010303080e0f0e0c0b;
    encBuf[331] = 256'h0b0a09080000020202040302040200080a0d0a0b0a080800000a0e0d0b0d0b0a;
    encBuf[332] = 256'h0a0a0b0b0c0c0a09080103040302030202040305030203030305040404030202;
    encBuf[333] = 256'h080a0c0d0b0b0a09080808080a09090900010108090c0a090107040503020201;
    encBuf[334] = 256'h0101020304030108090b0a0a020505030301080b0e0a0b0b0a0a0b0a0b090203;
    encBuf[335] = 256'h06040100080d0b0c0a09080000080b0d0d0c0b0b0a0909080a0d0c0b0c0a090b;
    encBuf[336] = 256'h090a0d0b0a0c0908090001080002040506050305040304050404040403030402;
    encBuf[337] = 256'h02000009090a0b0b0b0b0c0c0b0c0c0c0c0b0c0a0b0a09080002020403030304;
    encBuf[338] = 256'h020304020402030303020402030302030100090a0d0c0b0d0b0a0b0a0a080000;
    encBuf[339] = 256'h0000090b0c0d0a0b0b0a0a0a0b0c0d0b0d0b0b0c0b0b0c0b0b0b0b0a08000404;
    encBuf[340] = 256'h05040403040402030202010101010102010108090b0f0c0c0b0b0c0a0b0b0a0a;
    encBuf[341] = 256'h0a0a0809000000000000010102030402010100000203050503030200080b0909;
    encBuf[342] = 256'h0006050404040204030304030201000808080000020302000a0f0c0d0b0c0b0c;
    encBuf[343] = 256'h0b0b0c0a0b0a0a09080000010202030504050304040203040203020302010009;
    encBuf[344] = 256'h0c0b0d0c0b0a0b0b0b0a0b0b0b0b0b0b0b0c0b0b0a0a00020504040201000808;
    encBuf[345] = 256'h09090a0b0c0c0d0b0c0b0b0a0909000008000908000003070403040303040202;
    encBuf[346] = 256'h01000a0d0e0c0b0c0b0a0b0b0b0c0c0a0b0b0a09090909090008010404050403;
    encBuf[347] = 256'h03030302040202030101080909080002060202030100010800010808090f0d0b;
    encBuf[348] = 256'h0d0b0a0b0b090a0a090908020306050303030203050306040304030203020100;
    encBuf[349] = 256'h080b0b0d0b0c0a0a090809080809090a0d0b0b0c0a0900030604050403030302;
    encBuf[350] = 256'h00000a0b0c0c0b0c0b0b0b0b0c0b0b0d0c0c0b0c0b0b0a090001030603040304;
    encBuf[351] = 256'h02040302040305030603060304040302020101080a0a0b0b0c0b0b0b0c0b0c0c;
    encBuf[352] = 256'h0c0c0b0c0b0a0a09080101040303030402030303040303030403030304030304;
    encBuf[353] = 256'h0302010108090c0c0b0d0a0a0a09080001000009090c0d0b0d0b0b0c0b0b0c0b;
    encBuf[354] = 256'h0b0c0b0a0a0a0a0b0b0a0b0a0900020706030603040304020201010000000808;
    encBuf[355] = 256'h080808090a0b0c0c0c0b0b0b0b0b0b0a0a090800010203030302000c0c0e0c0b;
    encBuf[356] = 256'h0d0b0c0a0b0a0909000100010008080102060604050503050303030302020008;
    encBuf[357] = 256'h090a0a0b0b0b0b0b0a0b0d0d0c0b0c0b0a0a0908000101020203010200080a0a;
    encBuf[358] = 256'h0d0b0b0c0b0b0b09010307060304030303020000000801010305030403020100;
    encBuf[359] = 256'h0a0c0c0c0c0c0b0c0b0c0a0b0c0a0b0a0a0a0a0a090809080a0b0a0a01040704;
    encBuf[360] = 256'h03040202010009090a0a0a0a080002020202080809090b090b0c0a0b0c0b0d0f;
    encBuf[361] = 256'h0d0c0c0b0c0b0a0c0a0b0c0b0c0a090800010304040304020303020402040304;
    encBuf[362] = 256'h03040202020008090b0b0c0b0b0b0b0c0c0b0b0b0c0b0a0c0a0b0a0a09080003;
    encBuf[363] = 256'h04040404020303030403020100080b0c0b0a0a00010001020104060405040203;
    encBuf[364] = 256'h02000100000103040402010a0e0d0d0b0c0b0b0a0a0b0b0b0b0b0b0b0a0b0e0b;
    encBuf[365] = 256'h0c0c0a0909000204050403050305030305030304040305040304030302010009;
    encBuf[366] = 256'h0b0c0c0c0a0b0a0b0a0b0c0b0d0b0b0c0b0a0a09000203060304020303020202;
    encBuf[367] = 256'h0203030203030201030202040203020100090a0c0b0b0b0a0803040603020208;
    encBuf[368] = 256'h0c0e0c0d0c0b0c0b0c0b0c0c0a0b0b0a0a0a0809000000020204040404040304;
    encBuf[369] = 256'h040303030202010008090a0b0c0a0c0a0c0b0b0c0a0b0a090908000001010302;
    encBuf[370] = 256'h04030304020108090c0d0c0d0b0d0b0b0b0c0a09090801010304030404040304;
    encBuf[371] = 256'h030403030402020101010808080809090a0b0b0d0d0b0c0c0b0b0b0b0a0a0800;
    encBuf[372] = 256'h020202030303040203030503040402030202010000000809090b0e0c0b0b0c0a;
    encBuf[373] = 256'h08080002030402020200080a0e0c0d0c0b0b0b0a0b0a0b0d0a0b0c0a0a0a090a;
    encBuf[374] = 256'h090000030603050303030402020201000108080809090a0c0c0c0c0b0c0b0d0b;
    encBuf[375] = 256'h0c0b0c0b0b0b0d0b0a0c0a090a0909090909090a080808000008010001040101;
    encBuf[376] = 256'h010a09010407070503050203040202030202010001000000080b0d0d0e0b0b0d;
    encBuf[377] = 256'h0a0b0a0b0a0a0a080802040404050304030203030201000809090a0a0b0c0b0c;
    encBuf[378] = 256'h0b0a0b0b0b0a0a090304060404030403030302020100090a0c0c0b0d0a0a0a09;
    encBuf[379] = 256'h09080a0b0c0d0b0b0b09090808080a0a0a0a0a00090d0d0c0d0b0b0a08010305;
    encBuf[380] = 256'h040403040402050404050504040403040303010100090a0b0c0b0b0b0b0b0c0c;
    encBuf[381] = 256'h0c0c0b0d0a0b0a09090001020403040303030203020303030303020101010102;
    encBuf[382] = 256'h04030503030101090909090002050404020200080b0c0e0b0d0c0b0c0b0b0c0c;
    encBuf[383] = 256'h0b0c0b0b0c0a0908080001020201020303060403040304020302020101080909;
    encBuf[384] = 256'h0b0c0b0c0b0b0c0a0a0a090002040603050302020100090a0a0c0c0b0b0d0b0c;
    encBuf[385] = 256'h0b0c0b0c0b0b0b0b090900020404040304030404040304020302020000080a0a;
    encBuf[386] = 256'h0b0c0b0c0b0b0c0b0c0b0a0c0a0a09080104050404030303020100000009080a;
    encBuf[387] = 256'h0b0c0c0c0b0b0a0b0a0a090908000203070403040303030203010100080b0e0c;
    encBuf[388] = 256'h0c0c0b0b0a0a0b0a0a0b0b0a0b090001040404030503030303030100090a0a0c;
    encBuf[389] = 256'h0b0c0b0c0c0c0b0c0c0a090a0800000101020203040304030304020100090a0d;
    encBuf[390] = 256'h0d0c0c0c0b0b0c0a090a0a0a0a0a090800040405030502030304030203020101;
    encBuf[391] = 256'h08080a0c0b0d0c0b0c0b0b0b0a0a080800020303040503040303040201000808;
    encBuf[392] = 256'h09090908090a0d0d0c0c0a0b0a0a090908090001030504040305030303030302;
    encBuf[393] = 256'h01080a0c0c0b0b0a0a0b0b0c0d0c0b0b0b0a0900010201010000000102040303;
    encBuf[394] = 256'h01010a0d0d0c0d0c0c0c0c0a0b0a0a0800010103030503040403040403060405;
    encBuf[395] = 256'h04040403040202020808090b0c0b0a0b0a0a090b0b0e0b0d0b0c0a0a0a080002;
    encBuf[396] = 256'h0305030303020301020102020202010102020305030404030203010000090a0a;
    encBuf[397] = 256'h09080104030402010a0d0d0d0c0b0b0c0b0b0b0d0b0c0c0b0c0b0a0a0a090808;
    encBuf[398] = 256'h08000101020404040303040303030302010008090908090008090a0d0c0c0b0a;
    encBuf[399] = 256'h0901050504040203010108090b0d0b0d0b0c0b0c0a0b0b0b0c0a0b0a0a000104;
    encBuf[400] = 256'h040403040303040304030403030302010009090b0c0c0a0b0a0b0a0b0a0a0a0b;
    encBuf[401] = 256'h0b0a0a080205060403040202000008080909080909090b0d0b0b0c0a09080103;
    encBuf[402] = 256'h060405030403030202010008080a0a0b0e0b0e0b0c0c0b0a0b0c0a0b0a0b0a0a;
    encBuf[403] = 256'h090800010101010202060305030303010108080a0b0b0c0c0b0b0c0b0c0a090a;
    encBuf[404] = 256'h080000000108080008000200080a0f0c0d0c0b0c0c0c0b0d0b0b0c0b0b0a0a08;
    encBuf[405] = 256'h0800020204040204030403040304030304020201010108000809080909090900;
    encBuf[406] = 256'h01000101090a0c0d0c090a09000101030101010002050305030208090d0b0a09;
    encBuf[407] = 256'h0802000a0d0f0d0b0b0a010505040402030202020102030100080c0b0c0d0a0b;
    encBuf[408] = 256'h0b0c0b0c0a0a090801010202010008000803060405030200090c0f0a0a0a0908;
    encBuf[409] = 256'h090a0d0d0c0b0a0b090000020202030204040605050604040404030303020100;
    encBuf[410] = 256'h090a0c0b0b0b0a0b0a0a0b0d0c0c0c0b0a0b0908000204040304030202010100;
    encBuf[411] = 256'h0800080808080008000002030404030302020102030404050403030402020008;
    encBuf[412] = 256'h0b0d0c0c0b0c0b0c0b0b0c0b0c0b0c0a0b0a0a0a080900080001020306030404;
    encBuf[413] = 256'h0202020001080008090808000001020204020103010003050505040304030201;
    encBuf[414] = 256'h08090c0d0c0b0c0b0c0b0a0b0b0b0b0a0a0a0901020405040403040203020303;
    encBuf[415] = 256'h04030303020200080b0c0d0b0b0a0a0900020303050202010101030705050403;
    encBuf[416] = 256'h04020100090b0d0c0b0b0c0a090a090a09090909080001020404050404030203;
    encBuf[417] = 256'h010108090b0b0c0d0b0b0d0b0b0b0b0909000203040303040202010200000809;
    encBuf[418] = 256'h0a0b0e0c0b0e0b0d0b0b0c0a0a09090800000100020203040404030303030301;
    encBuf[419] = 256'h0008090b0c0b0d0a0b0c0a0b0b0b0b0a0b0c0a0b0a0901020404030303010001;
    encBuf[420] = 256'h0001020008080b0b080903060202020a0a090c01050307030202030101030203;
    encBuf[421] = 256'h040101020808010900050205050202010a0e0d0d0c0c0c0b0b0b0b0a0a0a0908;
    encBuf[422] = 256'h0801010203030404010203010303010102090a0a0f0b090c0a00000506040305;
    encBuf[423] = 256'h030203010000090b0b0c0c0c0c0c0b0d0c0b0b0c0a0a09090900000800010001;
    encBuf[424] = 256'h0202050404040403060405040404040403040202020008090a0b0c0b0a0a0b0a;
    encBuf[425] = 256'h0a0b0d0b0d0b0c0a0a080001040305030303010108080a0a0a0b090909080100;
    encBuf[426] = 256'h0203040404030403030503030404020303020108090b0e0c0b0d0b0b0b0c0b0b;
    encBuf[427] = 256'h0c0b0c0a0b0b0b0a0a09080800010102020201030203030201010a0b0e0b0b0a;
    encBuf[428] = 256'h0908010104030404040405030504030503040203020108090a0d0c0b0c0b0b0a;
    encBuf[429] = 256'h0b0b0b0b0b0a0a08000306040404040303020302010008000908090809090a09;
    encBuf[430] = 256'h0a09090800020406040403040302020202020202030100090d0d0c0c0b0b0a0a;
    encBuf[431] = 256'h09080001030404040304030303040304020301000b0d0d0d0b0c0c0a0b0b0b0a;
    encBuf[432] = 256'h0b0b0b0b0a0b0a0909090801010203030201010808090809090b0c0c0b0c0909;
    encBuf[433] = 256'h080101010201080c0d0d0c0b0a0a0908010000090a0b0c090900080a0d0d0c0c;
    encBuf[434] = 256'h0b0a0b0c0b0d0d0d0b0c0b0b0a0a090900000304050404030304030304030504;
    encBuf[435] = 256'h0203030201010100010101020000080b0b0c0d0b0b0d0b0b0b0b0a0b0a080901;
    encBuf[436] = 256'h030604050303050202020208080a0d0c0b0d0b0b0c0c0b0b0c0b0a0908000203;
    encBuf[437] = 256'h03050302030101000a090a0a09010205050302000a0f0c0d0b0c090900010203;
    encBuf[438] = 256'h0202090b0e0d0b0c0b0b0a0a090808000808090a0a0a08010407050504050405;
    encBuf[439] = 256'h0305040304030203020108090b0c0c0a0b0a090a090a0a0c0b0c0b0b0a090103;
    encBuf[440] = 256'h0604040303020108090b0d0b0b0b0a0908010304040304030303040302040303;
    encBuf[441] = 256'h0304020201000a0c0c0c0c0c0b0a0b0b0a0a0a0a090a0a0b0c0b0c0a0b0a0909;
    encBuf[442] = 256'h0900000800080a0a0c0e0b0d0b0c0b0b090a0800020305040203030303030403;
    encBuf[443] = 256'h0404040304040304020100090b0e0b0c0b0b0b09090000010001080008080002;
    encBuf[444] = 256'h05050404030303020000090b0a0c0a0b0a0b0b0b0b0a09000306040503040303;
    encBuf[445] = 256'h02020108000900000103030301090d0e0c0c0b0a090002040504030302030101;
    encBuf[446] = 256'h000100010008090b0e0d0c0c0c0b0c0c0b0b0b0b0c0a090a0908080801000000;
    encBuf[447] = 256'h08090a0b0d0b0c0b0b0b0b0b0c0c0b0b0d0a0b0a080001030503050303030202;
    encBuf[448] = 256'h0109090a0b0a0808000108090a0d0b0b0e0b0d0d0c0b0c0b0b0b0c0b0c0a0b0a;
    encBuf[449] = 256'h0908000103010203040405020303010101080801090801000106030505020203;
    encBuf[450] = 256'h030403010102090002010406030403040203020100090b0c0c0a080801020108;
    encBuf[451] = 256'h090d0d0d0d0b0c0c0a090900010101080b0c0c0c0a0808020503050402030201;
    encBuf[452] = 256'h010009090a0a0b090b0a0a0c0b0c0c0b0c0a0b090a09090908090a0a0c0c0b0d;
    encBuf[453] = 256'h0b0b0c0a09080103030404030306030406030504050404040404030403030202;
    encBuf[454] = 256'h0100090a0b0c0c0a0a0a0909090a0b0c0c0b0b0b0a0003050504030203000809;
    encBuf[455] = 256'h0b0e0b0b0b0a09080203060403030302030102010101020203020301080b0f0d;
    encBuf[456] = 256'h0b0d0c0a0b0a090a080800080008090b0c0b0d0b0a0b0a0b0b0b0b0c0a0a0909;
    encBuf[457] = 256'h0900090a0a0d0b0b0b0a0103050502010009090a090800020406040504040402;
    encBuf[458] = 256'h030101090a0c0c0b0c0a0a090000020202020008080800030704040402030302;
    encBuf[459] = 256'h00080a0c0c0c0b0b0a090908000808090800000103040302030108080a0b0901;
    encBuf[460] = 256'h03070503030200080a0c0b0b0a09010407040404030302030303040304020201;
    encBuf[461] = 256'h090a0c0e0b0e0b0c0c0b0b0c0a0b0a0a0a0a0908080808090a0b0b0d0b0b0a0a;
    encBuf[462] = 256'h0a090908090b0b0e0b0a09000206050304040304030302030201000000010102;
    encBuf[463] = 256'h040101080e0c0d0c0c0b0b0b0a0b0a090b0a0a0a0b0a0a090908000102050503;
    encBuf[464] = 256'h0503010100080002030704040403030303020203010303050304020201000000;
    encBuf[465] = 256'h080001090b0c0f0b0c0d0a0b0a0a09000103020404020202030204010008090a;
    encBuf[466] = 256'h0b0c0b0c0c0b0b0b0a09090a0b0e0c0a0a080305050402020000090a0a0a0a0a;
    encBuf[467] = 256'h0a0a0d0b0b0d0a090908000b0c0e0d0d0b0d0b0a0b0808010403040302020100;
    encBuf[468] = 256'h0809080103040604030304020403040503050403050303030402010008080a0b;
    encBuf[469] = 256'h0b0b0c0c0a0a0b0a0b0a090800020306040503040303040202010108090a0b0b;
    encBuf[470] = 256'h0a0a08010102030100090a0a0908040405040304030303040108000a0c0b0d0b;
    encBuf[471] = 256'h0b0c0c0b0b0e0c0b0d0b0c0b0a0a090900000202030304030303020303010108;
    encBuf[472] = 256'h0b0d0e0d0b0c0c0b0b0b0a0a0a080000020304050303050202020000080b0c0b;
    encBuf[473] = 256'h0d0c0a0b0b0a0a0908000102030503050404030403030202010000080a0a0c0c;
    encBuf[474] = 256'h0b0b0c0b0a0a0a0a0b090909080808000001040303050101080a0c0b0e0c0b0b;
    encBuf[475] = 256'h0c0b0a0900010205030403030404040404030402020200090a0c0e0b0d0b0c0a;
    encBuf[476] = 256'h0b0a0a0909090a0a0a0c0b0a0b09090808090a0c0b0d0b0b0b0b0b0d0a0a0b09;
    encBuf[477] = 256'h0900020405050404040203030201020202020100090a0e0b0d0b0c0c0a0b0c0a;
    encBuf[478] = 256'h0a0b090a0a0a0a0a0b0a0a0801040505040203020101090a0a0c0a0908020404;
    encBuf[479] = 256'h04030302010008000102060305030403030201000b0c0d0c0a0b090a09090b0b;
    encBuf[480] = 256'h0d0b0c0a0b090a0800010306040404030204020202020202020008090a0b0c0c;
    encBuf[481] = 256'h0a0c0b0a0c0b0a0b0b090a09080a0c0b0f0b0c0c0b0b0b0c0a0a0b0a0c0b0a0c;
    encBuf[482] = 256'h0c0a0a0a0908090108010205040603030303010200000100010202020208090b;
    encBuf[483] = 256'h0f0c0c0b0b0a0802060504050304030302030101000808080802020203010000;
    encBuf[484] = 256'h0801060505040403040303040304040203030203020102020102010201010000;
    encBuf[485] = 256'h090a0b0b0d080003070503050303030402020102010200010008090c0e0c0c0c;
    encBuf[486] = 256'h0b0b0b0a0a0a09090801020306030303020101090b0d0d0d0c0c0b0d0b0b0a0a;
    encBuf[487] = 256'h0a0808080008080008000102020200080a0c0b0c0c0a0b0b0b0b0b0c0c0c0c0b;
    encBuf[488] = 256'h0b0b090103050403020201000809090c0b0d0b0b0b0a080809090b0d0c0b0a00;
    encBuf[489] = 256'h040505030403020100080909090002040404010108090a080105060304040102;
    encBuf[490] = 256'h00080a0a0a0b090900010202040200080e0d0d0c0c0b0a0a0a090a0a0c0b0b0b;
    encBuf[491] = 256'h0a0a080102030503030403010201000a0a0e0c0b0d0a0b090800020306020402;
    encBuf[492] = 256'h030203010202000008090a090b080800010108090d0f0c0c0c0b0b0b0a090801;
    encBuf[493] = 256'h0204030300080a0d0c0a0c0a0a0b0c0b0d0b0909010204030303050304040302;
    encBuf[494] = 256'h020009090a0a0c0b0e0b0c0b0b0b090909090809090000010002020307060404;
    encBuf[495] = 256'h0304040201020008080a0c0a0c0b0c0b0d0b0d0c0a0b0b0b0909010103040203;
    encBuf[496] = 256'h0200010001020503030302000a0d0c0c0b0b0a0a0b0c0b0c0c0b0a0b09080004;
    encBuf[497] = 256'h0604040403030202010202020404030305020303030202020100010305050404;
    encBuf[498] = 256'h04030302040103030304040303050204030204020202010100080909080a0001;
    encBuf[499] = 256'h04060403040303030303040402040203020301020109090a0d0a0a0b08090901;
    encBuf[500] = 256'h0100030108000b0f0d0c0b0a0909010200020a0e0c0d0c0b0c0b0a0b0c0b0b0d;
    encBuf[501] = 256'h0a0a0b08090908090a0c0c0b0c0b0c0b0b0b0b0c0b0a0b0a0a0b0d0a0b0b0909;
    encBuf[502] = 256'h0901000801000001090c0c0f0c0a0b0b08080002010008090c0b0e0c0b0c0b0b;
    encBuf[503] = 256'h0a0900010405030402020000080a0a0a0a0a0a090908080809090c0c0d0c0c0b;
    encBuf[504] = 256'h0d0b0a0900030505040202020100000102030504030302020109090d0c0d0c0b;
    encBuf[505] = 256'h0c0b0c0a0b0a0a0a090a0909090a0b0d0c0c0b0c0a0b09090801020502030300;
    encBuf[506] = 256'h080a0d0b0c0b0a090808000809080b0a080005060403030208090e0b0d0b0b0b;
    encBuf[507] = 256'h0a0908000001090c0c0d0b09080205050305010200080a0a0c0c0a0a09000002;
    encBuf[508] = 256'h020208080c0c0c0b0b0a0a0800010206030403040204010202020101090a0a0d;
    encBuf[509] = 256'h0a0808010403020308090b0f0b0a0a09020206050203030008090c0c0a0a0901;
    encBuf[510] = 256'h0306040301010b0c0d0d0a0b0a08000002030302020108080809000908000c0c;
    encBuf[511] = 256'h0c0e0c0b0c0b0a0b0b0b0a0b090b090808020204050504040403030302010008;
    encBuf[512] = 256'h0800000305030503020201080808000307060403040304020202030203040302;
    encBuf[513] = 256'h0403030403030303020100080809080002020404030504040405030403040302;
    encBuf[514] = 256'h0101000808080900000800090c0c0c0b0c09090003050404030203010108090a;
    encBuf[515] = 256'h0c0b0b0c0b0a0b0a0b0d0d0b0c0c0b0a0b090a0a0a0a0c0a0c0b0a0a0a090909;
    encBuf[516] = 256'h090a0c0b0e0c0a0c0a0a0b0b0a0b0c0a0c0a0a0b09090801020202000c0f0d0c;
    encBuf[517] = 256'h0c0a0a09080102030301080a0d0c0b0a0900020404030302080a0e0d0c0b0b0b;
    encBuf[518] = 256'h0a09080801010101030303040201090c0c0c0a08010504050202080b0f0c0d0b;
    encBuf[519] = 256'h0c0a0a08010404050303030200090b0c0c0b090900010304030201080b0d0c0b;
    encBuf[520] = 256'h0a0a080205040403030200090b0e0b0c0a0a0800010402040201010809090b0b;
    encBuf[521] = 256'h0b0b09080001020301010008080003070404040302030100090a0c0c0c0b0b0b;
    encBuf[522] = 256'h0a09080800000808080800010303050200000b0e0b0e0c0b0b0c0a0b09090808;
    encBuf[523] = 256'h0000000101030504050304030304020201010108090809080102050403040303;
    encBuf[524] = 256'h03020203010100080808000207040305020200000a090a080103060404020201;
    encBuf[525] = 256'h00080a09080003060504040402030202010008090b0b0d0c0b0c0c0b0a0a0900;
    encBuf[526] = 256'h0103050203020101010001010002040305050404030402020101080800010205;
    encBuf[527] = 256'h050304040204020302040202030303030303020102000801010002020001080b;
    encBuf[528] = 256'h010203070707040302040202010108080808080100040403050302020109090b;
    encBuf[529] = 256'h0d090908040405040302020108080b0d0a0c0b0a0b0c090a0a09090a0a0b0e0a;
    encBuf[530] = 256'h0c0c0a0a0b0a0a0a090a09000909080b0e0b0e0c0b0b0c0a0b0a09090a090c0c;
    encBuf[531] = 256'h0b0d0c0a0b0b090a080000020200080a0f0d0c0c0b0c0b0b0b0b0b0b0a090908;
    encBuf[532] = 256'h08090a0b0e0b0d0a0c0a090a0a090a09090908080002020304010000090a080a;
    encBuf[533] = 256'h090a0f0e0c0c0b0b0b0a09090a090b0d0a0c0b0a0c0b0c0b0c0a0b0800020505;
    encBuf[534] = 256'h0404030304020202010000080b0a0b0b0a080104040303030001000801030505;
    encBuf[535] = 256'h050304030301000a0d0c0d0a0b0a090808000009090a0d0c0b0b0b0808020503;
    encBuf[536] = 256'h0503020303020305020403010201090a0c0d0b0b0c0b0a0b0b0b0d0a0a090802;
    encBuf[537] = 256'h03040401090c0f0c0c0b0c0a0a0a09080801080000090b0c0d0b0a0908030405;
    encBuf[538] = 256'h040303020201010000000000020102050101020001010101040800000c0a090a;
    encBuf[539] = 256'h00030102020b0b0b0f0d0a0c0b0a0d09080a0000080103030706030404030403;
    encBuf[540] = 256'h0304020303030303040202030203030304030102010001010307040405030304;
    encBuf[541] = 256'h0303040203020302030302020202040306040404030402030203030204030403;
    encBuf[542] = 256'h0503030503040402020100000a0b0b0d0a0a0909000000020000010001020504;
    encBuf[543] = 256'h040402030008090c0d0a0b0b0a0a0a0a0a0c0a0a0b0b0b0b0001040704030402;
    encBuf[544] = 256'h00000a0b0c0b0c0b0a0b0a0b0b0c0d0c0c0c0b0c0a0a090909080a0b0c0b0a09;
    encBuf[545] = 256'h09000100090a0e0b0c0c0a0a090800000101080a0c0e0c0b0b0b0b0b09090800;
    encBuf[546] = 256'h020202040100080b0d0b0e0c0b0c0c0b0c0c0b0c0c0a0b0a0908000001010100;
    encBuf[547] = 256'h00010203040301080a0d0c0b0b0a090001030503030201080a0d0b0b0c0a0909;
    encBuf[548] = 256'h0908080801090a0a0f0b0a090104040303080808000507030303090b0e0c0a09;
    encBuf[549] = 256'h0105050404030303030102000808080801020404030300080d0c0d0c0a0b0b0b;
    encBuf[550] = 256'h0a09080001030304030302010100000808010406050505030303030108090a0b;
    encBuf[551] = 256'h0b0a0a0808010203040202020201020103050404050305020200080c0c0d0c0b;
    encBuf[552] = 256'h0b0c090a090800080000090a0a0c0b0b0a090000020304040403040302040203;
    encBuf[553] = 256'h04040303030108090b0a0a00030504030300090d0d0d0c0b0b0c0a090909090a;
    encBuf[554] = 256'h0b0b0c0a0a09000003060306030402020100080a090808020301020101030707;
    encBuf[555] = 256'h0405030303030202010102020304020403040404030502020202010000000001;
    encBuf[556] = 256'h0002030204040204030403040203040204030405030305030202020008080a0a;
    encBuf[557] = 256'h0b0c090a0800020104020008090c0b0c0c0a0a0a0001010302080a0f0e0c0c0c;
    encBuf[558] = 256'h0a0b0b0a0909000000010809080b0a09000003040204020101090c0c0e0c0b0c;
    encBuf[559] = 256'h0b0b0b0d0c0c0c0b0b0c090a09090a0b0b0d0b0b0a0b0a0a0b0a0b0b0b0c0c0b;
    encBuf[560] = 256'h0c0b0c0b0b0b0b0b0b0a090908090b0c0c0b0a000406030301090e0d0b0d0a0a;
    encBuf[561] = 256'h0a0809090a0b0c0c0c0b0b0a0b0a090801020304050202030001080808000908;
    encBuf[562] = 256'h090e0c0c0c0b09090802020201080a0c0c0b080903060405030402030100090a;
    encBuf[563] = 256'h0b0b0c0a090908000a0a0b0e0b0a0b0900000002080104030706030504030302;
    encBuf[564] = 256'h0208080a0b0a0c0a080900020100000c0d0c0d0c0b0b0c090909090909090909;
    encBuf[565] = 256'h0100020300090a0f0b0b0b0b080a0a000a09020808020d0d0b0e0a0102070603;
    encBuf[566] = 256'h040303010100090a0a0908090800090b0b0f0b0a0b0c0a0d0b0b0b0b09080206;
    encBuf[567] = 256'h0305040202020101000808090908010405050304030302010800080001040404;
    encBuf[568] = 256'h0304030302030302040203040305040305020301010100000002040304020100;
    encBuf[569] = 256'h090a0a0a00030704040402020301010101020203040403050403040402030202;
    encBuf[570] = 256'h010100010101020303050402040304030302020109090b0c0a090a0801020505;
    encBuf[571] = 256'h0304040103010808090b0b0d0b0c0b0b0b0b0b09090b0a0c0c0a0a0a02040406;
    encBuf[572] = 256'h030101080b0c0c0c090900010108090c0f0b0c0b0b0b0c0a0b0c0a0c0a0b0a0b;
    encBuf[573] = 256'h0a09090002030703040303010208090a0b0b0a0b0a080c0c0c0e0c0a0c0a0a09;
    encBuf[574] = 256'h090800000808090b0e0b0c0a0a080103040301000b0f0c0d0b0b0c0a0b0b0a0a;
    encBuf[575] = 256'h0a0a090908080809090b0b0c0a09080801080b0c0f0b0b0b0a00000203010809;
    encBuf[576] = 256'h0d0b0a0b09000909080e0b0c0c0b0b0d0c0c0c0c0b0b0c090909010002020101;
    encBuf[577] = 256'h0009090909000504050503020200090a0d0b0a0a090002030603050302030301;
    encBuf[578] = 256'h010009090000030703040401010108090808000200090a0f0f0b0c0b0a0a0800;
    encBuf[579] = 256'h010103010201000001010104030406020303020100090b0a0c09020306050202;
    encBuf[580] = 256'h010a0b0d0d0b0a0b0a0a0a0b0b0d0b0c0c0b0a0b090100020301080a0f0b0a0b;
    encBuf[581] = 256'h0003050504020300080a0b0c0b0a080206040402030202000000090001000203;
    encBuf[582] = 256'h0404030203020001090901000407050306020303020203010203020305020504;
    encBuf[583] = 256'h0304050305030303030202010001020204050304040204020204020303040303;
    encBuf[584] = 256'h030203030203020102000808080a000000070403050402030202020301040402;
    encBuf[585] = 256'h05020203010000080a08090a000009030201050108000b0f0c0c0d0a0a0b0b0b;
    encBuf[586] = 256'h0d0a0c0b0c0b0d0b0b0d0a0c0a0b0a0b0a0a0a090a0b0a0b0d0b0c0b0b0b0908;
    encBuf[587] = 256'h0001030101080b0f0d0c0c0b0c0a0b0a0b0a0a0c0a0c0c0a0b0b0a0a0a090908;
    encBuf[588] = 256'h0909090a0d0c0b0e0b0b0c0b0b0c0a0b0a0b0b0b0b0a0a0a0808010201030304;
    encBuf[589] = 256'h05030504020302000a0a0f0c0b0c0b0a0a0a09080a090d0c0b0d0b0a0b090000;
    encBuf[590] = 256'h00020808090d0b0b0c0b0a0909080800010808000a09080a0904020607020403;
    encBuf[591] = 256'h030204010204020404020201080b0b0e0a090900020101010b0c0c0e0a090900;
    encBuf[592] = 256'h030305050202020101010101020202050203040204030203030201020808010a;
    encBuf[593] = 256'h09010903070405050203040001080a0b0b0c0a090801030302020b0e0c0e0b0a;
    encBuf[594] = 256'h0b090800000208080b0f0c0b0c0b0909000200010109090a0b0a020206050202;
    encBuf[595] = 256'h02080a0a0e0a0a0b09090a09090c0c0b0d0b0b0c0a0a0a08000800010808090a;
    encBuf[596] = 256'h0804060705030503020201000008000304050404020303020202010203040403;
    encBuf[597] = 256'h0404020304030403050303030403030304030403030303030403030304020302;
    encBuf[598] = 256'h0201020103050504040304030303030303050304040204020202030102020202;
    encBuf[599] = 256'h020103020003030305040104030102020001000a080b0f0a0b0e0b0b0d0b0b0c;
    encBuf[600] = 256'h0b0b0d0a0b0c0b0a0c0a0b0b0b0c0c090a0b08090900090b0a0e0c0b0b0d0a0a;
    encBuf[601] = 256'h0a0a0a0b0b0d0c0b0c0c0a0b0b0b0b0c0a0a0b0b0b0c0b0c0b0c0b0c0b0c0a0b;
    encBuf[602] = 256'h0b0a090a09000908080a0a090b0b080a0801000205020202090c0d0f0b0c0c0b;
    encBuf[603] = 256'h0a0b0a090800010102020002000908080900000103030103080d0d0e0d0c0b0c;
    encBuf[604] = 256'h0a0b09080002040403040201010809090a0900020307030204010000090b0c0c;
    encBuf[605] = 256'h0c0a0a0801010202090d0e0e0b0c0b0a090900000000080a0a0a0b0a00080103;
    encBuf[606] = 256'h0405040202040203040201020909090a0a000103070202020009080d0c0b0d0b;
    encBuf[607] = 256'h0a0a090101010408090a0f0b0b0c0a08000803000800090b0203060705020302;
    encBuf[608] = 256'h02010008020204070304040202030000000a0a090b0a00090a010a0d0a0e0c0b;
    encBuf[609] = 256'h0c0c090b0a080a09090c0a0a0c09080800020008090f0b0c0d09090901040204;
    encBuf[610] = 256'h030101000b0a0c0d09090800030205030304010108090b090a08060505050304;
    encBuf[611] = 256'h0302020101010002030405040303050202030202030202040302050304040303;
    encBuf[612] = 256'h0403020302010302020304030504020403020303020202010201020403040503;
    encBuf[613] = 256'h0204010100000900080803010305010101090a0a0e0b0a0c0a0a0c0b0b0e0c0a;
    encBuf[614] = 256'h0c0b0a0c0a0b0b0c0b0e0a0b0d0a0b0b0c0a0a0b0a0c0a0b0d0a0b0c0b0a0b0b;
    encBuf[615] = 256'h0a0c0b0b0c0b0b0c0b0b0d0a0a0b0b0a0c0a0a0c0a0b0c0b0b0c0b0a0b0a0a0c;
    encBuf[616] = 256'h0a0a0c0b0a0b090909010008080a0d0b0c0c090909080008000909080a0b0a0c;
    encBuf[617] = 256'h0a090b0803020507020303000800090804030705020304020001000001010304;
    encBuf[618] = 256'h020402080a0a0f0b0a0b0a00000102000a080f0b0a0c0a080a09010a0a090d0c;
    encBuf[619] = 256'h090d0b0a0c0c0b0c0b0b0b0b0a0b0a090c0c0a0d0b0a0b0a0008000401010308;
    encBuf[620] = 256'h00000909000a0804000607020404020202000000090002020605030403020302;
    encBuf[621] = 256'h0002020204050304030303040303050203030001080a09000004060303050101;
    encBuf[622] = 256'h0108000800010304040402030302020302040303040304030502020302030208;
    encBuf[623] = 256'h08080b0b0c0c0b090908020304040100080b0b0c0b08020506030201080c0c0d;
    encBuf[624] = 256'h0c0a0b0909090808090801010207030405030404030404020402030203030304;
    encBuf[625] = 256'h0403050203040201020202030305050204020302020203030305040204030204;
    encBuf[626] = 256'h0303050303040302030203030404030502030302030201030402040302040101;
    encBuf[627] = 256'h02020104030205020101000a000909020302050209000c0e0a0b0c0a0a0b090b;
    encBuf[628] = 256'h0e0a0b0d0a0b0c0b0b0d0b0b0c0b0b0c0a0b0b0b0d0b0b0d0b0b0b0d0a0b0b0b;
    encBuf[629] = 256'h0d0b0c0b0b0c0b0a0b0c0b0b0c0b0c0b0b0b0b0b0c0b0b0c0b0b0a0c0a0a0a0b;
    encBuf[630] = 256'h0a0d0a0b0c0b0a0a0908090808090b0c0c0a0c09080801030303040108080a0a;
    encBuf[631] = 256'h0a0b090008020502030502020401030201020300040602060403030502020201;
    encBuf[632] = 256'h02040204040204030204030202030101010909090b09000003060102080b0d0d;
    encBuf[633] = 256'h0c0b0b0a0a080808080b0c0c0c0c0a0c0a0a0b0c0a0b0a0a0908010101000b0e;
    encBuf[634] = 256'h0c0d0b0a0a080303040301080b0f0c0a0c0a090909080909090a0a080a0a090d;
    encBuf[635] = 256'h0c0b0e0a090800030204030008090c0908000306030303010102000307020304;
    encBuf[636] = 256'h0101010900030207050303040201000000010102040202020008010002050202;
    encBuf[637] = 256'h030800010005070504040202020000090a090800020403040302010108080008;
    encBuf[638] = 256'h0003040603040403030402010008090a0c0b0d0a0a0900020404040302020100;
    encBuf[639] = 256'h0103040706040305020303010202010303040503040304030303030303040303;
    encBuf[640] = 256'h0403050204020302030302040103030304030303030203050204040203020101;
    encBuf[641] = 256'h000800020207040304030202000000080001020103000b0b0f0d0b0c0c0a0c0b;
    encBuf[642] = 256'h0b0c0b0b0c0b0b0c0c0b0c0c0b0b0b0b0b0b0a0c0b0c0c0b0b0d0b0a0b0a0b0a;
    encBuf[643] = 256'h0b0b0c0c0b0c0b0c0b0c0b0b0b0b0b0c0a0b0c0b0c0b0b0d0a0b0b0a0a0a0a0a;
    encBuf[644] = 256'h0a0b0b0b0b0c0b0b0b0d0a0c0a0a0b0a090900010002020100080c0b0b0c0804;
    encBuf[645] = 256'h0406050303030203010101040307040304030304030202030202030102030102;
    encBuf[646] = 256'h050205040203030200010900000103060303030201000908000901020801010a;
    encBuf[647] = 256'h0a080d0b0a0f0d0a0c0b0a0c0a090b0c0b0e0c0b0d0a0b0a09090909090b0d0c;
    encBuf[648] = 256'h0b0c0a0b0a0a0a0b0b0c0c0a0a09000808000a0b0b0d0b000105060403030202;
    encBuf[649] = 256'h0000080808010203060403030302020208000101050603040402020101000000;
    encBuf[650] = 256'h0305050404020302020101000203040403030402010101010101010202010101;
    encBuf[651] = 256'h02050403060203010100080809080001020202030303060304020208090c0b0b;
    encBuf[652] = 256'h0a0104050402010a0c0e0b0c0a08000203030304020205040404040303030304;
    encBuf[653] = 256'h0304050402040202020101010203050404030302030202030502030402020401;
    encBuf[654] = 256'h0403030504020303020102000303050504020403010301010201010304020502;
    encBuf[655] = 256'h0204020202030001080909090b000000050208000c0e0b0d0c0a0b0a0a090b09;
    encBuf[656] = 256'h0b0c0a0c0d0a0b0d0a0c0a0b0b0a0a0b0b0b0d0d0b0c0c0b0c0b0a0a0a0b0b0c;
    encBuf[657] = 256'h0b0d0c0b0b0b0c0a0a0a0b0a0b0c0b0c0b0a0b0c0a0b0b0b0b0c0a0a0b0b0b0c;
    encBuf[658] = 256'h0c0b0b0c0b0b0a0b0b0a0b0b0a0b0b0b0d0c0b0d0b0b0a0a0000010402030200;
    encBuf[659] = 256'h0800090005030705030305020202020102010303030405030403030403010202;
    encBuf[660] = 256'h0002020104030403040203030202030204030305040204040203040202020100;
    encBuf[661] = 256'h010800010800010800000909080c0b0a0f0d0b0d0c0a0b0a0908000100090b0f;
    encBuf[662] = 256'h0e0b0b0b09080003020301080a0c0c0b0a0a08020101030000000909090d0b0c;
    encBuf[663] = 256'h0d0c0a0b09090800010808090a0a080903060204050104030405030402020100;
    encBuf[664] = 256'h00080103060503030300090c0b0c0a0102070303030208090b0b090206050404;
    encBuf[665] = 256'h0202010108080800020305040403020202020101010204030503030202010000;
    encBuf[666] = 256'h0900000205030303020000000407050404030402010100010205030603030202;
    encBuf[667] = 256'h0100080001020504030302010808090900030406030202010800080802050405;
    encBuf[668] = 256'h0402040202020202030503050304030302030108000000020403050201000a0d;
    encBuf[669] = 256'h0b0c0b080001030200090d0f0b0b0a0908000201000a0d0d0c0b0a0a08080108;
    encBuf[670] = 256'h080a0e0c0c0c0a0a0a09090a090b0d0c0b0d0b0a0b0b0a0a0b0a0c0c0b0d0b0a;
    encBuf[671] = 256'h0b0a0a09090a0c0b0c0c0b0b0b090a09080a0b0e0c0c0b0b0b0a090808080b0c;
    encBuf[672] = 256'h0d0c0b0c0a090808010100080a0c0c0b0c0908000303040301080a0c0c0a0900;
    encBuf[673] = 256'h0503050402010009090a0909010304040201080a0c0a0b090102040502010108;
    encBuf[674] = 256'h0800010407040304030203010101010304030503030203010200080808090900;
    encBuf[675] = 256'h080104010202090b0a0f0a080901040203030202030305070204030301020909;
    encBuf[676] = 256'h090b0a080800010a0c0d0e0b0c0c0b0b0e0b0c0b0b0b0a090008080a0d0c0c0c;
    encBuf[677] = 256'h0b0a080103040404020100080808080003040405020302020001090800080002;
    encBuf[678] = 256'h0204030203020202040305040204010100080802030705040304030201000000;
    encBuf[679] = 256'h0002040504030402030100010002030306030303020201030206040304040202;
    encBuf[680] = 256'h0101010303050603040304020201020100020304040402030302000009080909;
    encBuf[681] = 256'h01030307040103010808090a0801010604040304020201010201020404020502;
    encBuf[682] = 256'h0203020102020103030003000b090d0e0a0a0b09090b090a0e0a0b0d0a0a0a01;
    encBuf[683] = 256'h010105030204020001080a08090a020302070200000c0f0b0d0b0b0c0a09090a;
    encBuf[684] = 256'h090a0d0b0e0c0a0c0b0a0b0a09090909090b0c0c0c0b0b0c090a090008010108;
    encBuf[685] = 256'h08080c0c0c0c0b0b0c0a0a0a0a090a0b0d0d0c0c0b0c0b0a0b0a090908090a0a;
    encBuf[686] = 256'h0c0b0c0c0a0b0a0a0a0908080800000001090c0b0e0b0b0c0908000203020001;
    encBuf[687] = 256'h0a0d0a0d0b0a0a0a0a0a0a080900040203050108090d0c090900070306030303;
    encBuf[688] = 256'h030100010900000802020303050203040000080b0e0b0e0a0908010305040302;
    encBuf[689] = 256'h02000808000801040405030303040102020201020808080b0c09090802000008;
    encBuf[690] = 256'h0f0e0b0e0b0b0c0a09090a090a0b0b0c0b090908010800010800020002050001;
    encBuf[691] = 256'h010a0900090207020304080b0f0d0b0c0a09000103040101090c0c0c0c0a0908;
    encBuf[692] = 256'h0103040503030402010201000102030605030404020302010000080000000103;
    encBuf[693] = 256'h0304030303030304030302020000080106050505030403030302010101020205;
    encBuf[694] = 256'h040403030402020302020303020303020202030504040404030303020108090b;
    encBuf[695] = 256'h0c0b0a0801060403050200000a0c0b0c0b090002050304020108090b0d0a0b0a;
    encBuf[696] = 256'h09080808000900090901080901090c0a0d0c0808010604040304010208080909;
    encBuf[697] = 256'h0b080908020202040300000a0e0b0e0c0a0c0a0b0a0b0b0b0b0c0b0c0b0c0b0b;
    encBuf[698] = 256'h0c0c0b0c0c0a0a0a090800010008080c0c0d0b0c0b0b0b090a08090a0b0d0d0c;
    encBuf[699] = 256'h0d0b0c0c0b0b0a0b0b0a0b090b0b0d0b0e0a0c0a0a0a0a09080000000008090c;
    encBuf[700] = 256'h0b0d0c0b0b0b09090800010000090c0b0f0b0a0c0a090908010801010800010a;
    encBuf[701] = 256'h0a0a0f0b0a0b0a08080206020204020103000102090002090206020605030404;
    encBuf[702] = 256'h0201020808090a08000104050304040203020101000a0a0a0c09010105060304;
    encBuf[703] = 256'h0302020109090a0b0801030704030403020202010008090a0a0c080102070503;
    encBuf[704] = 256'h030402010809090b0a0a000104060203030100080b0c0b0c0b0a0b0900080202;
    encBuf[705] = 256'h0008090f0b0b0c0a0909000809090a0b0a020606050403030200000908080206;
    encBuf[706] = 256'h050404040202010101000808000001010403050303020301080a0a0d0a090802;
    encBuf[707] = 256'h0504050402030302010200000101040404050304040202020108000000020305;
    encBuf[708] = 256'h0403030502020203020303020203010302020406020503030502010101080800;
    encBuf[709] = 256'h0901030307050304030103010808090b080808040504040302020208080a0c09;
    encBuf[710] = 256'h0a0a010202070402040200000a0c0b0c0b0a0808040203040108090b0e0a0b0b;
    encBuf[711] = 256'h0a090902010004010000090e0b0c0d0a0a0a080801010108090d0d0a0c0a0a08;
    encBuf[712] = 256'h0908080a0a0d0c0c0b0b0a0a0a090b0c0b0d0c0b0c0c0a0b0b0a0a0a09080800;
    encBuf[713] = 256'h0a0c0c0d0c0b0c0b09090001010101090a0c0e0c0b0b0c0a090908080800090a;
    encBuf[714] = 256'h0c0e0c0b0d0b0b0b0a09090908090a0b0e0c0b0c0a0b0a0a0908080808080808;
    encBuf[715] = 256'h090a0b0b0e0b0b0b0c0a090900080101000a0c0f0d0b0c0b0b0a090102020501;
    encBuf[716] = 256'h00000b0c0b0d0a09090003020305020203000102080000090005020705030305;
    encBuf[717] = 256'h02010108090a0b090800020602040302020109090a0c0a080903070304040101;
    encBuf[718] = 256'h00090a0b0d0a080801030202020808090c09090a0a080b0a0009020703050301;
    encBuf[719] = 256'h090a0f0b0c0a09010206030302010a0c0b0d0a0800020404030201080a0c0c0b;
    encBuf[720] = 256'h0b0a0001030602030108090b0e0b0a0900020504050203020100000908010103;
    encBuf[721] = 256'h0704040303030202000808080001040503050302020000080809080102040603;
    encBuf[722] = 256'h0403030302020301020404040504030303030201010101020405030402020100;
    encBuf[723] = 256'h09090908010204030202000909090a0801000303000301040704040502020101;
    encBuf[724] = 256'h0900080005040404030102080a0a0c0c0a0a0a080800000109090d0e0c0c0c0b;
    encBuf[725] = 256'h0a0a000003040201000c0d0c0c0b0a090802010302000a0c0d0c0b0c0a090808;
    encBuf[726] = 256'h0008000009090c0c0c0b0c0a0b0909080800080a0b0d0c0c0b0a0a0908080909;
    encBuf[727] = 256'h0b0d0c0b0c0b0b0a0b090a0b0b0d0d0b0c0c0b0c0b0a0a0900010001080b0d0e;
    encBuf[728] = 256'h0c0a0b0a09000102030202090c0b0f0c0a0b0a0a08000102030400080b0f0c0b;
    encBuf[729] = 256'h0d0a0909000101020308090a0e0b0b0c0a08090102030305020102090a0c0c0b;
    encBuf[730] = 256'h0a09000303050301090a0f0b0a0b0801000203080a0b0f0a0800020702030201;
    encBuf[731] = 256'h08090b0900010604040303020202010304020303010203020506040305020201;
    encBuf[732] = 256'h0009090a08010205050203030302020002020102030306050404040303030100;
    encBuf[733] = 256'h090b0a08000505040402010108090a0808020404040303020201010102030304;
    encBuf[734] = 256'h0403030403050302020200080808020505040403030100090809000305050502;
    encBuf[735] = 256'h0302020101000202020503030503030404020303020301000101010405030503;
    encBuf[736] = 256'h0202010800000a00080901010006030404030202000a080a0b01040507030203;
    encBuf[737] = 256'h020000080a08080903010002000a020208070009090d0e0a0b0a080008040009;
    encBuf[738] = 256'h080c0d0a0b0b08080901090d090a0c000100040108080b0f0a09090201000309;
    encBuf[739] = 256'h0e0b0d0c09090900000a0a0d0e0a0b0a090808000009090b0e0a090a00080802;
    encBuf[740] = 256'h080a00000007040204000a0a0e0b0a090003050202000c0b0e0c090a08080108;
    encBuf[741] = 256'h000a0b0c0c0b09080900090c0c0c0c0a0a0900000000090b0c0d0c0b0b0b0a0c;
    encBuf[742] = 256'h0b0c0b0c0a0b0a0a0c0b0c0e0b0c0b0b0a0a09090808090b0b0d0c0a0b0c0b0b;
    encBuf[743] = 256'h0c0c0a0b0a090900090a0d0d0d0c0b0c0a0a09080008080a0b0c0d0b0c0b0b0a;
    encBuf[744] = 256'h0a0a090909000809080a0b0b0d0c0a0909010203060203020008080a0c0a0c0b;
    encBuf[745] = 256'h0b0b0b080800050100000e0c0b0e0a090a080101020300010209080108010508;
    encBuf[746] = 256'h01020a01050106040203030000080b09080b08020a08000d0902000407010201;
    encBuf[747] = 256'h090b0b0e09010307070304030302020201020203050304050204020203010008;
    encBuf[748] = 256'h090b0a090a000202040201090c0e0b0c0b0a08080202030101090a0b0c090800;
    encBuf[749] = 256'h0307030403040302020100090908000407040305020100090b0d0b0a08000405;
    encBuf[750] = 256'h030403020101080800000205040404030402030203010008090a090a08010205;
    encBuf[751] = 256'h04020200090c0c0d0b0b0a090000020203030402010100080808000405060403;
    encBuf[752] = 256'h04040202020102010001010808090a0b0a090003040402090d0e0d0c0b0b0a09;
    encBuf[753] = 256'h000103040202020008090a0b0b0c0a090002060403040200090d0d0c0b0c0b0a;
    encBuf[754] = 256'h09000000010108090b0d0c0b0c0a0a0908020305030403020000090908000204;
    encBuf[755] = 256'h06030502020101010808080a0a0b0d0d0b0c0c0a0b0a0b0a0c0c0b0c0b0b0c0a;
    encBuf[756] = 256'h0b0a0a0b0a090801030404040201000a0a0b0b0901060505030303010108090b;
    encBuf[757] = 256'h0b0b0b090002050503040201080b0e0c0b0b0a0801030404030100090b0b0b0b;
    encBuf[758] = 256'h090001020300080a0f0b0c0d0b0b0d0b0b0c0b0b0a0b0a0c0b0c0b0c0a090800;
    encBuf[759] = 256'h0203040101000a08080105050504040303030303030202000008000003060504;
    encBuf[760] = 256'h04030200090b0f0b0b0b0a0001030503020208090c0c0b0c0909010204040402;
    encBuf[761] = 256'h03020000090a0a0b0900010306030402030202000008090c0b0d0b0908020605;
    encBuf[762] = 256'h0403030202080a0a0b0a00030705040303030302010100000000000102030306;
    encBuf[763] = 256'h0303040202000a0b0d0c0c0a0b090800040404040303020100090a0a08010407;
    encBuf[764] = 256'h050403040203010008080a0909080104050305020200080a0c0d0a0b0a090801;
    encBuf[765] = 256'h02030101080b0d0c0c0a0a0901010203040101010801000002020101080b0b0e;
    encBuf[766] = 256'h0c09090901030204020a0b0f0e0b0b0c09090002030404020200080b0a0d0b09;
    encBuf[767] = 256'h08080305040403030300080a0d0d0b0c0b090908010001000a0d0d0d0b0c0a0b;
    encBuf[768] = 256'h090900000100010009080a0b090a09020202060201020102030203040109090e;
    encBuf[769] = 256'h0e0b0d0b0b0a0a08000001080b0e0d0c0c0b0b0a0a090800020202010208080b;
    encBuf[770] = 256'h0c0c0b0b0b080003070403040101090b0f0b0d0b0a0b09080001010108090e0c;
    encBuf[771] = 256'h0c0b0c0a0a0900010103030200080a0c0c0b0b0a09000102020301080a0e0d0c;
    encBuf[772] = 256'h0b0b0d0a0a0a0a0a0b0b0c0c0b0c0b090a0a09090a0b0c0c0a0a090004040604;
    encBuf[773] = 256'h0303030201010809080800030704040303030201090a0c0c0b0a090002040503;
    encBuf[774] = 256'h040101080a0b0e0b0b0b0a00010405030302000a0b0f0b0c0a0a080002040203;
    encBuf[775] = 256'h02000a0c0c0d0a0b0909000203050303020000090a0a0a000204060403030302;
    encBuf[776] = 256'h01010808080808010800000a0a080a09030102030e0d0d0f0b0b0d0b0a0a0800;
    encBuf[777] = 256'h00010208090c0e0c0b0d0a090900010302030200080b0d0b0b0b090802050403;
    encBuf[778] = 256'h05030203010100090a090a0003060605030304010100090a0a0a090801040503;
    encBuf[779] = 256'h030501010008090a0a0b0909010204060304040202020000090b0b0c0a090005;
    encBuf[780] = 256'h05040502020208090c0c0b0a0a000205050303030200090b0b0d0a0908020306;
    encBuf[781] = 256'h040303030200080a0b0e0a0a090802040404020200090b0d0c0c0b0a0a090001;
    encBuf[782] = 256'h02020202080a0d0c0c0c0a09090002030404030202010008090a0b0a09000206;
    encBuf[783] = 256'h05040403030200090b0d0c0a0a09000203040202080b0d0d0b0b0a0a08000101;
    encBuf[784] = 256'h010108080a0b0a09090000090a0d0d0d0b0c0a08000203050202090b0f0c0b0b;
    encBuf[785] = 256'h0a08010306030402020008090909090001020404040404030304020100090b0c;
    encBuf[786] = 256'h0c0b0908010306030201080b0f0b0d0b0a0b090800010203020100090c0c0c0b;
    encBuf[787] = 256'h0b0b0900030405040302020100090b0c0c0b0a09010306040403020200090b0c;
    encBuf[788] = 256'h0b0b0a08010405040303020200000a0a0c0b0b0b0a0003060504030301000a0c;
    encBuf[789] = 256'h0d0c0b0b0a09000103030301080b0d0d0c0b0b0a080801030306020303010101;
    encBuf[790] = 256'h0809090a0900000307050404030402020100090c0b0b0a090104060305020200;
    encBuf[791] = 256'h090a0d0b0c0b0a090001030305020200090b0d0c0b0b0a090003050403030201;
    encBuf[792] = 256'h090a0c0c0b0c0909000204040403020201000a0b0d0b0a090002050503030301;
    encBuf[793] = 256'h00090b0d0b0b0a0800020404040303020100090b0c0c0b0a0a08020306030302;
    encBuf[794] = 256'h00090c0c0d0a0b0a09080102040403020101090a0c0c0b0a0908020403040202;
    encBuf[795] = 256'h010009080808080009000808030505060303040100090b0d0b0c0b0908090100;
    encBuf[796] = 256'h01010201010108090c0f0c0b0b0b0900040503040301010a0c0d0c0b0b0a0a08;
    encBuf[797] = 256'h00020404020301090a0e0c0b0b0b090002050304020200080a0b0d0c0b0a0a08;
    encBuf[798] = 256'h0002050404020300080a0d0c0b0b0a08000203030300090c0d0c0b0c0a0b090a;
    encBuf[799] = 256'h09090002030405030202000a0b0c0c0b09000306040304030200090a0c0d0b0b;
    encBuf[800] = 256'h0a08000204030302080b0e0c0c0b0c090a09080808080808000800080a0d0c0d;
    encBuf[801] = 256'h0b0b090801040504020201080b0b0d0b0a09000204040302030100080a0a0a0a;
    encBuf[802] = 256'h0908020405040303030302000008090a0c0b0b0b0908030706030302000a0d0d;
    encBuf[803] = 256'h0c0b0b09090102030201080b0e0c0a0a09080102030202020001000000000000;
    encBuf[804] = 256'h0001000002040101010000010107050305030101080a0a0b0b08000304040100;
    encBuf[805] = 256'h000b0b090a09080a080a0c0a00020507030302010a0d0d0c0c0b0b0b0b0a090a;
    encBuf[806] = 256'h08080908090b0e0d0c0c0b0b0900020405020200080b0d0c0a0a090001030403;
    encBuf[807] = 256'h0201010808000101030403040303040202030201020008090c0e0c0d0c0b0b0a;
    encBuf[808] = 256'h090001040302020a0c0e0c0b0a0a00020404030201000b0c0c0b0b0909010203;
    encBuf[809] = 256'h05030304030202010008000800030405040201010a0d0b0e0c0a0c0a090a0808;
    encBuf[810] = 256'h0801010000080a0c0b0d0a090802040303020a0d0e0c0b0a0b08010104030202;
    encBuf[811] = 256'h00080a090a010304060402020208090b0d0c0a0b0b090b0908090a00090a0101;
    encBuf[812] = 256'h04060304020109090d0b0a0a0004030304080a0f0e0b0b0b0a00020504030402;
    encBuf[813] = 256'h0108090b0b0b0a080304050403020100090a0d0b0a0a08020404050203030100;
    encBuf[814] = 256'h0808090809000202040502020302020202020302020303070403050403040303;
    encBuf[815] = 256'h04010101000a090909090800030403040201090b0f0c0b0c0b09000203060303;
    encBuf[816] = 256'h030201080a0b0a0a000306060404020303010100080900000105030603030303;
    encBuf[817] = 256'h0100080a0a0b09080101040302020108090b0b09000007030205020102000801;
    encBuf[818] = 256'h0800030604050302030109090b0b08020407050304020100080a0a0b0a080003;
    encBuf[819] = 256'h050402030200080a0d0a0a0a08030307040203020001080b09090a0001010301;
    encBuf[820] = 256'h0801080b05040406030303030008090b09000007040305020101090c0c0b0c0a;
    encBuf[821] = 256'h090803040405020201000a0a0c0c090a0801020205010009090d0b0c0b090909;
    encBuf[822] = 256'h01020305040203030000080a0b0b0b09000206030302010b0b0d0d0a0a0a0802;
    encBuf[823] = 256'h0103030103030900080a08000c0a0d0e0a0c0d0a0a0b08010004030201080c0b;
    encBuf[824] = 256'h0e0b090800050403030200090c0d0b0b0b090801020208080b0c0c0b0b080002;
    encBuf[825] = 256'h0404020300080a0b0d0808010405030302090b0f0d0b0b0b0a00030504040201;
    encBuf[826] = 256'h08090b0d0b0b0b08010304040301000b0c0e0c0b0a0b08000103050302010009;
    encBuf[827] = 256'h0b0d0b0a0900010305020101090a0b0d0b0c0a0a0a090a080801000203060202;
    encBuf[828] = 256'h00090d0c0c0b0c0a09080800020000090b0f0d0c0a0b0a08080101030201080a;
    encBuf[829] = 256'h0d0d0c0b0a0b0a0a0a09090b0a090a0b0a0b0d0d0b0c0b0a0900010404030201;
    encBuf[830] = 256'h08090b0d0b0b0a090808000008090a0b080a0a090a0d0b0d0b0b0c0b08080800;
    encBuf[831] = 256'h0108090c0d0c0c0d0b0a0b090000010301010a0e0c0c0b0b0a0801020102000a;
    encBuf[832] = 256'h0b0f0c0a09090101020400080a0b0e0b0b0901020504020202090c0c0c0b0a0b;
    encBuf[833] = 256'h09020204040200090d0c0c0c0a0a090801010202080a0b0f0b0c0b0a08090001;
    encBuf[834] = 256'h0008010909090b0b090909000000010b0a090c0b0a0c0a090a0a010a0b080d0b;
    encBuf[835] = 256'h0a0c0a01000205020203080b090f0a0b0c0a080b0a090a09010908010b0b0b0f;
    encBuf[836] = 256'h0b080a090002050502020308080a0d0b0b0b0900080205020404000102080800;
    encBuf[837] = 256'h0900020106050204030202000808090b0b090a08030204070203040302030202;
    encBuf[838] = 256'h0200090201030703040503020108080a0d0c0a0a0a0800020504030302020009;
    encBuf[839] = 256'h0c0b0b0b00030607030304020108090a0b0b0908010505040304020202000808;
    encBuf[840] = 256'h090000020504040303020100090a0a0a0a080104040303030303020405040402;
    encBuf[841] = 256'h030301000009090808020403030301080c0d0d0a0a0900020604040402020201;
    encBuf[842] = 256'h08080808000104040402020100080a0908010604050303040201000808010000;
    encBuf[843] = 256'h030503030201080c0d0b0c0c0909000104050303020208090a0b0b0802040604;
    encBuf[844] = 256'h03020108090b0d0a0b0a08080002020202000000080802030106010100090b09;
    encBuf[845] = 256'h0d0b000205060403040100090b0c0a09000406040403020200090a0b0d090908;
    encBuf[846] = 256'h02030404030100080a0b0d0b0a090902040403040301000909090b0b09090008;
    encBuf[847] = 256'h09090a0d0a0b0b08090a00090f0b0d0c0a0a090203060403020200090a0d0d0a;
    encBuf[848] = 256'h0a09000104040403030100090c0b0c0b0901020504030302000a0c0c0d0a0b09;
    encBuf[849] = 256'h090800020102010100090b0e0b0b0d090908000103030201000a0d0d0c0b0c0a;
    encBuf[850] = 256'h09080801030403040200000b0d0c0b0a0a08000203040200090a0d0c0a0a0900;
    encBuf[851] = 256'h010204010102010800080a000a0b0b0e0b0a0c0a080900010008020201010000;
    encBuf[852] = 256'h000c0a0b0e0a0b090a090a0a0c0d0c0a0d0a0a0a090a080908090a0900020101;
    encBuf[853] = 256'h0801080b0b0c0d0c0a0b090b09080802040404040201080b0e0c0b0b09010405;
    encBuf[854] = 256'h040202000a0c0d0c0c0a0a0900020303040300090b0e0b0c0b0a080002030503;
    encBuf[855] = 256'h0200090c0c0c0b0b0a09080102020201010808090a0a0b0c0b0b0c0a08020604;
    encBuf[856] = 256'h04040201080a0d0d0b0b0b0b080102040404020200090c0d0b0b0a0908020403;
    encBuf[857] = 256'h040201080b0e0c0b0b0a09000103040303030202010008090a090b0b08010106;
    encBuf[858] = 256'h03030200090d0f0c0b0b0c0b0a080003050403030301080a0d0d0a0b09080103;
    encBuf[859] = 256'h05030301000a0c0c0b09090104040404020201000009090a0909090008000808;
    encBuf[860] = 256'h0a0a0d0a0a0a01020307040202010808080a00040405030301000a0c0d0b0a0a;
    encBuf[861] = 256'h0a0808080101000203020402010201090b0a0c0a090803060304030000000a0a;
    encBuf[862] = 256'h090d0b0b0b00010207070303030201090b0c0b0d09090001040403040101000a;
    encBuf[863] = 256'h0b0e0b0c0a0a080205040403030208090c0c0b0b0a0001030603020101090a0c;
    encBuf[864] = 256'h0c0b0b090900010204040202030108000b0d0b0c0b0a08000104040403040202;
    encBuf[865] = 256'h00090c0d0b0b0a0802070403040201000a0b0c0c0b090802030503040100080a;
    encBuf[866] = 256'h0b0b0c0a090801020304030201080a0d0b0c0a09090102030302020100010202;
    encBuf[867] = 256'h030301080c0d0c0b0c090802040404020008090b0c0a09000101030201030301;
    encBuf[868] = 256'h01080a0c0e0b0b0b0909010305030202020009000204030303010c0e0c0c0b0a;
    encBuf[869] = 256'h080003030401080a0d0d0b0b0a09080103050404020201080b0d0c0c0a0a0a00;
    encBuf[870] = 256'h000303040201090c0c0b0c0a090800010001010202030403080a0f0e0b0c0b0a;
    encBuf[871] = 256'h090002050303030201090b0d0b0c0a09000105030504020201080a0d0c0c0a0a;
    encBuf[872] = 256'h080102040402010109090b0c0b0a0a080103050403030201090b0e0b0c0a0a08;
    encBuf[873] = 256'h0001050203010008090a09080003040301000a080808040403050201090c0c0c;
    encBuf[874] = 256'h0b0b00010405050304020101000809090a0a0801040504030202090a0c0d0a09;
    encBuf[875] = 256'h0801040304020201080000000103020201090d0c0b0c0908030403030208090c;
    encBuf[876] = 256'h0c0a0a010205040303030201010a0b0b0e0c0a0800020304040108080a0a0004;
    encBuf[877] = 256'h04060402010109090b0c09010305040302000a0c0d0c09090001020304030000;
    encBuf[878] = 256'h000a090b0c0b090a00030306040201080a0b0d0c090a08010303030301090d0b;
    encBuf[879] = 256'h0a080205040101000a0a0a0a01010305030103010908090b0a0c0d0a0a090101;
    encBuf[880] = 256'h0505040202080a0c0d0c0a090800020404010108090b0a0b0c09090901020205;
    encBuf[881] = 256'h0502030100080b0d0c0b0b0a000103040202010a0c0a0c0b090b0b0a0b0c0909;
    encBuf[882] = 256'h080103050108090c0f0c0a0b0b080000030304020100090c0c0c0b0c0b090908;
    encBuf[883] = 256'h0304040201080a0e0d0a0b0908010305020201080a0b0c0a0a09010100010008;
    encBuf[884] = 256'h0d0b0a090a08030306030100080a0c0c0c0a08080102030400090e0d0d0b0b0a;
    encBuf[885] = 256'h08000404030302080a0c0c0a0b08000303050200090c0c0a0c0a080001020203;
    encBuf[886] = 256'h010008090909080801060203040200080c0d0c09090901030404020100090b0c;
    encBuf[887] = 256'h0b080802050502030108080b0d0b0a0b0a080901000002010a090a0a0b0b0908;
    encBuf[888] = 256'h08030403030301090b0c0a090a0803040302000a0b0b0e0b0a00010305040303;
    encBuf[889] = 256'h0101090a0b0d0b0a0001050503030301090b0f0c0a0a09000203050402020009;
    encBuf[890] = 256'h090a0b0a0801030403030109090b0b0b0a0a0000000001080a080b0901030406;
    encBuf[891] = 256'h03040302080a0c0d0c0a0a0900020404020200090c0c0b0b0b08020603050302;
    encBuf[892] = 256'h0101090b0c0c0a0a0900010304030201000a0a0d0b0a09090204030404000008;
    encBuf[893] = 256'h090c0a0b0c0b0a090909080909080100000908080b0b0a0a090a0909080a0a09;
    encBuf[894] = 256'h0c0c0b0b0c0a0b0908090a01000a0a0908080000020002020009090b0c0b0c0a;
    encBuf[895] = 256'h090801030202020a0a090d0b0a0a09000101080100090b0c0a0b0c0a08090b0a;
    encBuf[896] = 256'h09090a090108000102000808080a0d0a090a09010204040101000a0c0b0c0a0a;
    encBuf[897] = 256'h0a08020204030403020908090a0b0a0b0001000305030402020201090a0b0b0b;
    encBuf[898] = 256'h0b09030703030503020009090a0b0c090802050303050100080b0c0b0b090003;
    encBuf[899] = 256'h06040303020008090b0a0808050503030301000a0c0c0b0a0002040603040201;
    encBuf[900] = 256'h00080a0a080801040405040201010009090a0b08000003060303030201030203;
    encBuf[901] = 256'h030504010202080908090b000202040404020009090b0e0a0a08030604050302;
    encBuf[902] = 256'h020108090c0a0b0a08000404040303020009090b0d0a09000205040403040101;
    encBuf[903] = 256'h0009090a0a0b080001030703030402010009080a0b0801020704030403010100;
    encBuf[904] = 256'h0a0a0a0b0a080005030405020001090909090a010203070302020100080a0a09;
    encBuf[905] = 256'h090103020306010001080a08090b01020003030103020902000a010008010008;
    encBuf[906] = 256'h02010902010804010802020a08090d00080a02010105020103000b00090e0909;
    encBuf[907] = 256'h09080000040101030008090c0c0a0c0b090a0a010303040201020a0d0b0f0b0b;
    encBuf[908] = 256'h0a0a00010207020101080c0b0c0c0b0a09010203060201010a0b0c0d0b0b0909;
    encBuf[909] = 256'h020204030208000a0f0b0b0b0a090801010202000b0c0e0b0b0b0b0908000100;
    encBuf[910] = 256'h00000a0c0b0c0b0a0b0a090b0b0c0d0b0b0d0b0a0a0a09090a0b0c0a0b0c0d0a;
    encBuf[911] = 256'h090a090a090c0d0b0b0d0c0a0b0a0808090a0a0a0c0d0a0c0a09000101020202;
    encBuf[912] = 256'h080b0e0c0c0b0a0b0a09000108000a0b0d0c0c0a0b0a0900080103000901090c;
    encBuf[913] = 256'h0c0c0b0b0d0b0b0b0c0b0a09090908000a0a0b0c0b0c0c0b0a08000103010200;
    encBuf[914] = 256'h0a0b0e0d0a0b0b0a0908020202040100000b0b0b0b0a080a0003010103090101;
    encBuf[915] = 256'h090d090b0c090c0a080908020802040100080b0b0b0c0a090002050203030009;
    encBuf[916] = 256'h090c0d0b0a0900080106010801090b0c0a0c0809020401030309090a0d0b0b0b;
    encBuf[917] = 256'h08010002030000080c0b0a0b0b080103050304020101080900000a0002000100;
    encBuf[918] = 256'h0901010908010a08020908000900000802050203040102000b0b0a0e0a080901;
    encBuf[919] = 256'h030205020800090f0a090a0001020504030201080a0a0c0b0900020603030303;
    encBuf[920] = 256'h00080b0d090a0803050504020201080a0a0b0a000003070304030100080a0b0a;
    encBuf[921] = 256'h0a080304070303010209090a0b0b000005040404020101010809090003040405;
    encBuf[922] = 256'h02020200090b0b0b08010204060202030109090a0a090002070403030300080a;
    encBuf[923] = 256'h0d0b0a0b08000306040203010000090a09080307030603020302000809090b09;
    encBuf[924] = 256'h0002020603040202010009080901050304040403010108080a0b0a0a01000303;
    encBuf[925] = 256'h0201000b0c0b0b0b08040504030503010208090a0a0a0002040504040201080a;
    encBuf[926] = 256'h0a0c0a0a000206040403030200080a0a0a0a0003060503030201080a0c0b0a0a;
    encBuf[927] = 256'h08040404040302010009090b09010106050304020201080a090a0a0002040603;
    encBuf[928] = 256'h03030200000a0b09010206050403040102000808090a00010105040203020001;
    encBuf[929] = 256'h0809000108050503050303040302020201030303060201030401020202030302;
    encBuf[930] = 256'h0503000404010404020304020401010200080100000201010701080101080001;
    encBuf[931] = 256'h0806040206030204030101020001020004040204030103020801080803050206;
    encBuf[932] = 256'h040205020002010801000902030105020103010a010a0e000009050301060200;
    encBuf[933] = 256'h020009000009030402060301030109080a0e00080805030305020001090c090a;
    encBuf[934] = 256'h0c08010005020103020d0a0b0e0a0a0a01010004030801090e0a0c0b0a090902;
    encBuf[935] = 256'h030105010a080a0e0a090b00010004020101090d0a0c0d090909000008010a0e;
    encBuf[936] = 256'h0a0c0c0a0a0a00000802080a0a0e0e0a0c0b090908000108000b0d0c0d0b0b0b;
    encBuf[937] = 256'h09080101030300080c0f0b0c0b0a0a0801020201000c0c0d0d0b0b0a09080002;
    encBuf[938] = 256'h0201000a0e0c0c0b0c0a080800000100090b0d0d0b0c0b0a090800000100090a;
    encBuf[939] = 256'h0d0c0c0b0a0a0a08000808080a0c0d0c0c0a0b0b090a09090a0a0c0d0c0b0b0b;
    encBuf[940] = 256'h0b0b0b090b0b0b0e0c0b0d0b0a0a0b090a090a0b0d0b0e0b0b0b0c090a080809;
    encBuf[941] = 256'h09080c0c0b0d0b0b0a0a090908000a0b0c0f0b0c0b0c0a0a0a08090a080b0c0a;
    encBuf[942] = 256'h0e0b0a0b0b090b0a090a0a0a0f0b0a0c0c0a0b0b0a0c0a090c0a090a0b080b0a;
    encBuf[943] = 256'h080c0b090e0a090c0a000b09080b0c0a0f0b0a0d0b090a09000900030a0a080f;
    encBuf[944] = 256'h0b090d0a080908020800010b0e090f0a090b09080801030000030b0b0a0f0b08;
    encBuf[945] = 256'h0b08040002050808000d0b090d0a080a00020102030809000f0b080b09020802;
    encBuf[946] = 256'h060001020b0b090e0a080a08040003050800020a0a010a000501030701010208;
    encBuf[947] = 256'h08000a08030803070302050000010a08010902070102050101020808010a0004;
    encBuf[948] = 256'h0004050203040001020900020902050304050202040001010000030105040303;
    encBuf[949] = 256'h0502020301010300010402040502030402020301020301040402040502030303;
    encBuf[950] = 256'h0304010203020305020404010304020303020403020403030503020403020403;
    encBuf[951] = 256'h0203040203030303040305030304030403030303030304030403050304030303;
    encBuf[952] = 256'h0402020202030205040304030403030302030203030305050204040203020302;
    encBuf[953] = 256'h0201030202050403050402020301020208020102040404040303030301020108;
    encBuf[954] = 256'h0204020604020403020301000000080303030705020302010201080101000503;
    encBuf[955] = 256'h0405030203020001080902010106040204030202020901000903040207030204;
    encBuf[956] = 256'h020101010900000a03030207040103020001000b010809050302070301030209;
    encBuf[957] = 256'h00090c08080a05020205030002080b090c0c000008050301050109010a0d0909;
    encBuf[958] = 256'h0b00010004020002000e080b0d08090901010804010a000a0e090a0c00090902;
    encBuf[959] = 256'h080a010a0e090a0e08090b00090b010a0d080a0d09090c08090b080a0d080a0d;
    encBuf[960] = 256'h09090c08090c08090c080b0b090b0d08090b080a0e080b0c090a0c08090b0809;
    encBuf[961] = 256'h0c090c0d0a0a0d09090a000909000a0c0b0c0d0a0b0c080909000009090b0f0b;
    encBuf[962] = 256'h0c0c0a0a0b0808000108090a0d0d0c0b0b0b0a0900000002090b0e0d0c0b0c0a;
    encBuf[963] = 256'h090908000000000a0c0c0c0d0a0a0a090008010008090c0d0b0c0c0a0a0a0808;
    encBuf[964] = 256'h000000090a0d0c0c0b0c0a090a08000000080a0b0e0c0c0b0b0a0a0900000000;
    encBuf[965] = 256'h090b0e0c0c0c0a0b0a090800000108090c0d0c0b0c0b0a0908000000010a0b0e;
    encBuf[966] = 256'h0d0b0b0c0a090808010000080c0b0d0c0b0a0b0a08080000080a0b0e0d0a0c0a;
    encBuf[967] = 256'h0a0a09080809080a0c0a0d0b0a0c0b080b09080b0b0a0f0b0a0c0a0a0b0b090b;
    encBuf[968] = 256'h0b0a0e0b090d0a090c09080a09080b0b0b0f0b0a0c0b090a0a000b09000d0b0a;
    encBuf[969] = 256'h0e0b0a0c0a000a00020908000d0b0b0f0b090b09010900040908000d0b0a0e0a;
    encBuf[970] = 256'h08090802080102090a080f0a090b0a000900040800020c0a000d09010a08040a;
    encBuf[971] = 256'h08030c0a010d09020901070000030909000d09000902060102050000010b0b08;
    encBuf[972] = 256'h0e09010003070103030000010b0a090b00040206050201030808080c0a080900;
    encBuf[973] = 256'h050204050102020000080a08010802060204030201020908010b080301040702;
    encBuf[974] = 256'h0205010203000203000304010104000204000305020304010302000203000307;
    encBuf[975] = 256'h0305040303040102010808010802040306040202030201010000020205050304;
    encBuf[976] = 256'h0402020201010100010203050402040302020201030204040403050203020101;
    encBuf[977] = 256'h01010103050306030304020100000808010205050404030202010009090a0900;
    encBuf[978] = 256'h030704040402020000090a0a0908010505040402020108090a0b0b0900020605;
    encBuf[979] = 256'h0304020101090a0a0b0a080105050403030200080a0c0a0b0a00030505040202;
    encBuf[980] = 256'h0100080a0b0b09090205040503010200080a0a0c0a080803050305030102000a;
    encBuf[981] = 256'h090a0a09000205050204010101090a090a0900010307030203020000080a0808;
    encBuf[982] = 256'h0804030306020102080908090a02020207040003010900090b01000907020103;
    encBuf[983] = 256'h0208000a0f080a0a020101070201020109080a0d090a0a01010006020002080c;
    encBuf[984] = 256'h080b0e09080901020206020102000b090c0d0a090b00010804010002080d090b;
    encBuf[985] = 256'h0e08090902030106020001080c0a0b0f09090a08000802020801090c0a0c0c09;
    encBuf[986] = 256'h090a02020206020000090e0a0d0b0b0a0b000008030208010a0f0a0b0e090909;
    encBuf[987] = 256'h010101040108080b0f0b0c0c090a0a000100020108000c0d0b0c0b0b09090102;
    encBuf[988] = 256'h0203020a0b0f0f0a0b0c09090901010101010a0a0e0c0b0c0a09090002020102;
    encBuf[989] = 256'h080c0c0d0c0b0b0a090801020101010a0d0d0c0b0b0b09080001030108090c0e;
    encBuf[990] = 256'h0b0d0b0a09090000000100090b0d0d0b0b0c0a090908080008090b0c0c0c0b0b;
    encBuf[991] = 256'h0c0a0a0908090a090c0b0d0b0c0c0a0b0b0b0a0b0b0a0b0c0b0c0c0b0b0c0a0b;
    encBuf[992] = 256'h0c0a0b0b0b0d0b0b0d0b0b0c0b0b0b0c0a0b0b0b0d0b0a0b0c0a0a0b0a0c0b0b;
    encBuf[993] = 256'h0c0c0b0d0b0a0c0b090b0b090b0b0a0d0b0a0d0b0b0c0a090b09080a09090d0c;
    encBuf[994] = 256'h0a0e0b0a0c0b090909000800010b0b0b0f0d0a0a0b080900020000020a0d0a0f;
    encBuf[995] = 256'h0b0b0b0a08080004020103090b0a0f0d090b09000801030102030a0c0a0f0a0a;
    encBuf[996] = 256'h0a0a0100030501020309090a0f0b090b09010802040102030a0a090f0a090a08;
    encBuf[997] = 256'h030003070101020a08080c0a080b080208010608010309000309010600010408;
    encBuf[998] = 256'h01030901050002070002020800020b09000a02070205050202030001010a0901;
    encBuf[999] = 256'h0902060205040203020108000a0a010a01070304060202020100010a09000901;
    encBuf[1000] = 256'h040306040303030001000b09090a010504040503030301000009090809000602;
    encBuf[1001] = 256'h0504020303010000090909080104040504020304000101080800080104030504;
    encBuf[1002] = 256'h0203030201010900000802050305040303030302020001020304050305030203;
    encBuf[1003] = 256'h0302020202030403060203040202020302040305030403040202020101010103;
    encBuf[1004] = 256'h0503060303040202010100000001030604040304020202000008000800030504;
    encBuf[1005] = 256'h0404030302010100090908080205040503040202010000090909080205030603;
    encBuf[1006] = 256'h0304020000080a08090902030406040202020100000908080802050305040203;
    encBuf[1007] = 256'h0200010009080009020303070501030201020108020101030501050301040200;
    encBuf[1008] = 256'h03010003020104030004020005020106030204040003010801080b0102000704;
    encBuf[1009] = 256'h0105020002000a08090b01020107050204020000000a090a0a00010107030204;
    encBuf[1010] = 256'h020001080a080a0a01030107040104010001080908090b010009050201050300;
    encBuf[1011] = 256'h03020a03080d01090b01010a07010004010902080d080a0c08080a0303000703;
    encBuf[1012] = 256'h0002000b080b0f0a090c00000804020003010a080c0f090a0b00000805020104;
    encBuf[1013] = 256'h0109090b0f0a0a0b090800030303050109080c0e090b0b08080803030104000a;
    encBuf[1014] = 256'h0a0e0d0a0b0c09080801010003000b090d0d0a0c0b09090a00000900080c090c;
    encBuf[1015] = 256'h0d0a0b0d090a0a08090a08090b090b0f090c0b0b0c0c0a0a0b09090a08090c09;
    encBuf[1016] = 256'h0b0d0b0d0c0a0b0b090a0a08090b0a0d0d0a0d0b0b0c0a0a0a09080909080a0d;
    encBuf[1017] = 256'h0a0d0c0a0c0b0a0b0a090a09080a0b0c0d0c0c0b0c0a0b0a0908080008080a0c;
    encBuf[1018] = 256'h0e0c0c0b0b0b0b0a0908000808090d0c0c0c0c0a0b0a090800000008090c0b0f;
    encBuf[1019] = 256'h0c0a0b0b0b090908000800090b0c0e0c0b0b0c0a0909080008010a0a0c0e0b0c;
    encBuf[1020] = 256'h0c0a0a0a090008000009090b0e0b0c0c0a0a0a09000908000a0b0b0f0c0a0b0b;
    encBuf[1021] = 256'h090b09080909080b0b0b0f0b0a0d0a090b0a090c0a090c0a090c0a090b0b090d;
    encBuf[1022] = 256'h0b0a0d0a090b0b000b09010c0a090f0b0a0d0a090a09000800020908080f0b09;
    encBuf[1023] = 256'h0d0a090a08020800040908000e0b090d0a090a08020802040900010d0b090e0a;
    encBuf[1024] = 256'h080a09020908040808020b0a010f0a000c09010900040802040800020c0a080e;
    encBuf[1025] = 256'h09000a01040103060101020909000d09000901060103050102010809000c0900;
    encBuf[1026] = 256'h0802060204040102020808000a09010802070203060101020900000a08010804;
    encBuf[1027] = 256'h0502040401020200000009000200040602030501020300010201020403040602;
    encBuf[1028] = 256'h0204010203010103020306020303030404010303020403030404020303020304;
    encBuf[1029] = 256'h0103040303050203030302040102030305040304030402030102020103030306;
    encBuf[1030] = 256'h0403030403030202020302040404030503040203020201020102040305040303;
    encBuf[1031] = 256'h0303030202020303060304040303030302010201020403050403030402010200;
    encBuf[1032] = 256'h0001010306030503030402000200080202010604030403030303010202010404;
    encBuf[1033] = 256'h0306030304040103020102020203040305030205020203030103030203040103;
    encBuf[1034] = 256'h040004030103030103030903010b02010c04020806020802010b000a0f08090b;
    encBuf[1035] = 256'h01020a06020803020a01090e01080a04040105030204020801000a0101090703;
    encBuf[1036] = 256'h0106030003020801000a01010807030105020803000b08090d08080a03020005;
    encBuf[1037] = 256'h010a010a0f080a0c00080a03010803080b080b0f090a0a02020007030003000a;
    encBuf[1038] = 256'h01080c02020207050204020102000900000a04030207040103010000090b090a;
    encBuf[1039] = 256'h0b02020107020001090e0a0d0b0b0b0b090909000a0c0b0e0d0b0b0d0a0a0b08;
    encBuf[1040] = 256'h0a0a080a0c0a0c0c0a0c0b090a0a09090908090b080b0d090b0c080a0a000009;
    encBuf[1041] = 256'h03010804000901090c080a0c010808050201040009080c0e0a0c0c090b0a090a;
    encBuf[1042] = 256'h0b090b0f0a0b0e0a0c0a0b0a0c090a0b0a0a0c0a0c0c0a0b0c0a0b0c090a0a09;
    encBuf[1043] = 256'h0a09090a0a0a0b0d0a0b0c090a08000001020101010a0c0b0e0c0a0a0a090800;
    encBuf[1044] = 256'h0009090a0e0e0c0c0b0d0b0b0b0b0b0c0b0c0b0d0c0b0c0b0d0b0a0b0c0a0a0b;
    encBuf[1045] = 256'h0a0c0b0b0b0e0a0b0c0a0b0a0b0a0a0a0a0b0a0c0b0b0d0b0a0b0a0909080100;
    encBuf[1046] = 256'h01030000000b0b080c0904010506020303020101090b090c0a080a0003090002;
    encBuf[1047] = 256'h0e0c0b0f0c0a0c0b0a0c0b0a0b0c0a0c0b0a0c0c0a0b0c0b0c0b0a0b0c090b0a;
    encBuf[1048] = 256'h080a0a090c0b0a0d0b090b09010802040202030808000d0a000a010702040501;
    encBuf[1049] = 256'h02020008000a0b000c08020801050809000f0b0b0f0b0a0b0b0a0b0b090c0b0b;
    encBuf[1050] = 256'h0f0b0b0d0b0a0b0c090a0a090a0b090d0b0a0c0b0a0b0a000a00020801040001;
    encBuf[1051] = 256'h0300020701020601030501030402020402020402020302030501020402030401;
    encBuf[1052] = 256'h02030000010909000a08020901050808000f0b0a0f0a0a0b0a080a0800090908;
    encBuf[1053] = 256'h0e0a0b0d0b090b09010002050103030100020800050104070303060203030202;
    encBuf[1054] = 256'h0401020303040502040303030303020302020302030602020401020200010109;
    encBuf[1055] = 256'h01010a00020a00000b09000d09000c09000c09080d0800080307030505020403;
    encBuf[1056] = 256'h0203030204040304050304040203030303030303050304040304030304020102;
    encBuf[1057] = 256'h020101020203040304030102010809090b0a090a00000000090b0e0d0c0c0b0c;
    encBuf[1058] = 256'h0a0b0a0a0a090a0a0b0c0b0b0c0a0a0809010202050303050402040502040304;
    encBuf[1059] = 256'h0303040403030404030305020303030402030304030305020304020203010302;
    encBuf[1060] = 256'h0203030205030203040102020001000802010803040104030004020805010005;
    encBuf[1061] = 256'h0301060202040302040201040302050202050302040302030402030302050302;
    encBuf[1062] = 256'h03030203020801000a00080b02080d080c0f0a0d0c0a0c0b0a0b0b0b0b0d0b0d;
    encBuf[1063] = 256'h0b0c0c0b0c0a0b0b0b0b0a0b0c0b0c0c0a0c0a0b0a0a090a0909090a0a0a0d09;
    encBuf[1064] = 256'h0a0a080008040302050302040302050302060302040302040302040303040402;
    encBuf[1065] = 256'h0303020402020303030503020403020302000201000203020603030502010200;
    encBuf[1066] = 256'h0900080a02030107050103020101000900080a04030307050104010101010800;
    encBuf[1067] = 256'h000802020105020003010a000c0e090b0d090a0a0a0a0c0a0c0c0c0c0b0c0c0b;
    encBuf[1068] = 256'h0b0c0b0c0b0b0b0c0c0a0c0b0b0c0b0b0c0b0b0c0a0b0b0c0a0b0c0a0c0a0b0b;
    encBuf[1069] = 256'h0b0b0b0b0b0c0a0a0a0a090a0a0a0a0a09090802040405040304030203030303;
    encBuf[1070] = 256'h0503050503030503030303030303030403040404030304020302010201010203;
    encBuf[1071] = 256'h0405020402030201010000000001020305030403020201000100090101010503;
    encBuf[1072] = 256'h0205020102010001080b080c0d090b0c090a0b090b0c0c0d0c0c0d0b0c0b0c0a;
    encBuf[1073] = 256'h0c0a0a0c0a0c0b0c0b0d0b0c0b0b0b0c0a0b0c0a0b0c0c0a0c0b0b0c0a0c0a0a;
    encBuf[1074] = 256'h0b0b0b0b0c0b0c0b0c0a0b0b0c0a0a0a0a0a0b0a0b0b0b0b0c0a0a0a08080801;
    encBuf[1075] = 256'h0201040303050403040503040304030502030402030402040302030403030303;
    encBuf[1076] = 256'h0403030403030403030303030303020303030502030303010202000800090801;
    encBuf[1077] = 256'h0102040202020b0c0d0d0b0b0b09000003050100000c0c0c0c0c0a0909000008;
    encBuf[1078] = 256'h01090b0d0f0b0c0b0c0a0b0b090b0c0a0d0c0b0d0b0b0c0b0b0c0b0a0c0c0a0c;
    encBuf[1079] = 256'h0b0b0d0b0a0c0a0b0b0c0a0b0c0a0c0b0a0b0b0b0c0b0b0b0c0a0c0a0a0b0b0a;
    encBuf[1080] = 256'h0a0a090a0a000908010801050104060204030403050203040303040304030403;
    encBuf[1081] = 256'h0403030402030402020303040303040302030302020201020201020401010200;
    encBuf[1082] = 256'h09080e0b0a0d0a0a0a0a0a0a0b0b0f0b0b0d0a0b0b0a090908000908080a0a09;
    encBuf[1083] = 256'h0b09020307060303050202030202040203060204030303030202020800020900;
    encBuf[1084] = 256'h030801030b0b0c0f0f0a0c0c0a0b0b0b0c0b0b0c0c0b0c0c0a0c0b0b0b0b0c0a;
    encBuf[1085] = 256'h0b0a0c0a0b0b0b0b0d0a0a0a0a09080801010204020304030404030603040403;
    encBuf[1086] = 256'h0403030403040303030404030303040304030203030303040203030204020201;
    encBuf[1087] = 256'h020001000908090b0b0b0e0b0b0d0b0c0c0b0b0d0b0b0b0c0b0b0c0a0b0b0a0b;
    encBuf[1088] = 256'h0b0b0a0b0a0a0908020305050503030503040304030403040403040303040303;
    encBuf[1089] = 256'h03040303030402040203020303030302030102010008090a0b0c0c0c0b0c0c0b;
    encBuf[1090] = 256'h0d0b0b0d0b0b0d0a0b0b0b0b0c0a0b0b0b0c0b0b0c0b090a0900000102030305;
    encBuf[1091] = 256'h0302050304050304040304030402040203020403030304030402030203020302;
    encBuf[1092] = 256'h020302020201020008090b0c0d0b0d0b0c0c0b0b0d0b0b0d0a0b0c0b0b0b0c0b;
    encBuf[1093] = 256'h0b0b0c0c090b0a0a0b0a090a0a00080801020105040204050204030306030204;
    encBuf[1094] = 256'h0304030304030402040303030403030402030302030303040202030302030201;
    encBuf[1095] = 256'h02000a080b0d0b0c0c0b0c0c0a0b0d0a0c0b0c0b0c0a0c0b0a0b0b0b0b0c0a0b;
    encBuf[1096] = 256'h0c0a0a0c090a0b09090900000802010003010004020207040305040203030202;
    encBuf[1097] = 256'h020101010002030204030201080c0d0d0c0c0b0b0c0a0c0a0a0c0b0d0b0d0b0c;
    encBuf[1098] = 256'h0a0c0a0a0b0a0a0b0b0b0c0b0c0b0c0a0b0b090a0a0808080000000101080303;
    encBuf[1099] = 256'h0307040306030403040304030304020303040204030304030304030202020102;
    encBuf[1100] = 256'h0201020303040403030200000a0d0c0b0d0a0b0a0a0a0a0a0b0e0c0c0c0b0c0c;
    encBuf[1101] = 256'h0a0a0b0a0a0a0a0b0c0b0d0c0b0c0a0b0b0a090a09090a0a0b0e0b0c0b0b0a0a;
    encBuf[1102] = 256'h09080000010008090c0c0b0d0a0a0a080000010100000a0d0c0c0c0b0b0c0a0a;
    encBuf[1103] = 256'h0a0a0b0d0a0d0b0c0c0b0c0b0b0b0b0b0b0c0b0b0b0d0a0c0b0b0c0b0b0b0a0a;
    encBuf[1104] = 256'h0a08080000020001020001030307050404040304040203030202030305030403;
    encBuf[1105] = 256'h05030304020202020201020103030405020203010100090a0a0d0a0a0a090008;
    encBuf[1106] = 256'h08010b0c0b0f0d0b0c0b0b0b0b0a0a0b0b0d0b0c0c0c0a0c0b0a0a0b090a0a0a;
    encBuf[1107] = 256'h0a0b0b0e0b0b0c0c090b0a090a09080a09080a0a080c0b090c09080900030204;
    encBuf[1108] = 256'h070101040000000809000a08030105060102040800010a0a080c080109020400;
    encBuf[1109] = 256'h02010a0c0b0f0b090b0901000504020402010202080103020605030504020402;
    encBuf[1110] = 256'h0303040204030304030404030303040303030303040203040203040203030202;
    encBuf[1111] = 256'h020101000808080908080a09090d0c0b0f0b0c0c0b0b0b0c0a0a0a0a0a0b0a0b;
    encBuf[1112] = 256'h0c0a0c0a0a0a0a09080808000801000001010404030505030404030403020402;
    encBuf[1113] = 256'h0202020101020002020103040102030808090c0c0a0b0b090901010001090e0c;
    encBuf[1114] = 256'h0c0d0b0a0a090801020304040203030403070304050304040303040302040303;
    encBuf[1115] = 256'h0403030503030502040303030502030304020302030402040203040203020302;
    encBuf[1116] = 256'h0201020202030303030202090a0d0e0b0d0b0c0b0b0b0d0b0b0d0b0c0b0c0a0c;
    encBuf[1117] = 256'h0a0a0b0b0a0b0c0a0c0b0a0b0b0a0a0a08080900010803030406030504040304;
    encBuf[1118] = 256'h0303030403030402030402030303030402020301020201020008090a0d0b0d0c;
    encBuf[1119] = 256'h0b0c0c0b0b0d0b0b0c0c0b0b0b0c0b0a0a0a090a0a090a0a09090b0001000405;
    encBuf[1120] = 256'h0206030305030304040204030304040203040303030303040202030202020202;
    encBuf[1121] = 256'h020202000008090c0c0c0c0b0c0b0b0b0d0b0c0c0b0c0c0b0c0b0b0b0b0a0b0c;
    encBuf[1122] = 256'h0a0b0c0b0c0b0b0c0a0a0a0909090a090a0c0b0c0b0b0a090002020703020402;
    encBuf[1123] = 256'h0202020102030206040305030304030204020202030204030304040203030203;
    encBuf[1124] = 256'h010808090b0c0a0c0a090b0a0b0d0c0c0d0b0c0b0a0b0c09090908080a090b0d;
    encBuf[1125] = 256'h0a0b0c0909080103020703020404010402020403040304030304020202020102;
    encBuf[1126] = 256'h000101010101000009090d0d0c0c0c0c0c0b0b0c0c0a0b0b0b0c0b0c0c0b0c0a;
    encBuf[1127] = 256'h0c0a0a0b0a0a0a0a0a0a0a090a0b0a0a0a080000040403060303040303030503;
    encBuf[1128] = 256'h04030305030403030203030302010102010201020203020008090c0e0c0c0c0b;
    encBuf[1129] = 256'h0c0b0b0b0c0b0b0b0d0b0c0b0c0b0b0a0b0a0a0a09090a090b0a0c0a0a090002;
    encBuf[1130] = 256'h0306040402040202010202030403060304040304030203020202020001000100;
    encBuf[1131] = 256'h00000108090a0d0d0b0e0c0a0c0b0c0b0b0c0c0b0b0d0b0c0c0b0b0b0c0b0b0c;
    encBuf[1132] = 256'h0b0b0c0b0b0c0a0c0a0b0a0b0b0a0b0a090b0a090a0909090808010203040503;
    encBuf[1133] = 256'h0405030503040403030403030304020304020303020303020402020203000002;
    encBuf[1134] = 256'h09090a0f0b0c0d0b0b0c0b0b0c0b0b0c0b0b0d0b0b0d0b0a0c0a0a0b0a0a0b0b;
    encBuf[1135] = 256'h090b0a0909000000020401030601030502040402040304030303040402020302;
    encBuf[1136] = 256'h02040101020001010800010800000b0b090f0d0a0d0b0b0d0c0a0b0c0a0c0b0a;
    encBuf[1137] = 256'h0b0c0a0b0b0a0b0b0b0d0b0b0d0a0b0b0a090908000102030203030002030104;
    encBuf[1138] = 256'h0503060403050303040402030402030403030303030401030201020401030501;
    encBuf[1139] = 256'h03040203030201020900000c09080a00010004050102020808080e0a0a0d0a08;
    encBuf[1140] = 256'h0a08000801020801040105040305040303030203020001000103070405040305;
    encBuf[1141] = 256'h0303030401020201010001010302030603030403020202010009090a0c0b0b0c;
    encBuf[1142] = 256'h0b0a0c0b0b0b0b0c0b0b0b0b0a0b0b0c0e0b0b0e0b0c0a0a0908020504040404;
    encBuf[1143] = 256'h0204020102020102020304040404040304030304020303030302030303030302;
    encBuf[1144] = 256'h030203030305030404030304020201090a0c0d0b0d0b0a0a0a08000003030103;
    encBuf[1145] = 256'h000a0a0c0f0a0a0b090808040402050402030303040301030302040201030302;
    encBuf[1146] = 256'h05030307030305030305020202010000080a0a0b0b0a09080204030602020202;
    encBuf[1147] = 256'h09080a0f0a0c0c0a0a0c0a0a0a09080a000008020809000a0f090b0e090a0a08;
    encBuf[1148] = 256'h0000040403060303040302040200030101020302070303060303050302030302;
    encBuf[1149] = 256'h03010101010800010902010003030105020002090e0a0d0e0a0c0c0b0b0d0a0a;
    encBuf[1150] = 256'h0b090a0b09090b0a0a0c0a0b0e0a0b0c0a0b0c09090a00000004030305030103;
    encBuf[1151] = 256'h0200020100030303070503040303040303030201020009080b0d0a0b0c090b0a;
    encBuf[1152] = 256'h080a0a080a0d0b0f0c0b0d0b0c0c0b0b0c0b0b0b0b0b0a0b090a0a090a0b0b0c;
    encBuf[1153] = 256'h0e0a0b0c0a0a0a09000002030405030204030203030204020203020304040306;
    encBuf[1154] = 256'h030305030203020101080b0a0d0c0b0c0b0a0b0a0b0b0b0b0d0c0b0d0c0c0c0b;
    encBuf[1155] = 256'h0c0c0b0b0c0a0b0b0a0a0b0b0b0c0b0b0d0b0b0c0b0b0b0c0a0b0b0a0b0a0909;
    encBuf[1156] = 256'h0800000302030202010109090000010704040504030402040201020101000009;
    encBuf[1157] = 256'h0a090b0b0a0c0a090b0b0a0e0c0c0d0b0d0c0c0a0c0b0b0d0a0b0b0b0a0b0c09;
    encBuf[1158] = 256'h0b0a0a0b0c0b0d0b0c0b0c0a0b0a0a0a08080000010100020801020001050103;
    encBuf[1159] = 256'h070102030203060103040202040102030008010a0a080d0a080c0a080b0a080d;
    encBuf[1160] = 256'h0b0a0f0c0a0d0b0c0b0c0b0b0c0a0a0a0a0a0b090c0b0b0c0c0a0b0c090b0b0a;
    encBuf[1161] = 256'h0b0b0a0b0b080a09020003070101030001030900040003070304060203030303;
    encBuf[1162] = 256'h040202030001040101050102040202050101030000020908000900010a00030a;
    encBuf[1163] = 256'h09010e0b080d0a010a08020b09080f0d0a0d0b0a0b0900080206020204020102;
    encBuf[1164] = 256'h0900000800020105070202050203040203040203030204030204030304030204;
    encBuf[1165] = 256'h040103030303050102040101010000000900020003060205040102020000000a;
    encBuf[1166] = 256'h09090a0801010306020403020403030403040305020303020402020403040403;
    encBuf[1167] = 256'h0404030304030303040203030204030204030404030404030303030302020201;
    encBuf[1168] = 256'h0102030404040305030203040202020202020103020002010002030307050204;
    encBuf[1169] = 256'h0401030201010109000808000101050402050402030402040301030201020108;
    encBuf[1170] = 256'h0303030704030503020403020402020302020303010402000304020504030503;
    encBuf[1171] = 256'h02030302010009080a0c08000903030107040103020104020003010900090d08;
    encBuf[1172] = 256'h090b010300070601040301030301020108020208040301060302050401040202;
    encBuf[1173] = 256'h02020001010a00080b00000904020905010901080d000b0d090b0e0a0c0c0b0b;
    encBuf[1174] = 256'h0e090a0b080909000009000a0d0a0c0c0b0b0c0a0a0a08080901010804010002;
    encBuf[1175] = 256'h010a020a0e080a0c08080a03040107030103020002000b090c0d090b0d090b0c;
    encBuf[1176] = 256'h08090a00080901000c080d0e0a0c0d0a0b0b0a0a0b09080a08090a09090d090b;
    encBuf[1177] = 256'h0d0a0b0c0a0c0b0a0b0b090908030202070301030100010a0c090b0c0a0b0c08;
    encBuf[1178] = 256'h000804030306030201000b0c0e0d0b0c0b0a0b0b0a0a0a080a0c0b0d0c0c0b0d;
    encBuf[1179] = 256'h0b0b0d0a0b0b0b0c0b0a0b0b0a0b0b0b0b0c0b0c0c0b0c0c0a0b0b0a0b0b090a;
    encBuf[1180] = 256'h080000010302030402010108090a0b0a0801030705050303030302020000090b;
    encBuf[1181] = 256'h0c0b0c0d0a0c0b0b0c0b0b0d0b090b0c0a0d0b0c0c0c0b0c0b0b0c0b0a0a0a09;
    encBuf[1182] = 256'h09080908090a0a0d0b0c0c0b0a0b090900010304050402030203020101010001;
    encBuf[1183] = 256'h030101060102040101040002030000020a0c0a0f0e0a0c0c0a0c0a0a0b0a0a0b;
    encBuf[1184] = 256'h0b0a0d0b0b0e0b0b0d0b0b0c0b0a0b0a0a0b0a090a0a0a0b0b0b0d0a0b0c0b0a;
    encBuf[1185] = 256'h0b0a080900030206050304040304030202030001030801030204060204050202;
    encBuf[1186] = 256'h040102010000000a0a080b0b090b0a000b0a090f0b0a0f0a0b0c0c0a0b0b0a0d;
    encBuf[1187] = 256'h0b090c0a0a0a0b090a0a080a09000b0a080c0a090b0802010705030604020304;
    encBuf[1188] = 256'h0303030203040202030303060203040303050202030101020800000a0a090c0b;
    encBuf[1189] = 256'h090d0a090d0a090d0a0a0c0c0a0b0d0a0c0b0a0c0a0a0a0a090a09080a09090b;
    encBuf[1190] = 256'h0b0a0e0a09090801000505020405020304020304020203020304030305030305;
    encBuf[1191] = 256'h0303040303040203030202040101010001000800010802030204040002020b0c;
    encBuf[1192] = 256'h0b0f0c0a0c0b0a0b0a080909080908080b0a0b0f0a0b0c0b090b0a0000030504;
    encBuf[1193] = 256'h0504020403020304010303020304030404030404030403040304020303020202;
    encBuf[1194] = 256'h0101010100020202050203040203020008080b0d0b0d0b0c0b0b0b0c0b0a0b0b;
    encBuf[1195] = 256'h0a0c0b0a0c0b0c0c0b0b0c0a0b0a090a08010005040305030403040203030202;
    encBuf[1196] = 256'h0203040503060304040304030303030202020102010203030503030503030303;
    encBuf[1197] = 256'h03030202010009090b0d0c0b0c0b0b0a090b000100010208000b0f0c0d0b0c0a;
    encBuf[1198] = 256'h0c09090901010306030304030203020002000802030307050304040304040203;
    encBuf[1199] = 256'h030303030303020102020102040205040306020304020202020000080b090b0c;
    encBuf[1200] = 256'h0a090a010000050202030208010b0f090c0d0a0a0b0a090a0000000302000503;
    encBuf[1201] = 256'h0801010801090d01000a04020107050205030304040103030003010001010003;
    encBuf[1202] = 256'h040207030304030304030103010801080a00090a00080a050201060201040108;
    encBuf[1203] = 256'h01080c090b0e090b0b09090b02010805030004020804000b01090c000a0d0101;
    encBuf[1204] = 256'h0904040106020204010003000901080a00080a05020107040105020103020102;
    encBuf[1205] = 256'h010901090a00000b05030106040104030104020003000902080c080a0c090a0d;
    encBuf[1206] = 256'h00080902000904000b000c0f0a0b0f090a0c09090b08090a08090c080a0d090a;
    encBuf[1207] = 256'h0d0a0a0b0a0a0c09090a00080902000804000902000a03080c01000a02010007;
    encBuf[1208] = 256'h030207040104020102010800090c090b0d09090a00000902090c080c0f0a0b0d;
    encBuf[1209] = 256'h0a0c0c0a0b0b0b0c0b0a0c0c090b0b0a0c0a0b0b0c0a0c0b0b0c0b0b0b0c090a;
    encBuf[1210] = 256'h0a09090900080900090c090a0b0a090901030506040304020203020002090800;
    encBuf[1211] = 256'h090a00090c090b0d090c0c0a0c0b0d0b0c0b0e0b0c0c0c0b0c0b0b0c0b0b0c0b;
    encBuf[1212] = 256'h0a0b0c0a0c0a0c0a0c0a0b0b0c0b0b0a0b0b0b0b0a0b0b0b0b0b0c0a0b0b0b0b;
    encBuf[1213] = 256'h0a0909000000030405040303070201030202030101020009010a080209080408;
    encBuf[1214] = 256'h09020f0b0a0f0d0a0d0b0b0d0b0a0c0b0a0c0b0a0b0c0a0c0b0a0c0b0b0c0c0a;
    encBuf[1215] = 256'h0b0b0a0c0a0a0b0a090a0a080a09000909020a08030900070001060103050303;
    encBuf[1216] = 256'h050202040102020102030002030103060002030801030a0a010f0c0a0c0c0a0d;
    encBuf[1217] = 256'h0b090c0b0a0c0a0a0b0c0a0b0c0a0c0b0b0c0b0b0c0b0b0b0c090b0a080a0900;
    encBuf[1218] = 256'h0909010800020801040004060103060203060202040202040202030203040103;
    encBuf[1219] = 256'h050102040102040101040001020000020808000a08080c09000c09000a0a000c;
    encBuf[1220] = 256'h09080e0b090d0a090c0a090b0801090205000305020304020305020305020403;
    encBuf[1221] = 256'h0305030305030304030305030203040203030303050202040202030303030303;
    encBuf[1222] = 256'h040101020000010801010800010801030908080c0a0c0d0a0b0e090a0b0a0909;
    encBuf[1223] = 256'h0001010406020503020503030304030403040304030503030503030403030403;
    encBuf[1224] = 256'h0303030403030304030305020303040203030303020303020303020304020203;
    encBuf[1225] = 256'h0203050203040302030202030901030a08030103060206040203040204020203;
    encBuf[1226] = 256'h0301050202040401030502030402040303040302040302030302030302040301;
    encBuf[1227] = 256'h05020204020203030103020803000a03010b04010b02080e00090e090a0c090b;
    encBuf[1228] = 256'h0b090b0c090a0c000a0b010a0c04000a05020004020904010802020905020006;
    encBuf[1229] = 256'h020205030104020103020104030004020004020802010b02090d00090d08090c;
    encBuf[1230] = 256'h08090c090a0e09090c0a0a0c09090c080a0b0a0a0d090b0b0a0b0d080a0a0009;
    encBuf[1231] = 256'h0b01090c01090d02080a04010805020805010003000803080b04000902080b02;
    encBuf[1232] = 256'h0a0f080a0c090b0d080b0c080a0c090c0c090a0d0b0b0c0b0b0e0a0a0c0a0b0c;
    encBuf[1233] = 256'h0a0b0b0b0b0d0a0a0b090b0b0a0b0b0b0c0c0a0a0c090b0b0a0a0c080a0a0809;
    encBuf[1234] = 256'h0a01090903010004020206020102010104010002090b080b0e0b0c0c0c0b0d0a;
    encBuf[1235] = 256'h0c0b0a0b0c0a0c0b0b0c0b0c0b0c0b0d0b0b0c0b0b0c0b0b0c0b0b0b0c0b0b0b;
    encBuf[1236] = 256'h0b0c0a0b0b0b0a0c0a0a0a09090a000008010302030303040401010202040305;
    encBuf[1237] = 256'h040203050202040202040100020008000a0b0b0f0d0a0d0b0b0c0c0a0c0b0a0c;
    encBuf[1238] = 256'h0c0a0b0b0c0b0c0b0b0c0a0b0c090b0a0a0b0a0b0d0a0b0c0a0a0b0a0a0b0908;
    encBuf[1239] = 256'h0808020203050205040304040203040203040103030103030303050103040002;
    encBuf[1240] = 256'h030001010908010b0a010e0b000d0c0a0d0c0a0d0c0a0b0c0b0b0d0a0b0b0b0c;
    encBuf[1241] = 256'h0b0a0c0a0a0b0b090b0a0a0b0b0a0c0b0a0c0a090a0900000204030604020305;
    encBuf[1242] = 256'h0203050203050303050204030203040202030302030303030203030202030001;
    encBuf[1243] = 256'h020900020c0a000d0a0a0f0b0b0e0b0b0d0b0b0c0b0b0c0b0a0c0a0a0b0b0a0b;
    encBuf[1244] = 256'h0a080a0801010306030603040304030403040304020304030304030403030404;
    encBuf[1245] = 256'h0203040303040203030204020201030101010100000808090c0a0b0d0b0b0d0b;
    encBuf[1246] = 256'h0b0b0b0c0b0a0b0c0b0a0c0b0c0b0a0d0b0a0b0c0a0a0a0a0a0a000801030405;
    encBuf[1247] = 256'h0503050304030403040303040304020402020402030303030502030402030304;
    encBuf[1248] = 256'h02030304030304030303030303020201020808000a0a0a0b0b0b0a080909080a;
    encBuf[1249] = 256'h0901000802010804020104020004020005030803050103040206030205030305;
    encBuf[1250] = 256'h040204030304030304030303030203030202010202000000010808000908090a;
    encBuf[1251] = 256'h080a09080b0c0a0c0c0b0d0c0b0d0c0a0b0c0a0c0a0b0b0d0a0a0b0a0b0b0a0a;
    encBuf[1252] = 256'h0a08080801000903000b000b0d090b0d090a0b00090a01000902010005020004;
    encBuf[1253] = 256'h040105020204020203030004020001020803000903000a020200040302070402;
    encBuf[1254] = 256'h0503030403020502010302010202010202000201000502010305020403020502;
    encBuf[1255] = 256'h0103020103010003000901080b080c0e0a0c0c0b0d0b0a0c0b0b0b0b0a0b0b0a;
    encBuf[1256] = 256'h0b0c090c0b0b0c0c0b0d0b0b0c0c0b0c0b0b0c0b0a0c0b0a0a0b0b0a0b0b0c0a;
    encBuf[1257] = 256'h0a0c0a0a0b0b0b0c0c0a0c0b0c0c0b0b0c0c0b0b0c0b0b0b0b0c0a0b0b0b0b0b;
    encBuf[1258] = 256'h0b0b0c0b0b0d0b0b0e0b0b0d0b0c0b0c0a0b0b0b0a0b0a0b0b090b0a0a0b0a09;
    encBuf[1259] = 256'h0809020303060303040203030302040304030504040304040403030404030304;
    encBuf[1260] = 256'h0304030304030303020303020203020202040202030203030102010808080a0b;
    encBuf[1261] = 256'h090b0b0c0b0e0b0c0c0c0b0d0b0b0c0c0b0b0b0c0b0b0c0b0b0b0b0a0b0a0b09;
    encBuf[1262] = 256'h0a090b0b0b0e0b0d0b0c0b0c0a0b0b0b0b0b0b0b0b0d0b0b0c0b0c0b0a0b0c09;
    encBuf[1263] = 256'h0b0d090b0d0b0c0c0b0c0c0a0c0b0a0c0b0b0c0b0c0b0b0b0c0b0b0b0c0a0a0b;
    encBuf[1264] = 256'h0a0b0c0a0c0b0b0c0b0b0c0b0b0b0a0a0b090809000100030503060403040403;
    encBuf[1265] = 256'h0403040304030403030502030403030403030502030304030403030403030403;
    encBuf[1266] = 256'h0303030304030203030304020203020302030203020303030204020302020101;
    encBuf[1267] = 256'h0908090d0a0b0d0a0b0c0b0b0c0b0c0d0a0b0b0b0c0b0a0a0a0a0909090a0b0c;
    encBuf[1268] = 256'h0c0c0c0d0b0c0c0b0c0b0c0b0c0b0c0b0b0d0b0b0b0d0b0b0c0b0c0b0b0c0b0c;
    encBuf[1269] = 256'h0b0c0a0c0b0a0c0b0b0b0c0b0c0a0b0b0c0a0b0b0b0b0b0b0c0a0a0a0a090a09;
    encBuf[1270] = 256'h0809080008020301060402050403040403040403040303050303040304030304;
    encBuf[1271] = 256'h0304020402030304030304020402030303040303040303030502030302040203;
    encBuf[1272] = 256'h020402020202030202030302030302040201020201020200020109000a0e090d;
    encBuf[1273] = 256'h0c0a0d0b0b0d0b0b0d0b0b0c0b0c0b0c0c0b0b0c0b0c0b0c0b0b0c0b0c0b0b0c;
    encBuf[1274] = 256'h0c0b0b0c0b0b0c0c0a0b0b0c0b0b0c0b0b0b0c0b0b0c0b0b0c0a0b0c0a0b0b0b;
    encBuf[1275] = 256'h0b0c0b0b0b0b0c0a0a0b0a0a0a0a090909080801020206030306040204030403;
    encBuf[1276] = 256'h0403050203040402030403030403050203040303040303040304030303040303;
    encBuf[1277] = 256'h0502030303040304020402030302040203030304020402020302030302030401;
    encBuf[1278] = 256'h020201010100010809090a0d0a0d0b0c0c0b0b0d0c0a0b0d0a0c0b0b0c0b0c0b;
    encBuf[1279] = 256'h0c0b0b0c0b0c0b0b0c0b0b0c0b0b0c0b0b0c0b0b0c0b0b0c0b0a0c0b0a0c0a0b;
    encBuf[1280] = 256'h0b0b0c0b0b0b0c0a0b0c0a0b0a0b0b0b0a0c0a0a0a0b0a0a0b0a0a0b090a0a00;
    encBuf[1281] = 256'h0900040104050304050204030404030305030305030304030404020304030403;
    encBuf[1282] = 256'h0304030304040203040303030404020304030303040303040203040203030303;
    encBuf[1283] = 256'h0403030402030302040202020201020100010008000a0a0b0d0c0b0d0c0b0c0b;
    encBuf[1284] = 256'h0c0c0b0c0b0c0b0c0b0b0c0b0b0d0b0a0c0b0a0c0b0b0b0c0b0c0b0b0c0a0b0c;
    encBuf[1285] = 256'h0a0b0b0b0c0b0b0b0b0c0b0b0b0c0b0b0b0c0b0a0c0a0a0b0a0b0b0a0c0a0a0b;
    encBuf[1286] = 256'h0b0b0b0c0a0a0b0a0a0a08090001010205020306020304030404030404030404;
    encBuf[1287] = 256'h0303050304030304040204030303040403030403030404020304020402030304;
    encBuf[1288] = 256'h0203040203040203030304030304030203040203020302030203020302020102;
    encBuf[1289] = 256'h010001080a090b0f0a0d0b0c0c0c0a0c0b0b0d0a0b0c0c0a0b0c0a0c0b0a0c0b;
    encBuf[1290] = 256'h0b0d0a0b0b0b0c0b0c0a0b0b0c0b0b0b0c0b0c0b0b0b0c0a0c0a0b0b0b0b0c0b;
    encBuf[1291] = 256'h0b0b0c0b0b0b0b0c0c0a0a0b0b0b0c0a0a0b0b0b0b0a0b0b090b0b0a0b0a090b;
    encBuf[1292] = 256'h0a00090005010506020306020305020403030403030503030403030503040303;
    encBuf[1293] = 256'h0403040303040304020304030204030303040304030303040303030403030304;
    encBuf[1294] = 256'h0303030403030303040303040203030203030203030201020001010808080a0a;
    encBuf[1295] = 256'h0c0c0b0e0b0c0d0b0c0c0b0b0d0b0c0b0b0c0c0a0b0c0b0c0b0b0c0c0a0b0c0b;
    encBuf[1296] = 256'h0b0d0a0b0b0b0c0b0c0b0b0b0c0b0b0c0b0c0a0c0a0b0b0a0c0b0a0b0c0a0b0b;
    encBuf[1297] = 256'h0a0c0a0a0b0b0b0b0b0b0c0a0a0b0a0909090808000201030602030602030403;
    encBuf[1298] = 256'h0404020403040304030403030404020402030304020402030402030403030403;
    encBuf[1299] = 256'h0304030303040304030204030303040304030304030304020402030303030403;
    encBuf[1300] = 256'h03040302040203030402030303030303040202020202010100010808090b0c0b;
    encBuf[1301] = 256'h0e0b0c0d0c0a0d0a0c0b0b0c0c0b0b0c0b0b0d0a0b0c0b0b0c0c0a0b0c0a0c0a;
    encBuf[1302] = 256'h0b0b0b0c0b0b0c0b0b0b0c0a0b0c0a0b0b0b0c0a0b0b0b0b0b0b0b0b0b0b0a0b;
    encBuf[1303] = 256'h090a0a0809000101020502060304040304040402040303040303050203040302;
    encBuf[1304] = 256'h0403030304030403040303040304030303040303040303040303040402030303;
    encBuf[1305] = 256'h0403030403030305020303030305020303040303030403020402020303020303;
    encBuf[1306] = 256'h0203020203020202020002080a090d0d0a0d0c0b0d0b0c0c0b0b0d0b0b0d0b0a;
    encBuf[1307] = 256'h0d0a0b0c0b0b0c0b0c0b0c0a0c0a0b0b0b0c0b0b0b0d0a0b0b0c0a0b0c0a0b0b;
    encBuf[1308] = 256'h0c0a0b0b0a0b0b0b0c0a0a0a090a0a0909090808080101020306030404040205;
    encBuf[1309] = 256'h0203040303050204020304030304040203040203040303040203030304030303;
    encBuf[1310] = 256'h0402030402030402030402030402020303030303030402040202030303030402;
    encBuf[1311] = 256'h03030203030104020003020102020003010a00090d080c0d0b0c0d0a0d0b0b0d;
    encBuf[1312] = 256'h0b0b0c0c0a0c0b0b0b0d0a0c0b0b0c0b0c0b0c0b0c0b0b0c0b0c0b0b0c0b0b0c;
    encBuf[1313] = 256'h0b0b0c0b0c0a0b0c0a0b0b0b0c0a0b0b0b0b0c0a0b0b0a0b0b0b0c0a0a0a0909;
    encBuf[1314] = 256'h0a08000103040404050303050304030403040304030305020304030304030304;
    encBuf[1315] = 256'h0303040303040303030403040203030304030303030304030202040102020101;
    encBuf[1316] = 256'h020201020101020002010009090a0c0c0c0b0d0d0a0c0b0b0c0b0b0d0b0b0c0b;
    encBuf[1317] = 256'h0b0b0d0b0b0c0b0b0c0b0c0b0b0c0b0b0c0b0c0b0b0c0c0b0b0b0d0a0c0a0b0c;
    encBuf[1318] = 256'h0b0b0b0c0b0b0c0b0b0b0c0c0a0b0c0a0c0a0b0b0c0a0b0c0a0b0b0b0c0a0b0b;
    encBuf[1319] = 256'h0b0a0b0b0b0b0b0a0c0909090800080204020405020404030404030403040304;
    encBuf[1320] = 256'h0403030404030303050303040204030204020303040204020203030402030304;
    encBuf[1321] = 256'h020303030304030203020302030202020101010008080b0c0b0d0c0b0c0c0b0c;
    encBuf[1322] = 256'h0b0c0b0c0b0b0c0c0a0c0a0b0b0c0b0b0d0a0b0b0c0b0b0b0c0b0b0c0b0b0b0b;
    encBuf[1323] = 256'h0c0b0a0c0b0a0b0b0b0c0b0b0c0b0b0b0c0a0b0c0a0c0a0a0b0b0b0c0b0a0c0b;
    encBuf[1324] = 256'h0a0b0c0a0a0c090a0c090a0b0a0a0c0a0b0b0a0c0b090a0a0909000100030602;
    encBuf[1325] = 256'h0307020304030404020403040304030305030305030303040403030403030502;
    encBuf[1326] = 256'h0304030204030204030204020303040203030303040203030303040302030302;
    encBuf[1327] = 256'h0303020201020100090a090d0c0a0b0e0b0b0c0c0b0c0a0c0b0b0c0b0b0d0b0a;
    encBuf[1328] = 256'h0c0b0a0c0a0b0b0b0c0a0c090b0b0a0b0c0a0a0b0b0a0b0b0b0b0a0a0a090908;
    encBuf[1329] = 256'h0101000201030502020202040502020303040403040303040203040302030302;
    encBuf[1330] = 256'h0203040201020301010100000101080a090a090a0b0c0a0c0b0a0c0b0a0a0c0b;
    encBuf[1331] = 256'h0a0c090a0a090b0b08090a090809000200080204030303050402040402030304;
    encBuf[1332] = 256'h0403030403030602020403030403020403040202030402020304020203030304;
    encBuf[1333] = 256'h0204020203020104020003010002020801010802080a01000a02080c08090a00;
    encBuf[1334] = 256'h0a0c01080b02000a030400030301070300040400030202040301050301040302;
    encBuf[1335] = 256'h040302040203040101030300020109010809080d0d0a0b0e0a0b0e0a0c0b0b0d;
    encBuf[1336] = 256'h0b0b0d0b0b0c0c0a0b0c0b0c0a0c0a0b0c0b0b0b0d0a0b0c0a0b0c0a0b0b0b0b;
    encBuf[1337] = 256'h0c0b0b0b0b0c0a0b0b0b0a0b0b0a090b0a090800000203040504030404040303;
    encBuf[1338] = 256'h0503030503030503030305030304030304030303040304020303040203030403;
    encBuf[1339] = 256'h0203040302040202030202030402010302020202020302020103010801080900;
    encBuf[1340] = 256'h080b080b0b090a0b080d0b080b0d0a0d0b0a0f0a0a0c0b0b0d0b0b0c0c0a0c0b;
    encBuf[1341] = 256'h0a0d0a0b0c0b0b0c0b0c0c0b0b0c0b0c0b0c0b0c0a0b0c0b0c0b0a0c0b0b0b0d;
    encBuf[1342] = 256'h0a0b0b0c0a0c0a0a0b0b0b0b0c0a0c0a0a0a0b0b0a0a0b0b090b090908000102;
    encBuf[1343] = 256'h0307030404030404030404030305020403030305030304030304030403020403;
    encBuf[1344] = 256'h0304020304020303040203030304030203030204020202020202020102010000;
    encBuf[1345] = 256'h0008090a0b0c0c0c0d0a0c0b0c0b0c0c0a0c0b0a0c0b0c0b0b0b0c0c0a0b0c0a;
    encBuf[1346] = 256'h0c0a0b0b0b0c0b0c0a0c0a0a0c0a0b0b0b0c0b0c0b0b0b0c0b0b0c0b0b0c0b0b;
    encBuf[1347] = 256'h0b0d0a0b0a0b0d0a0a0c0a0a0b0b0b0c0b0a0b0c0a0b0b0a0b0b0a0b0b090b09;
    encBuf[1348] = 256'h000a010202060303070402040304030503040303050303040402040303040303;
    encBuf[1349] = 256'h0502030403020403030304030304030303040303030403020304020303020303;
    encBuf[1350] = 256'h020303010202020000080a0a0c0c0c0c0c0b0c0c0b0c0b0c0b0c0b0c0b0c0b0b;
    encBuf[1351] = 256'h0c0b0b0c0b0c0b0b0c0b0b0c0b0b0c0a0b0c0a0b0b0c0a0b0b0b0b0c0b0b0a0b;
    encBuf[1352] = 256'h0c0a0b0b0b0b0b0b0c0a0a0a0b090b0a090b09000a0802090106000206020204;
    encBuf[1353] = 256'h0304030306030204030205030204040203040204030305020304030304030305;
    encBuf[1354] = 256'h0203040303040204030303040303050203030402030402040202030304020303;
    encBuf[1355] = 256'h04020303020402020203020302020202020100000008090a0d0b0c0d0b0c0c0b;
    encBuf[1356] = 256'h0c0c0b0b0d0b0b0b0d0b0b0c0b0c0b0a0c0b0b0c0b0b0b0c0b0c0a0b0b0c0a0b;
    encBuf[1357] = 256'h0b0b0b0c0a0b0b0a0b0c090b0a090a0a08080901000004040204040204040303;
    encBuf[1358] = 256'h0502040303040402040302030502030402030402030304020402030302040302;
    encBuf[1359] = 256'h03030304030204020203030203030203030203040101010001010901000c0809;
    encBuf[1360] = 256'h0c08090d080a0c08090b080a0c000a0c00080b02080b03080b07000903020904;
    encBuf[1361] = 256'h0308060208040301030402050201040202040201050101030202030201040201;
    encBuf[1362] = 256'h04010004010003010803020904000b06000b01000b00080d00080b00090c0809;
    encBuf[1363] = 256'h0c01090a04090b05000902010005000905010803020905010904010802010903;
    encBuf[1364] = 256'h090a03090c020a0f08090c090b0d0b0c0b0c0c0b0b0e0b0b0c0c0a0c0b0b0c0b;
    encBuf[1365] = 256'h0b0c0c0a0c0a0b0c0a0b0c0b0b0b0c0b0b0c0b0b0b0c0b0b0b0c0b0a0b0c0a0a;
    encBuf[1366] = 256'h0a0a0a0a09090908080000020306030403060204030305030304030403040304;
    encBuf[1367] = 256'h0303040402030402030304030302040303030402030303030402030302030302;
    encBuf[1368] = 256'h030302030200010108000a0c0b0d0c0b0d0b0c0c0c0a0c0b0b0c0c0a0b0c0b0c;
    encBuf[1369] = 256'h0b0b0b0d0a0c0a0b0c0b0b0b0c0c0b0b0b0d0a0c0b0a0b0d0a0b0b0b0c0c0a0b;
    encBuf[1370] = 256'h0c0a0b0c0a0b0c0b0b0b0c0b0c0a0c0a0b0b0c0a0c0a0b0b0b0b0b0d0a0b0b0a;
    encBuf[1371] = 256'h0b0c090b0a0b0b0a0a0b0a090a09000a08030104050205040204050203040304;
    encBuf[1372] = 256'h0403030404030303050303030502040203030304030403030304030303050203;
    encBuf[1373] = 256'h03030304030304020302030303030303030202030101020009010a0b0c0d0c0a;
    encBuf[1374] = 256'h0d0b0c0c0c0a0b0d0a0c0b0b0c0c0b0b0c0b0c0b0b0c0c0a0b0c0a0b0c0b0b0b;
    encBuf[1375] = 256'h0c0b0c0b0b0c0a0b0c0b0b0c0a0b0c0a0b0b0b0c0b0b0c0b0a0b0b0b0c0b0a0b;
    encBuf[1376] = 256'h0b0a0c0b090b0a090a0a090a0801090005080307010204020404030305030403;
    encBuf[1377] = 256'h0403040204030304040203040204020303040304030204030303050203030403;
    encBuf[1378] = 256'h0303040302040303030402030304020303030303040302030303030303020302;
    encBuf[1379] = 256'h010101000a0a0b0d0d0c0b0c0d0a0c0b0c0b0c0b0c0b0c0b0c0a0c0b0b0b0d0b;
    encBuf[1380] = 256'h0b0b0c0b0c0b0b0d0a0a0c0a0a0b0c0a0b0b0b0b0c0b0b0b0b0c0a0b0b0a0b0b;
    encBuf[1381] = 256'h0b0b0b090a0a080a080101020403060403050402040403030403040403030403;
    encBuf[1382] = 256'h0403030403040303040304020402030304020402030303040303030502030303;
    encBuf[1383] = 256'h0305020203030304020402020203030204020303020304010302030203020302;
    encBuf[1384] = 256'h0003010801080b09090f0a0b0e0a0c0b0a0d0c0a0b0c0b0b0d0a0c0b0b0b0e0a;
    encBuf[1385] = 256'h0a0c0a0b0c0a0c0a0b0b0d0a0a0c0a0a0b0b0c0b0a0c0a0b0a0c0a0a0b0b0b0b;
    encBuf[1386] = 256'h0a0c0b090a0b080a0a0800080203020603040504020404020403030404030305;
    encBuf[1387] = 256'h0203040303040303050203030403030304040203030303040303040302040202;
    encBuf[1388] = 256'h0302020302040201020200020108000009000b0d090b0f090a0c0b0b0c0b0c0d;
    encBuf[1389] = 256'h0a0a0c0b0a0d0a0a0c0a0b0b0c0b0b0b0c0c0a0b0b0b0c0b0b0c0b0a0c0b0b0b;
    encBuf[1390] = 256'h0c0a0b0c0a0b0b0b0c0b0a0b0c0a0a0c0a090b0a0b0b090c0a090a0b08090b09;
    encBuf[1391] = 256'h080b00010a010302030403070201050302050303040402030502030303060202;
    encBuf[1392] = 256'h0403010403020402020403020304020304010303030304010303010303010301;
    encBuf[1393] = 256'h0802090b090d0c0a0d0c0b0c0c0b0d0b0b0c0c0b0c0b0b0d0b0b0d0a0b0c0b0b;
    encBuf[1394] = 256'h0c0b0c0b0c0a0b0c0a0c0a0b0b0c0a0c0a0b0b0b0c0b0a0c0b0a0b0c0a0b0b0b;
    encBuf[1395] = 256'h0b0c0a0b0b0b0b0b0b0b0b0b0b0b090a0a000800030204050306030403040403;
    encBuf[1396] = 256'h0403040303050303040304030402030403030402040203040203030303050202;
    encBuf[1397] = 256'h03040202030303030303040203030202020202010001000a0a090e0b0b0f0b0a;
    encBuf[1398] = 256'h0d0c0a0b0c0b0c0b0c0b0c0b0c0b0b0d0b0a0c0b0b0c0c0a0b0b0b0d0b0a0c0b;
    encBuf[1399] = 256'h0a0c0b0b0b0c0b0b0c0a0c0a0b0b0b0b0d0a0a0b0c0a0a0b0a0b0c090b0b0a0a;
    encBuf[1400] = 256'h0b0a0b0a090b0900090002000406010405020205020403030503030503030403;
    encBuf[1401] = 256'h0403040303040304030304040203040203040203030403030304030303040303;
    encBuf[1402] = 256'h03030403030303030304020203010202000001080a0a0c0b0c0e0b0b0d0b0c0b;
    encBuf[1403] = 256'h0d0b0b0c0b0c0c0a0c0a0b0c0b0b0b0d0a0b0c0a0c0a0b0a0c0a0b0b0c0a0b0b;
    encBuf[1404] = 256'h0c0a0b0b0b0b0b0d0a0a0a0b0a0a0a0b0a0a0a09090908010802060103040305;
    encBuf[1405] = 256'h0403040402040304030304040303050302040303040304030304030403030304;
    encBuf[1406] = 256'h0402030403020403020403030303040402030303040302040302030402030302;
    encBuf[1407] = 256'h03040202030302030202030102010801080b0a0c0d0c0c0b0b0e0b0b0d0b0c0b;
    encBuf[1408] = 256'h0c0b0c0b0c0b0c0a0c0b0b0c0b0b0c0b0c0b0b0c0b0b0b0d0a0b0b0c0a0b0c0a;
    encBuf[1409] = 256'h0b0b0b0c0b0a0b0c0a0b0b0a0c0a0a0a0a0a0a0a0a0909090900080202020503;
    encBuf[1410] = 256'h0504030404030305030404020304030403030403040303040304030204030304;
    encBuf[1411] = 256'h0303040303040303030403030403030304030402030303040203040202030303;
    encBuf[1412] = 256'h030304030203030203030203020102010802090b080e0c090c0d090c0c090b0d;
    encBuf[1413] = 256'h0a0b0c0a0c0c0a0b0b0c0b0c0a0c0b0b0c0b0b0c0b0b0c0b0b0c0b0b0c0c0a0b;
    encBuf[1414] = 256'h0b0a0c0b0b0b0b0c0b0c0a0b0b0a0b0c0b0a0c090b0a0b0a0a0b0a0a090b0a09;
    encBuf[1415] = 256'h0900000901030303040503030604020204030403030403040402030304030402;
    encBuf[1416] = 256'h0304030304020304020303040303020403020304020203030303030403010302;
    encBuf[1417] = 256'h0202030201000801080b00090c08090e090a0a0b0c0c0a0b0e0a0a0b0b0c0c0a;
    encBuf[1418] = 256'h0a0c0a0b0b0b0c0b0b0c0b0b0b0c0b0b0b0b0d0c090a0b090a0c0a0a0a090b0b;
    encBuf[1419] = 256'h0b0a0b090a090a0d09000a0b09080809090a080a0a0a080a0a09090a0a0a0a0a;
    encBuf[1420] = 256'h0b0b0a0b09090c0b090b0b0b0d0b080b0b0b0b0c0a0a0e0a080b0b090b0c0a0b;
    encBuf[1421] = 256'h0a0a0b0d09090a0a0b0b080a0b09090909090a09090908090a08080908090908;
    encBuf[1422] = 256'h090909090808090908090a08090c09080a0a0a0a0a0c0b080b0d08090b0a090b;
    encBuf[1423] = 256'h0b0c0b080b0e09090a090a0a09090c0a090a0a0a09080a08000b0b0000000809;
    encBuf[1424] = 256'h0901000802000902010802000002010001000001000801000000000800000809;
    encBuf[1425] = 256'h0908080b0a090c0b080b0d090b0d090b0c0a0c0a0b0c0c0a0c0b0a0c0b0b0b0d;
    encBuf[1426] = 256'h0a0b0c0a0c0a0a0c0b090c0b0a0b0c0a0b0b0b0c0b0a0c0b0a0b0b0b0c0b080a;
    encBuf[1427] = 256'h0a0a0b0a0a0a0808080801010101020403010404020304040304020404030303;
    encBuf[1428] = 256'h0404030305030303040304030403020403030304040303030404020303040203;
    encBuf[1429] = 256'h0403030304030402030402030402020402030203040203030403020402020302;
    encBuf[1430] = 256'h030304020202040102020201020201010809080909090b0a0a0c0b0a0d0c0b0c;
    encBuf[1431] = 256'h0c0b0c0b0b0c0c0b0b0c0b0c0b0c0b0c0b0b0c0b0c0b0b0c0b0c0a0c0a0b0b0c;
    encBuf[1432] = 256'h0b0b0b0c0b0c0a0c0a0b0b0b0b0c0b0b0b0b0c0b0b0b0c0b0b0a0b0a0b0a0a0b;
    encBuf[1433] = 256'h0b09090808080803000304030404030504030305030304030404030304030403;
    encBuf[1434] = 256'h0304030403040303030404020304020304020304020303040302040303030304;
    encBuf[1435] = 256'h0303030404020203030402030203030304030203030304020202040102010100;
    encBuf[1436] = 256'h010001000900090a090b0e090a0b0c0c0b0b0c0c0b0d0a0b0c0a0b0c0b0c0b0b;
    encBuf[1437] = 256'h0c0c0b0a0c0b0b0c0b0a0c0b0b0c0c0a0b0a0b0c0b0b0b0d0a0b0a0b0c0b0b0b;
    encBuf[1438] = 256'h0c0b0a0a0b0b0b0b0d0a0a0a0a0a0a0a0a090a00000800080100020403040303;
    encBuf[1439] = 256'h0306020403040303050303030503030403030403040203040303030403030403;
    encBuf[1440] = 256'h0402030303040203030403030203040304010203020203020103020302010001;
    encBuf[1441] = 256'h01080108000809090a0a0a090a090a0b0c090b0c0b0b0c0c0b0b0b0c0a0a0b0c;
    encBuf[1442] = 256'h0c0c0b0c0b0a0a0a0c0b0b0b0c0a0b0c0b0b0b0c0b0b0a0c0b0b0c0b0b0b0a0b;
    encBuf[1443] = 256'h0c090a0b0a080a09080a0a080a08000909080800000900010001000001020008;
    encBuf[1444] = 256'h0201020102020203020102020101020202010101020202020302030102030200;
    encBuf[1445] = 256'h020100020202030100010201010801010808010002010808000808010a090009;
    encBuf[1446] = 256'h0a000809080a090809090a09080a0b09080a0a090a0a0a0a0a0b0a0a0a0a0a08;
    encBuf[1447] = 256'h0a08090a090a0909090909090a08000809000809090800080900000800010808;
    encBuf[1448] = 256'h0001020100000008010100010200010808000008000000010808000009080808;
    encBuf[1449] = 256'h090809090809090b0a0a0b0b09090a0b0c0b0b0a0c0a0c0b0b0c0c0a0a0b0c0b;
    encBuf[1450] = 256'h0c0b0b0b0a0d0b0b0a0b0c0c0a0a0b0b0d0a0a0b0b0b0a0b0c0a0a08090a090a;
    encBuf[1451] = 256'h0b090a0808000008000000000000000100010202020303010301040303030403;
    encBuf[1452] = 256'h0304020403030502020203030403020502030403020403030502010202020303;
    encBuf[1453] = 256'h0403030303020302020102010103020201000000000101000000090808090a08;
    encBuf[1454] = 256'h0a09090a09080c0a0b0c0a0b0e090a0a0a0b0e0a0b0a0b0b0d0b0b0c0c0a0b0b;
    encBuf[1455] = 256'h0b0c0b0b0d0b0b0c0a0b0c0b0a0c0a0b0b0b0c0b0b0c0b090b0c0a0a0c090b0a;
    encBuf[1456] = 256'h0a0a0a0b0b0a09090b0808000101000100080201020302020502010401020502;
    encBuf[1457] = 256'h0203040303030306020104020303040404010203020202030305030304020202;
    encBuf[1458] = 256'h030304020304010102030203010203020201000001000800000800080808090a;
    encBuf[1459] = 256'h09090a090a0a0a0b0c0a090b0a080b090a090b0b0b0c0a0b0b0b0c0a0b0c0b0c;
    encBuf[1460] = 256'h0b0a0a0c0a0b0c0a0b0b0b0b0c0a0b0a0a090b0909090a0b0a09090a090a0a08;
    encBuf[1461] = 256'h0908000800000801010800020800020201020302040203040202030303050202;
    encBuf[1462] = 256'h0304030403040302020304040303040402030303040402030302030502020302;
    encBuf[1463] = 256'h0403030304020302030502010203040401010302020201010201010000000108;
    encBuf[1464] = 256'h00010801010809080909080808080a080809080a0b09090a0b0a0b090a0b0a0a;
    encBuf[1465] = 256'h0b0a0a0b090a0b0b0b0c0a090a08090b080a0d09090808080a08080a00090a0a;
    encBuf[1466] = 256'h090a080009080100010001020200020100020101020303050302030301030301;
    encBuf[1467] = 256'h0403030602010203040404020303020402030202030504030403020302010203;
    encBuf[1468] = 256'h0104050304030304020202030204020102020203030504040203020800090808;
    encBuf[1469] = 256'h010002010204020204010908000a00080900080b00020801000b090c0d0a0b0b;
    encBuf[1470] = 256'h0b0b0b080a0b0a0c0b0b0d0c0a0b0c0a0c0b0c0a0a0a090b0a0c0c0c0c0c0b0c;
    encBuf[1471] = 256'h0a0a0a090008090a0c0c0b0c0b0a0c09090a09080a0900090b0b0d0a0c0b0c0a;
    encBuf[1472] = 256'h0a0a000801040102000909080908020801020002030203040203010001080a09;
    encBuf[1473] = 256'h000104030205030202020000080003020104020102020103010008090c090b0b;
    encBuf[1474] = 256'h090000020100010b0b0a0a0b08080001000b0b0e0b090a0a01080a090b0c0b0f;
    encBuf[1475] = 256'h0b0a0b0b080909000a0b090b0a090a0b0b0f0b0b0b0b0800010209090a0f0b0c;
    encBuf[1476] = 256'h0b0b0a0a09000909090b090909080100090a0f0b0a0c0a08000002020000090c;
    encBuf[1477] = 256'h0c0d0b0b0b09000002050202020002000b0d0b0f0a090800030403030000090d;
    encBuf[1478] = 256'h0b0b0d0a090800020303040202010b0b0b0e0b0a0d0909090003030402080a0d;
    encBuf[1479] = 256'h0f0b0b0d0a090000020102020800090b0c0c0f0b0a0b08010103030108090e0c;
    encBuf[1480] = 256'h0b0d0a09090002020303010100090b0a0d0a0908020303040200040202050202;
    encBuf[1481] = 256'h0108090001010604040503030304010200080800000306040403030402010101;
    encBuf[1482] = 256'h01000000030404060402040101010008080002030504040202000009090a0800;
    encBuf[1483] = 256'h0205040303030200000809090a000103060502030108090b0d0b0b0c0a090900;
    encBuf[1484] = 256'h000801000808090c0b0d0b0b0b0d0c0b0c090908010100090d0f0c0c0c0a0908;
    encBuf[1485] = 256'h0002030302000a0c0d0c0c0b0a0900020404030200090b0e0c0a0b0a08010204;
    encBuf[1486] = 256'h04020300080a0b0c0a0a0800030503040202010000080000090a0b0d09010207;
    encBuf[1487] = 256'h0503050203020000090b0a0a09010505040403030301080b0d0b0c0908020504;
    encBuf[1488] = 256'h04030301000a0a0c0b0a080102040404020100080a0a0d0b0a0a080003040402;
    encBuf[1489] = 256'h0200090c0b0d0b09090801010009090b0a0a0a00080b0f0e0d0b0c0b08080203;
    encBuf[1490] = 256'h0303010a0f0d0b0b0b080003030302080a0d0d0b0c0a09090000010101000809;
    encBuf[1491] = 256'h0b0c0d0c0a09080205030301080b0e0c0b0a0a08010305020201080a0c0b0b0a;
    encBuf[1492] = 256'h080103030403010102000800090900080801000a08000003050405020200090c;
    encBuf[1493] = 256'h0b0d0b09090107060404030201080c0d0c0b0b0908030604030201090b0d0b0c;
    encBuf[1494] = 256'h0a0901030404030301080a0c0d0b0a0b0808020403040301080a0c0c0b0b0908;
    encBuf[1495] = 256'h020403030208080b0b0b0a080000000b0f0c0b0900030703040200080c0c0b0c;
    encBuf[1496] = 256'h0a090102050304030101080b0d0c0b0b0a08030505040201000a0b0d0b0a0901;
    encBuf[1497] = 256'h030503040200080a0b0b0b0a080103040403020108090b0b0b09010306040302;
    encBuf[1498] = 256'h01000a0b0d0b0a00040505030200090c0d0b0a0801040404030108090c0c0b0a;
    encBuf[1499] = 256'h0801030503020208090a0c0b0a0908010304030302080b0d0c0b0a0901040403;
    encBuf[1500] = 256'h040200090b0d0c0a0900030504020208090d0c0b0b0a00030603040200080a0b;
    encBuf[1501] = 256'h0b0b0a09080103040404020201080b0f0b0d0a0900030405030201090b0d0b0a;
    encBuf[1502] = 256'h0800030304020008090a0a0808010201080a0c0d0a0802060403040108090c0a;
    encBuf[1503] = 256'h0b090900010203030504020300090d0d0c0b0b0902040603040200080a0c0c0a;
    encBuf[1504] = 256'h0a08010304030301000a0c0b0c0a0908010204040202010008090a0a0a0c0b0c;
    encBuf[1505] = 256'h09080205030402080a0b0d0a0a08080102040305020200080b0c0c0b0b0b0a09;
    encBuf[1506] = 256'h08020405030200090c0b0b0a0908010205030401080b0e0b0b0a0908080a0b0c;
    encBuf[1507] = 256'h09000406040200090b0e0b0b0a0800030403040200080b0d0d0b0b0c09090103;
    encBuf[1508] = 256'h0703040208090d0c0b0b08000305030302000a0c0c0c0a0a0000020402030101;
    encBuf[1509] = 256'h08090a0d0b0c0a09000206030303010a0c0d0c0a0a08020305030200080b0c0b;
    encBuf[1510] = 256'h0a090205030401090a0d0b0b09010204030200080b0a0b080003040402020008;
    encBuf[1511] = 256'h0a0b0c0c0b0b0c0b0b09010506030302000a0d0b0c0a08010306040303000b0f;
    encBuf[1512] = 256'h0c0b0c09000204030201000a0b0b0b0a0002030403020009090c0b0b0d0b0b0b;
    encBuf[1513] = 256'h0a09020604030301090a0d0a09080002030101090a0c0c0a0a0802030402000c;
    encBuf[1514] = 256'h0f0c0b0a0802050404020108090b0c0b0b0a0901030504030301080c0d0c0c0a;
    encBuf[1515] = 256'h0900020404030301080a0c0c0a0a0901030403020108090b0c0c0b0a0a080002;
    encBuf[1516] = 256'h0503040202000808090809090a0b0b0c0c0a0a0908020505030302080b0e0c0b;
    encBuf[1517] = 256'h0b09000406040302000a0c0e0b0b090802040303030100090b0b0c0c0a0a0900;
    encBuf[1518] = 256'h020304030300090b0e0b0b0b080003050403020100090b0c0c0b0b0908000201;
    encBuf[1519] = 256'h00090908020706030201090c0c0b0a0004040302080a0d0b0b08020505030200;
    encBuf[1520] = 256'h090b0c0a0a09010204030402010008090900010201000809000406050202000a;
    encBuf[1521] = 256'h0c0b0c0a0a08010204050404020303030201080b0f0d0b0a0901040403030009;
    encBuf[1522] = 256'h0c0d0b0a090203070303020200090b0b0c0b0a090900020203030100090a0b0a;
    encBuf[1523] = 256'h090002050405030403030100080c0c0c0908000201090f0c0c0a000206040302;
    encBuf[1524] = 256'h000a0d0b0b0a010405030301080b0c0c0a0908000203020201000909090a0908;
    encBuf[1525] = 256'h09000104060404020201090a0c0c0b0b0b0a00030604040101080a0b09080305;
    encBuf[1526] = 256'h030301080a0b0a0800030201090d0d0b0b00030704030201010808000100080a;
    encBuf[1527] = 256'h0b0c0a000204030108090909020402010a0d0a0804070703040200090c0c0c0a;
    encBuf[1528] = 256'h0a0800020404020301080a0c0c0a09000305040302080a0c0c0c0a0900020305;
    encBuf[1529] = 256'h020008090b0a09080001020202020404030301090e0c0d0a0b09090000010203;
    encBuf[1530] = 256'h03030402020200080b0d0d0c0b080105050303010a0c0e0c0b0a0a0801040504;
    encBuf[1531] = 256'h020208090c0b0b09000203020100090a09080000090c0d0d0c0a080002060304;
    encBuf[1532] = 256'h0200000a0b0d0a0a0908000203020200080b0d0c0b0a09000102030303040304;
    encBuf[1533] = 256'h02000a0c0f0b0b0a0801020201080c0b0c0b0900010303030502010200010008;
    encBuf[1534] = 256'h0b0d0e0c0c0a0a08000002010808090900010000080a000307070302000a0e0c;
    encBuf[1535] = 256'h0c0a0a09000204030201090a0c0c0a0a0001040504020100090b0d0b0b0a0a0a;
    encBuf[1536] = 256'h09080001040404040301090c0d0d0a08000404030201090b0d0b0b0a08080101;
    encBuf[1537] = 256'h03020201000a0a0b0900030303010809090105050402080d0e0d0c0b0a080203;
    encBuf[1538] = 256'h0602020100090a0a0a00010201090d0c0b090106030401090b0e0b0c09080203;
    encBuf[1539] = 256'h0404030200090c0c0a0a080002030200080a0b0c0a09080305050201080a0c0b;
    encBuf[1540] = 256'h0a0003060301000a0c0b0a09010201080b0e0b09000306040201000a0b0b0a0a;
    encBuf[1541] = 256'h00020403030202010a0d0d0c0b0a0002040302000a0d0b0a010605040201090b;
    encBuf[1542] = 256'h0e0b0909000201020100000800080101020301080b0f0a0a010506040302080b;
    encBuf[1543] = 256'h0e0c0c0a09080103040402010008090a090001030301000b0e0c0a0a08010202;
    encBuf[1544] = 256'h00080c0b0c09080205040504030302080a0c0d0a0a0808010101010008090a0b;
    encBuf[1545] = 256'h0c0a0901020504030403040303000a0f0b0c0a0801030303000a0d0b0a090204;
    encBuf[1546] = 256'h040302010009090808010108090b0e0c0b0a09080102040302080a0b0a000104;
    encBuf[1547] = 256'h0403050406030402080a0d0c0c0b0a0a0800030504030301000a0b0c0b090002;
    encBuf[1548] = 256'h03030301090b0d0b090000080a0d0d0b0a010407030402000009090a08080801;
    encBuf[1549] = 256'h0808090b0c0a0908020504030301000c0c0c0b09000306040301000b0c0b0b08;
    encBuf[1550] = 256'h0002030208090a0b0804070703030200090c0b0c0a090001030204020201090b;
    encBuf[1551] = 256'h0f0c0b0a09080103020303040504030301080a0d0c0a0b090001020303020200;
    encBuf[1552] = 256'h00080a0c0d0b0a00020503030303040402010a0e0d0b0a090908090b0a080106;
    encBuf[1553] = 256'h040303000808000204040201090c0a0901050402010a0d0d0c0a0a0800030304;
    encBuf[1554] = 256'h0201000808080808080808090a0d0d0b0b0803060403020809090a0802050404;
    encBuf[1555] = 256'h0302000a0b0c0d0a0a080908080a0c0b0b080307050402010008090909080909;
    encBuf[1556] = 256'h090b0b0c0b0a0a0003050503030201080b0a0a000506030402000909090a0b0e;
    encBuf[1557] = 256'h0d0b0c0b0a090001020203040402020108090a090106040302000b0c0c0a0900;
    encBuf[1558] = 256'h00000a0d0c0b0a010307030201080a0b0a0a080000080a0b0e0c0a0a08010304;
    encBuf[1559] = 256'h0300090b0c0901050504020201080809080000080a0f0c0d0c0b0a0a00030604;
    encBuf[1560] = 256'h030200090b0c0b0a0800010108090b0a0805050403000a0e0b0c0a0801020304;
    encBuf[1561] = 256'h04040201080a0b0c0b09090808000800080101000108090c0d0b0b0a00080000;
    encBuf[1562] = 256'h09010406040201080d0b0c0a00020503030108090908010202000d0d0c0a0a09;
    encBuf[1563] = 256'h08090a09090808090b0d0b0a030707030301000a0b0c0c0a090001020301000b;
    encBuf[1564] = 256'h0c0c0b0802050402080a0d0c0a0802040304020009090b0a0a0909090c0c0a09;
    encBuf[1565] = 256'h010302090f0f0a0908020401010101020604030200090d0c0b0b0a0808000008;
    encBuf[1566] = 256'h080002030303080a0c0b0b0a0c0c0c09000506040302000a0b0d0a0808000101;
    encBuf[1567] = 256'h010103040300090c0c0a09080a0c0e0c0a08010204030008080801030403080a;
    encBuf[1568] = 256'h0d0b0801050302080c0d0a0a0002030208090a0801020202010306040302090c;
    encBuf[1569] = 256'h0d0b0b08010302010b0f0b0b09020402090e0d0a0004050302000a0b0b090001;
    encBuf[1570] = 256'h0102020305050202080b0d0b0b090800090b0b0a020704030200090b0a080001;
    encBuf[1571] = 256'h00000008080801020404010a0e0d0c0b090802030504040202020009090b0b0b;
    encBuf[1572] = 256'h0d0c0b0b08030704020200080808000101080a0d0c0b0c09090001030300090c;
    encBuf[1573] = 256'h0b0b0004040302030504050302020808090808080b0d0d0b0b0a090808080002;
    encBuf[1574] = 256'h0203040403040301090d0d0c0a090102040304020204040202080c0c0b0b0908;
    encBuf[1575] = 256'h08080909020406030300080a0a0a0b0b0c0b080206040200080a0a0a00080202;
    encBuf[1576] = 256'h050503040201000800090a0d0e0b0c0b0a090908010307050303030202000809;
    encBuf[1577] = 256'h0a0b0c0b0b0d0b0d0a090801020202000001020504040403030201090c0c0a0a;
    encBuf[1578] = 256'h0808090c0d0c0a0908010102020305040403020208090b0d0b0b0a0002040201;
    encBuf[1579] = 256'h090b0b0802070301090b0d0a080404040100090909080a0d0d0d0a0900020302;
    encBuf[1580] = 256'h010100020504020100090908000002000a0c0d0c0c0a0a090102030503030301;
    encBuf[1581] = 256'h000a0a0b0a0103050200090c0b0c0b0b0d0c0b0a090205040401000b0c0c0a00;
    encBuf[1582] = 256'h020303000a0d0b0a00020200090007070703030301080b0c0d0b0b0b0a090001;
    encBuf[1583] = 256'h04020201090c0b0d0909000303040303040200090b0d0b0a0800000000080102;
    encBuf[1584] = 256'h050302020101010108090809080b0f0e0c0a0a00030402080b0f0a0900020302;
    encBuf[1585] = 256'h080b0d0a08010201080a0c0a09000200090c0a00060704030401010809090a0a;
    encBuf[1586] = 256'h0a0b0b0b0909080001080a0c0c0a0002040302080a0b09080c0d0d0b08040503;
    encBuf[1587] = 256'h01080b0e0c0b0b0a09010306030303020203010a0f0d0b090205050302000909;
    encBuf[1588] = 256'h0a0b0a0c0c0a0a0003040301090c0c0b0b0a0a0800020405030201080a0b0b08;
    encBuf[1589] = 256'h0103040201090b0b0804070503020108090b0b0c0b0c0b0b0902040503020809;
    encBuf[1590] = 256'h0d0b0b0b0a0909000002020200090b0a0003070402000a0c0a08030706030200;
    encBuf[1591] = 256'h090c0d0b0b0a09080104050403020208080a0b0c0d0b0c0a0802030602010009;
    encBuf[1592] = 256'h0a0a0808000001010008090c0c0b0c0b0a0a0900020405030304020303020208;
    encBuf[1593] = 256'h0a0b0b01050502000a0e0b0b0b0a0b0909000206030303020101000a0d0d0b0c;
    encBuf[1594] = 256'h0a0a0a0a0a09080204020302040505040301080908000203000a0f0b0a080101;
    encBuf[1595] = 256'h000b0d0a08020301080a0a0307050200090b0b0908090b0e0c0b080203040200;
    encBuf[1596] = 256'h08000204040301000008080a0e0c0c09000405030200090a0b0b090908090a09;
    encBuf[1597] = 256'h0803070303000a0e0b0a00030402020008080808090b0b0b0a0b0c0e0c0b0901;
    encBuf[1598] = 256'h070503030200000909090808080100000809090005050302090d0d0b0b0b0a0c;
    encBuf[1599] = 256'h0a0b0901030504030404030402010008010201000d0e0d0a0a09000101010008;
    encBuf[1600] = 256'h080002040504020200090c0b0a0900010008090b0a0a0a0a0c0b090207060304;
    encBuf[1601] = 256'h02030302000a0e0d0c0a0a000102020100010101020100090a000102000a0d0b;
    encBuf[1602] = 256'h090101080f0d0b0b080102020203060403020201030504030301090c0d0d0b0d;
    encBuf[1603] = 256'h0a0a08000100010000020504030402010008090a0a0b0a0a0a0a0a0c0b0a0207;
    encBuf[1604] = 256'h050302000a0b0c0a0a09000002040402020809090808090d0d0c090205040401;
    encBuf[1605] = 256'h08090908010203000a0d0b0c090909090a08080100080c0b0905070504010008;
    encBuf[1606] = 256'h0b0b0a0808010008080a0801030405030201090a0c0c0b0b0a0a0a0900030603;
    encBuf[1607] = 256'h020101020605040202080c0c0d0b0b0a0801030403020109090a090900000306;
    encBuf[1608] = 256'h04040201090b0e0b0a0900000108090b0b0b090105050403030403030200080c;
    encBuf[1609] = 256'h0e0d0b0b0b0900020304020008080a0a0a0a08030706030200090c0b0a0a0800;
    encBuf[1610] = 256'h0000000000000900010307040200090c0b0a09010300090c0e0a0a0002030200;
    encBuf[1611] = 256'h0a0c0d0a0a0a08000106050504030200090b0d0b0b0a0a090909010205040402;
    encBuf[1612] = 256'h02020008080008090a0d0c0c0b0b09000800000a0a0c0a090104050503040301;
    encBuf[1613] = 256'h0008080a0a0a0a0a0a09000202010a0f0f0b0c09000204030301010800090b0e;
    encBuf[1614] = 256'h0c0c09080204030300090b0b0b08010305030301090d0c0c0b09080102040202;
    encBuf[1615] = 256'h0008090b0b0a0002050403030000090a0b0d0e0c0b0b0b08020405030301080a;
    encBuf[1616] = 256'h0a090800010100020201000a0e0b09020503000b0e0b0b09090b0e0c09000404;
    encBuf[1617] = 256'h0302000808020302090f0c0c0900010101000801030301090e0c0a000103010b;
    encBuf[1618] = 256'h0e0c0b09010102030205050302010a0c0c0a0900010201010000090d0d0c0a00;
    encBuf[1619] = 256'h02040201080a09000204040303020200090f0d0c0a0a0908090a0c0a08020705;
    encBuf[1620] = 256'h03030101000008080a0a0c0a0b090a090a09080001010108080809080a0a0901;
    encBuf[1621] = 256'h07070302010909090908080a0c0b000606040302080a0c0b0a0a0a0b0b0b0a08;
    encBuf[1622] = 256'h01030203020304030203050406030301090b0c0a0a090c0e0c0b090104040200;
    encBuf[1623] = 256'h08090801040200090a0a00030503020808090a0b0d0c0b0003070402000a0c0b;
    encBuf[1624] = 256'h0a08010201000a0b0c0a090102030302080b0901070402000b0e0b0902040402;
    encBuf[1625] = 256'h0100000104040301000a0d0c0d0b0c0909010102010101020404030202000008;
    encBuf[1626] = 256'h0d0d0d0b09000306030108090a0a0a09080a0a0800020300090a000706040301;
    encBuf[1627] = 256'h0009090900000202020303000c0e0d0c0b0b0a0b090801050405020100080000;
    encBuf[1628] = 256'h020301080c0b0900040401090c0c09080000090d0b0a02060502010809090800;
    encBuf[1629] = 256'h00080b0d0b0a08010304030101080b0b0d0a080305050302010008090a0c0c0c;
    encBuf[1630] = 256'h0b0b080002040203020404050302000a0b0d0b0a0b0a0908010404030200090a;
    encBuf[1631] = 256'h0a090908000307060302080d0d0c0a0800030302010000080102030403020108;
    encBuf[1632] = 256'h0c0d0b0c0a090a0a0a09010605030401000808090a0c0b0c0900020403010008;
    encBuf[1633] = 256'h08020502000a0d0b0a000101090c0e0a0003050401000909090809090b0c0a08;
    encBuf[1634] = 256'h010304020203050301000b0d0a080101080d0e0c0a0802030503010008080103;
    encBuf[1635] = 256'h030400090c0c0a0a0800000008080909090b0e0b0d0a09000307050403030101;
    encBuf[1636] = 256'h090a0b0b0b0c0b0c0a0900020402020009090b0b0c0c0a080004050303030202;
    encBuf[1637] = 256'h01090b0e0d0a09000100080800030707020100090b09090800090a0d0b0a0908;
    encBuf[1638] = 256'h010008090a090900020604030301090b0c0901030302080a0801040400080002;
    encBuf[1639] = 256'h07070301090d0d0c09090002020201010200010108090b0c0c0a0a0a0a0b0c0b;
    encBuf[1640] = 256'h0902050402010a0b0b0a0103050305040404040301000a0d0c0c0b0c0a0a0908;
    encBuf[1641] = 256'h020305040200000909090809090a0b0a080103040203030302090c0d0c090001;
    encBuf[1642] = 256'h00090c0d0a0002050201080a09090000090b0e0c0a0908010404030301000808;
    encBuf[1643] = 256'h080100090b0a0a0002090f0f0e0a09000103020201090a0d0b0b0a0900020404;
    encBuf[1644] = 256'h0504030301080d0d0c0b0b0a080000020303030303050304020008090b0b0a08;
    encBuf[1645] = 256'h080a0d0b0c09080101000c0f0d0c0a09090002000100010306030300080a0901;
    encBuf[1646] = 256'h030401090d0b0a000306030200090b0b0c0b0a0b0c0a0a08030705030301090c;
    encBuf[1647] = 256'h0c0b0b09080009090a09090800080808000505050403030200080a0b0d0a0909;
    encBuf[1648] = 256'h000108010002040502010b0e0c0b0b0909090c0b0c09010306030200080a0a0b;
    encBuf[1649] = 256'h0b09080103050404030503030402010109090c0c0c0c0c0b0b09090103040302;
    encBuf[1650] = 256'h01080a0a0c0a0a08000002040405030401000a0a0a0003040300090c0c0a0908;
    encBuf[1651] = 256'h080000040504040108090c0c0a0a0a0a0a090800000100020606050402010809;
    encBuf[1652] = 256'h0a0a0a0a090a0b0a0a090102050504040302020809090b0b0d0b0e0a0a090101;
    encBuf[1653] = 256'h000008080003070304010100000000000a0c0c0b090901040304020108000801;
    encBuf[1654] = 256'h030201090e0d0b0a08000101090b0d0c0a090204060303030302020101000b0e;
    encBuf[1655] = 256'h0c0a09000008090d0c0b0901030702020100080104040301080b0d0c09090008;
    encBuf[1656] = 256'h090b0c0b0908010102040604030403020000080a0c0c0c0a0a08000202040304;
    encBuf[1657] = 256'h0201090c0c0b0b0b0a0a0a090804060402010809080808000808090002030401;
    encBuf[1658] = 256'h0100030603030108090800000c0f0d0b0b08000202030604040402010008080a;
    encBuf[1659] = 256'h0a0b0e0b0b0a00010200090b0a020705030200090908010202080b0e0c0b0a09;
    encBuf[1660] = 256'h000101020202010100000304050302030306040303080c0e0c0b0a0a09090a0b;
    encBuf[1661] = 256'h090004060503030100090b0a0a090001010100090a0b0c0b0e0b0c0a08020705;
    encBuf[1662] = 256'h03040101080808080000080a0a0c0a0b090800020405030201000b0c0b0c0900;
    encBuf[1663] = 256'h02040301000a0902060503020008090b090a0b09080205030303030406040202;
    encBuf[1664] = 256'h090c0b0c0b0b0b0d0b0a0902050303030001020306030302010a0c0d0b0c0b0c;
    encBuf[1665] = 256'h0a0a090908000102030505040404020008090a0a0808090b0e0b0b0a00000100;
    encBuf[1666] = 256'h080105050402080a0d0d0b0a0a0908090000000202030203020100090b0f0d0c;
    encBuf[1667] = 256'h0b0b0a0900010202080a0c0d0a0908010201080000020306020108090a0b0c0c;
    encBuf[1668] = 256'h0b0a0b090a0e0d0b0a000606030301080b0c0b0c0a0b0a090801020203030301;
    encBuf[1669] = 256'h00080808010406040301090d0c0b0a0002050302080b0f0d0a0b0a0a08080001;
    encBuf[1670] = 256'h030405030302020200000a0c0d0c0a0a080008000a0a09080206030302000a0a;
    encBuf[1671] = 256'h0c0c0c0b0c0a0a08080100010103050301080c0c0a0901030300080803070602;
    encBuf[1672] = 256'h000b0c0c0a090008090801050604030300090a0b0c0c0b0c0a09080808090909;
    encBuf[1673] = 256'h0204050302000808010305020302010102000a0d0d0b0b0a0001030502010009;
    encBuf[1674] = 256'h0c09000307030201080908000201080908010706030201080a09080205050504;
    encBuf[1675] = 256'h040202010108090809080100010202020203050503030301080800000202000a;
    encBuf[1676] = 256'h0d0c0b0a0a0b0c0c0b0b00030704030201080b0c0a0a09080a0e0c0e0b0b0c0a;
    encBuf[1677] = 256'h0909000000000809090808080c0d0d0c0a0b0a0b0a0b0b08010203010b0e0c0b;
    encBuf[1678] = 256'h0b09090a0c0a0a090000090b0d0a0902040402010102020402080b0f0b0b0802;
    encBuf[1679] = 256'h0404020302020305020302020101020604030403010202010001080102050505;
    encBuf[1680] = 256'h0202020100080b0c0a0902050402080a0c0a0a0008090d0d0c0a090800000009;
    encBuf[1681] = 256'h080b0b0b0c0b080102060202000a0d0c0c0b0b0b0a080908080a0d0b0b0a0002;
    encBuf[1682] = 256'h0305020001000101080d0e0e0c0b0a0900000202010205040503030201080a0a;
    encBuf[1683] = 256'h0d0b0c0c09080202040101000002040402020000010000090e0d0b0b09080001;
    encBuf[1684] = 256'h0001010405040304020100090b0c0d0b0b0c0a0a0a09090a0c0b0b0b08020304;
    encBuf[1685] = 256'h030203070505040304030302020100080a090a09080103040303030100000000;
    encBuf[1686] = 256'h090b0f0c0a000307030402010103030502000809090800010001010305040401;
    encBuf[1687] = 256'h01080809090a0b0b0a0804050202080908080202000c0f0c0c0a0b0b0d0c0c0b;
    encBuf[1688] = 256'h0b0a0a090a0a0b0b0d0a0b0a0b0b0a0901040402020a0c0c0d0b0b0d0c0a0b0b;
    encBuf[1689] = 256'h0909090000000203040304030304020300080a0b090005040403030101010002;
    encBuf[1690] = 256'h0000010307060305030303030403030403040303040201020000000809080001;
    encBuf[1691] = 256'h0201000a0c0b090002000b0d0a08040602000c0e0c0b09080808000909090b0c;
    encBuf[1692] = 256'h0c0d0c0b0b0b0a0b0d0c0b0c0909000808090b0d0b0b0b09090b0a0c0c0b0b0b;
    encBuf[1693] = 256'h0a0a0b0a0c0d0b0c0b0b0a08020203010109000103050100090c0a0a09000001;
    encBuf[1694] = 256'h0305050505030404020101090809000102020202000205060404020302000908;
    encBuf[1695] = 256'h0908020306030201080b0d0c0b0b090908090a0d0b0b0a0909090b0d0b090002;
    encBuf[1696] = 256'h0502080a0d0d0c0b0c0b0b0a090800010100010100010a0c0c0c0c0a0a0a0b0b;
    encBuf[1697] = 256'h0c090908010103040403040100000c0c0d0c0c0a090802040201080a0b0a0908;
    encBuf[1698] = 256'h090a0d0c0b0b0c0b0d0c0b090105040503030304040403050304020201010000;
    encBuf[1699] = 256'h00000203020101080a0b0d0c0b0b0a0800010404040404030304030303030301;
    encBuf[1700] = 256'h080a090a090800000205040403030302010008090d0d0b0c0900010304020108;
    encBuf[1701] = 256'h080b0a0c0c0c0c0d0b0c0b0b0c0b0a0b0b0a0b0c0b0d0b0c0b0b0a0b0b0b0a09;
    encBuf[1702] = 256'h090001020201020200090d0e0d0b0c0b0b0b0c0a0a0909090800020404030402;
    encBuf[1703] = 256'h0102030504030302020202020202020305030502030403040403040303030502;
    encBuf[1704] = 256'h0302020001000103060404040203020202020108090a0a0b090909090a0c0b0c;
    encBuf[1705] = 256'h0a080001030200090c0d0b0c0b0d0d0c0b0c0b0a0a0c0c0c0b0b0c0a0a0a0a09;
    encBuf[1706] = 256'h0a090008010008090b0d0c0c0a0b0a0b0c0c0c0b0c0a09090008000808080002;
    encBuf[1707] = 256'h030402010a0b0d0b0b0b0b0b0d0a0a080105060404020302000101020202000b;
    encBuf[1708] = 256'h0d0e0b0a0908000001020304050303030202040202030102000a0b0c0c0b0c0c;
    encBuf[1709] = 256'h0c0b0c0b0a0b090a0b0a0a080002010202020305000b0f0f0b0b0b0c0a090801;
    encBuf[1710] = 256'h0404040100090a08000305040202000008080a0b0b0e0b0c0b0a080003050304;
    encBuf[1711] = 256'h03030404020200090b0c0b00010301090f0d0b09080204030403040303010109;
    encBuf[1712] = 256'h0a0a0a0001000a0e0d0b0a0a08000100080a0c0c0b09090800080a0c0c0c0a0c;
    encBuf[1713] = 256'h0a0909090a0d0b0b0a0307070703030402020202020201010002010403020301;
    encBuf[1714] = 256'h0809090a09080800010908020507060303020201020202030303030405030203;
    encBuf[1715] = 256'h030203030302090d0c0d0b0b0c0b0a0a09000800090a0b0c0b0b0b0b0c0b0e0d;
    encBuf[1716] = 256'h0b0e0b0b0c0a090a090a0b0b0c0d0b0b0c0b0d0b0c0b0c0a0a0909090808090a;
    encBuf[1717] = 256'h0a0b0b0a0a09090809090a0c0c0a0a0a0801000000090a0a0903070704040201;
    encBuf[1718] = 256'h0101010305040404020302020202030505040303030402020201010200020202;
    encBuf[1719] = 256'h0303030405040304030202010101010009090a0a09080008090b0c0b0a0a090e;
    encBuf[1720] = 256'h0e0d0d0b0c0b0b090a0a0a0c0b0c0c0a0b0b0b0b0c0a0b0a0a0808010200090d;
    encBuf[1721] = 256'h0f0c0c0a0b090b090b0a0909090a0a0c0a0b080001020100000809090a0a0003;
    encBuf[1722] = 256'h0707040202020100000002020406030403020008080001050405030302020008;
    encBuf[1723] = 256'h000002030303030305030301080a0b0909090a0f0b0901040502090e0d0b0b0a;
    encBuf[1724] = 256'h0a080808080a0a0b0c0a090102020b0f0f0c0b0b0a0b0a0a09090000080a0c0c;
    encBuf[1725] = 256'h0b0b0a0b0c0c0c0a000003030201000102020100080d0b0b0a08020404050108;
    encBuf[1726] = 256'h090d0c0a0a08030304030302030304040100080d0b0a0a02050504030201080a;
    encBuf[1727] = 256'h0909000002080a0c0d0a0a0908080b0d0e0c0c0b0a0a0809090a0b0c0c0b0c0a;
    encBuf[1728] = 256'h0a0a080102040403050404050403050303040202020101000101020303030301;
    encBuf[1729] = 256'h00090b0d0c0a0a08010203060403040403040203030203040303050304030304;
    encBuf[1730] = 256'h030303010108090c0a0c0b0b0b0b0c0a0c0b0c0b0b0b0a0a0b0c0b0c0a0b0d0b;
    encBuf[1731] = 256'h0d0c0a0a0a090a090b0c0e0b0d0c0b0b0c0a0a0a0a090a090a0a0b0b0c0a0a0a;
    encBuf[1732] = 256'h0a0a0a0b0b0a0a0b0c0c0b0b0901040603030201000909080001030402040404;
    encBuf[1733] = 256'h0503040201010204050503030304030404020303030304030603030402010201;
    encBuf[1734] = 256'h010101010000080001030302010009090102070303030303040302000a0e0d0b;
    encBuf[1735] = 256'h0c0a0a090a0a0b0a0c0c0c0d0d0b0b0c0b0b0a0a0b0a090b0a0b0b0b0b0a0a0b;
    encBuf[1736] = 256'h0d0b0b0b0c0a0c0b0d0b0c0a0b0a0a0b090a0b0b0c0c0b0b0b0a080203030302;
    encBuf[1737] = 256'h09090b0b0a0b0c0a000407070403040102020304030302000800010505040203;
    encBuf[1738] = 256'h0101010002020404040302030101020201080b0e0b090004050201090b0e0a0b;
    encBuf[1739] = 256'h0b0b0c0c0a0b0909000100080b0e0c0b0b0a0808000000020201080c0d0c0c09;
    encBuf[1740] = 256'h0a08080809090c0d0b0a09000203030208000800080c0f0b0d0a0909090b0e0c;
    encBuf[1741] = 256'h0a0a0002040403030303020201080a080004060402020808090a0a0909090809;
    encBuf[1742] = 256'h08010000080e0d0b0b0a080000090d0c0c0b0909090a0f0c0b0b0b0a0a090002;
    encBuf[1743] = 256'h04070405040403050302040202020101010002020403030100090b0b0a0b0b09;
    encBuf[1744] = 256'h0a00030704030303030305040404040203030304030304040203030202000809;
    encBuf[1745] = 256'h0b0d0c0c0b0b0a090808080a0b0c0c0b0b0c0b0b0b0b0b0b0e0b0c0c0a0a0a0a;
    encBuf[1746] = 256'h090a0b0c0d0b0d0c0b0b0d0b0b0b0a0a0a0a0a0b0c0b0b0a0a090809080a0a0a;
    encBuf[1747] = 256'h0b09090801030605050303030100000800010202030202030404060304050204;
    encBuf[1748] = 256'h030305040303030403040405030304020302020102010101030203040100080a;
    encBuf[1749] = 256'h0908000103030403010208090c0c0c0b090900010101080d0c0d0c0a0b0b0a0c;
    encBuf[1750] = 256'h0c0b0c0a0a0b0d0b0e0b0c0b0b0a0c0b0a0b0a0b0c0c0c0c0b0b0a0908080909;
    encBuf[1751] = 256'h0a0a0a0908000108080b0b0e0b0b0a090908090a0b0b0c0b0e0c0d0b0b0c0908;
    encBuf[1752] = 256'h0002020304050403030302030203030201000a0b0a0804070404030304020201;
    encBuf[1753] = 256'h00080909090908000801010405040304020202020203000a0c0f0c0c0b0b0c0a;
    encBuf[1754] = 256'h0a090809000909080a0a0c0d0c0c0b0a08080001000008090a0a0a0003070403;
    encBuf[1755] = 256'h01080a0e0b0b0b0b090a0a080a08090a0c0b0e0b0b0b0b000003070203020008;
    encBuf[1756] = 256'h010104050301010a0a0000050400080b0e0a0808020201080008030604040402;
    encBuf[1757] = 256'h0100080a0b0b0a0001050301090d0e0b0b0b0800010305030603040304030503;
    encBuf[1758] = 256'h06030403020202020001020204040304030202000008090b0b0c0b0a0a080002;
    encBuf[1759] = 256'h02050403060403040303040202010100010103050503030401010008090b0c0b;
    encBuf[1760] = 256'h0b0c0b0c0b0c0b0b0a0b0b0b0d0a0a0b0b0d0c0b0c0b0b0b0b0c0b0b0a0b0b0c;
    encBuf[1761] = 256'h0c0c0b0b0c0a0b0a0b0c0b0b0a0c0b0d0b0c0c0b0a0b0a0a0a0a080900000102;
    encBuf[1762] = 256'h0404030402010100000000010103060504040303030203020303050403040303;
    encBuf[1763] = 256'h0303020402030504040404030402020303030403030303020303020200090b0f;
    encBuf[1764] = 256'h0c0a0b09090a0a0b0b0c0a090808000100010208080a0c0c0b0c0c0b0c0b0c0c;
    encBuf[1765] = 256'h0d0b0d0b0a0a0a0a0c0b0c0b0b0b0c0b0d0b0c0b0b0b0c0c0b0b0c0a08090800;
    encBuf[1766] = 256'h000001010201000000000009090a0b0c0b0c0b0b0a0b0b0e0c0b0a0802020202;
    encBuf[1767] = 256'h0908010307040305040404030304030204040303040203030302000809090900;
    encBuf[1768] = 256'h010203030405040304020201000008080a09090b0b0d0b0a0803070603030201;
    encBuf[1769] = 256'h08090a0c0b0e0b0b0c0b0b0b0b0c0c0a0b0b090909080809090a090004050405;
    encBuf[1770] = 256'h0304020301010008090c0c0c0a0a0801010200090b0d0c0a0b0b0c0b0c0b0c0a;
    encBuf[1771] = 256'h090a09090909010206040404020302020203040303020200080808090b0d0c0b;
    encBuf[1772] = 256'h0a0a0a0d0d0c0b0908010100000808010303010b0f0c0b000506060403040403;
    encBuf[1773] = 256'h03030304020101020002020303030100080a0b0c0b0b0a0a0000010404030504;
    encBuf[1774] = 256'h03030403040304040302030302020404060403030302010008090b0d0b0c0b0b;
    encBuf[1775] = 256'h0c0a0a0a0b0a0c0c0c0b0d0b0b0b0b0b0b0b0c0b0909080008090a0c0b0d0b0d;
    encBuf[1776] = 256'h0b0c0b0b0b0c0b0b0d0a0b0a0b0b0c0c0b0b0c0a0a0a090909090a0b0b0a0a09;
    encBuf[1777] = 256'h0802040404040405030503030202010100010000000002040404040202030303;
    encBuf[1778] = 256'h0502040304040403050203030203030303020304030304030303020202020008;
    encBuf[1779] = 256'h08090b0b0c0d0c0d0b0c0b0b0b0b0b09090900090808080001090a0c0d0a0a09;
    encBuf[1780] = 256'h09090b0e0c0e0b0d0c0b0c0c0b0b0d0a0a0b0a0a0b0c0c0b0a0b0a0b0b0b0b0b;
    encBuf[1781] = 256'h0a0900080100010203010100000001020301080d0f0e0b0c0a0b0a0909080801;
    encBuf[1782] = 256'h0102020101030204050404040306040303050203020303030304030303030201;
    encBuf[1783] = 256'h01000102020402000b0f0d0c0a0b0a090909090a0a0a0b0a090b090808010202;
    encBuf[1784] = 256'h010108080303020400000201080a0f0f0f0f0a0b0a0a0b0a0b0b0b0c0b0d0a0a;
    encBuf[1785] = 256'h0a09090a08000003040202010801030304040009090d0d0b0d0b0a0a08010203;
    encBuf[1786] = 256'h030100010a0a0b0f0f0a0c0b0a0b0a0808010303040402050403050202020100;
    encBuf[1787] = 256'h00010000080b0d0d0c0a0b0a0909090800090009080001030604030504050404;
    encBuf[1788] = 256'h040402030202030303040304030304020202020100000809080809090a0c0b0b;
    encBuf[1789] = 256'h0b09000103060404040304020303040503050304030303020201010808090908;
    encBuf[1790] = 256'h090a0c0e0c0c0b0d0b0b0b0b0c0b0c0b0b0c0b0c0a0a0a090909000908080a0b;
    encBuf[1791] = 256'h0b0c0b0a0c0b0b0d0a0a0b0a0a0c0c0b0e0b0c0c0b0b0c0b0a0b0a0b0a090801;
    encBuf[1792] = 256'h0102020304030504030303050303060303050303030402010201020103030202;
    encBuf[1793] = 256'h0201000101040604040403030404030303030402020304030402030402020200;
    encBuf[1794] = 256'h00000808090809090b0b0e0b0c0b0b0b0b0d0c0c0b0b0b0a09090b0b0c0b0b0a;
    encBuf[1795] = 256'h0a090b0b0c0d0a0b0c0c0b0c0c0a0c0b0c0b0b0c0c0b0b0c0b0c0b0b0d0b0b0b;
    encBuf[1796] = 256'h0b0c0a0b0b0b0a0a090001010304040305030203020100000008010103040404;
    encBuf[1797] = 256'h03040203020108090b0d0b0c0b09000305050403040303040403050203030303;
    encBuf[1798] = 256'h030304020201010000000908090a09090c0b0e0b0c0b0b0b0d0b0c0c0b0a0b0b;
    encBuf[1799] = 256'h0b0a09080101000100080001040402080a0f0d0a0b09000800090a0b0c0d0b0d;
    encBuf[1800] = 256'h0c0c0b0b0b0b0a0a0b0b0c0a0a09090a0908090001020101090b0b0b02070706;
    encBuf[1801] = 256'h030203030202020100090b0b0c0c0b0a0b0a000003050108090b080405050401;
    encBuf[1802] = 256'h00010102040304020102020204020108090a0c0c0c0b0d0a0b0a080103070504;
    encBuf[1803] = 256'h0405030304020303010302020304030502030302020100080900080102020208;
    encBuf[1804] = 256'h0a0d0b0e0a090801030406030202010101030505050303030302010002010102;
    encBuf[1805] = 256'h0100090b0d0c0d0c0b0d0b0b0b0d0b0b0d0b0b0c0a0b0c0b0b0a0b0a0a0a0a0a;
    encBuf[1806] = 256'h0a0b0a0908010208090d0d0c0b0c0b0b0b0c0b0b0b0b0c0b0b0d0c0b0b0b0c0a;
    encBuf[1807] = 256'h0b0b0a0909000000000002050505030403030404040304040203020303040102;
    encBuf[1808] = 256'h0100000000010203050305030304030203030404030502030202020203030303;
    encBuf[1809] = 256'h0403030303020201080a0c0d0b0d0c0b0d0b0b0c0b0b0b0b0c0a0a0a090a0b0d;
    encBuf[1810] = 256'h0c0c0b0c0a0b0a0b0a0b0b0c0b0b0d0b0a0a0a0b0b0c0c0b0b0b0c0a0c0b0d0b;
    encBuf[1811] = 256'h0c0b0b0c0b0b0c0a0b0b0b0b0b0b090901020404030402030203010202030604;
    encBuf[1812] = 256'h0404030303030203020303040201010800080002050205020303050204020303;
    encBuf[1813] = 256'h0403050403030403040303040202010108080808090b0c0d0b0c0b0a0b0a0b0c;
    encBuf[1814] = 256'h0b0b0d0b0b0b0b0b0c0b0b0a09000203070202010009090b0a09090b0b0f0d0b;
    encBuf[1815] = 256'h0d0b0b0b0a0a0b0c0b0d0b0b0b0b0b0c0b0b0c0a090908000001030404050203;
    encBuf[1816] = 256'h03030203020101000801080205030704030403030303000100090a0a0d0b0c0d;
    encBuf[1817] = 256'h0b0b0b0a08010404040303030202020108090b0c0b0901050703030303020603;
    encBuf[1818] = 256'h0604040304030305020302010102020305030503020303020202010101000203;
    encBuf[1819] = 256'h0304020108090b0b0a0b01010101020903070506040404040304030302020101;
    encBuf[1820] = 256'h00080809090a0a0a0b0d0c0d0b0d0b0b0c0b0b0c0c0b0c0b0c0b0b0b0b0b0c0a;
    encBuf[1821] = 256'h0b0b0b0c0b0b0b0b090a090a0a0c0a0c0b0c0b0d0b0c0b0a0a0b0a0c0b0c0c0b;
    encBuf[1822] = 256'h0b0b0c0a09090908080800000002030404040403050304040304030304040304;
    encBuf[1823] = 256'h0303040303020303030202030304040403040304020302020303040302030402;
    encBuf[1824] = 256'h0202010203030504020202000809090a0a0c0c0c0c0b0c0c0b0b0c0a0c0a0b0b;
    encBuf[1825] = 256'h0a0b0b0b0b0c0b0c0c0c0b0c0b0b0c0b0a0b0b0c0c0a0a0b0a0a0b0b0d0b0c0a;
    encBuf[1826] = 256'h0c0a0b0c0b0b0c0b0a0b0a0b0a0a0b0b0c0b0b0b0b0800030504020201020305;
    encBuf[1827] = 256'h0604040403030402030102000001000202030303040304040303040304020202;
    encBuf[1828] = 256'h010202020202020104040503040203020303040202000800080101000b0f0e0c;
    encBuf[1829] = 256'h0b0c0b0a0b0b0b0b0b0d0a0a0b0b0b0d0b0c0b0c0b0c0b0c0a0a0a0a09090808;
    encBuf[1830] = 256'h0908090b0c0b0b0c0a0b0c0b0e0c0b0d0b0a0b0b0a0908000008080b0c0b0d0c;
    encBuf[1831] = 256'h0a0a0a0800010302040303020502040302030502050303030302030303050201;
    encBuf[1832] = 256'h010809090909010404040402020101000008090a09000102010a0c0c0c090202;
    encBuf[1833] = 256'h0706030604030305030404040403030403030203020402040203020302010101;
    encBuf[1834] = 256'h00080808000108080a0d0b0b0b0b0b0c09080106040204010202030405030504;
    encBuf[1835] = 256'h030304020202020203030200090c0b0e0c0b0c0c0b0c0b0c0c0a0c0b0b0c0b0b;
    encBuf[1836] = 256'h0b0c0a0a0b0a0b0b0a0b0c0b0b0b0a0a090808090a0a0c0b0b0b0a0b0b0d0b0c;
    encBuf[1837] = 256'h0c0b0d0c0b0d0a0a090908090a0a0b0908000000010306060304030404030404;
    encBuf[1838] = 256'h0402030402030304020402040203020303030303030402030303030100080000;
    encBuf[1839] = 256'h010200010002040503050203020302010100020102080a0e0b0c08080008090c;
    encBuf[1840] = 256'h0d0c0d0c0d0c0c0a0c0b0a0c0b0b0b0c0b0c0b0c0b0a0b0a090a0a0a090b0b0c;
    encBuf[1841] = 256'h0c0a0b0a0a0b0b0b0c0a0a0a0908090800090809090809090a0a0c0b0a0c0908;
    encBuf[1842] = 256'h0902070405040304030404030403030203030604030403030403030402030302;
    encBuf[1843] = 256'h03030303020302020000090a0a0c0a090901030101010d0c0d0d0b0b0b0c090a;
    encBuf[1844] = 256'h0a080a0b0b0c0b0b0e0b0c0d0b0c0a0b0b0d0b0c0b0c0a0b0b0a0b0a09090908;
    encBuf[1845] = 256'h0a0b0a0d0c0a0c0c0b0c0b0b0b0b0b0b0a090900020304050204030302030102;
    encBuf[1846] = 256'h0303050403040402040202020100010101020403040401020102060504040302;
    encBuf[1847] = 256'h020201020305030403030302020000080000010000080809090c0c0d0c0c0c0a;
    encBuf[1848] = 256'h0a09080001010203020406040403050304040403030403020303040304020403;
    encBuf[1849] = 256'h03030303020100000008080809080b0d0c0d0b0b0a0a00010002010103050205;
    encBuf[1850] = 256'h030305040304030304030305030403020202020008090b0d0d0c0b0d0b0b0d0b;
    encBuf[1851] = 256'h0b0c0b0c0a0b0b0b0b0c0b0b0b0c0a0b0b0b0a0b0a0909080000000200080008;
    encBuf[1852] = 256'h01020306030200090c0f0b0d0c0b0b0b0a0a09080909090b0b0b0a0901030605;
    encBuf[1853] = 256'h0504040403030404030305030304030303040304020303030304020401020200;
    encBuf[1854] = 256'h010000000008090909090909090a0a090001050201020008000008010908000a;
    encBuf[1855] = 256'h0e0b0f0c0b0e0b0b0d0b0c0c0b0c0b0d0a0c0b0c0c0b0b0c0b0c0b0b0b0c0a0a;
    encBuf[1856] = 256'h0b0a0a0a0a0a090a090a0b0a0a0a090909090908010306030303020008090b0c;
    encBuf[1857] = 256'h0c0b0b0c0a0b0a0a080803060305030305040307030404030303030305030305;
    encBuf[1858] = 256'h030304030303040302030202010100000808090809080909090b0a0a0d0b0e0d;
    encBuf[1859] = 256'h0c0b0c0b0b0b0c0b0b0b0a0b0a0c0b0c0b0a0c0a0c0c0b0b0c0a0b0b0c0c0b0b;
    encBuf[1860] = 256'h0b0b0c0b0c0c0b0c0b0c0c0a0a0a090a090a0a0a080a09090900010304030101;
    encBuf[1861] = 256'h030206040203040103020109090d0a0000040503040404030402020301020208;
    encBuf[1862] = 256'h00000a00010003060203040103030104040204030203030303030000090b0a0a;
    encBuf[1863] = 256'h0d0b0d0a09010404030202010307030505030504040304040203030203030404;
    encBuf[1864] = 256'h0303050203030202020001010101010008090b0b0c0b0b0b0c0b0a0a08010105;
    encBuf[1865] = 256'h0303050402060305030403030303030403020202030202010a0b0f0c0b0d0b0d;
    encBuf[1866] = 256'h0b0d0b0c0b0c0b0b0c0b0c0b0a0b0b0b0c0a0a0b0b0b0b0b0b0c0a0b09090808;
    encBuf[1867] = 256'h000000010302020108090a0b0c0d0d0c0b0c0a0b0c0b0c0b0a0b0a0a0a0a0801;
    encBuf[1868] = 256'h0203050503060404030404030403030403040303040303030403040302040302;
    encBuf[1869] = 256'h03040201020101020101010809080809090a0b0b0b0a0a0d0b0d0a0a0909090a;
    encBuf[1870] = 256'h0c0a0c0a0c0c0b0d0b0c0b0c0b0c0c0a0b0b0b0b0d0b0b0d0b0b0d0b0b0d0a0b;
    encBuf[1871] = 256'h0b0c0a0b0b0c0a0b0a0b0a0a0b0b0a0c0a0a0b0b0d0a0a0a0808080008000203;
    encBuf[1872] = 256'h0404020304040304030203030404030303040305030403020204040304040303;
    encBuf[1873] = 256'h050303040204020303040203010201020101010001000000080808000000080b;
    encBuf[1874] = 256'h0b090b0c0c0f0e0b0d0b0b0c0b0b0b0c0b0b0c0b0c0b0c0a0b0b0b0d0a0b0b0c;
    encBuf[1875] = 256'h0a0b0a0b0c0a0b0b0b0b0c0a0a0a0909090100010208080a0b0d0b0d0c0b0c0b;
    encBuf[1876] = 256'h0a0a0a0008030504040302020108000009080001060504040404030403030402;
    encBuf[1877] = 256'h02030202020101020001020203040306030303030009090a0a0a08010203010c;
    encBuf[1878] = 256'h0f0e0b0c0a090a08090900080305040605040305030402030303030303040304;
    encBuf[1879] = 256'h03050203020202010202020203030502030200080a0d0b0b0c0a090908080a08;
    encBuf[1880] = 256'h000104050406040305030403020203030302030203020301080b0d0d0c0b0c0b;
    encBuf[1881] = 256'h0c0b0c0b0d0b0d0b0b0b0b0c0b0b0c0b0b0c0b0c0a0b0b0a0909090908000000;
    encBuf[1882] = 256'h01000008080000020000090c0c0c0c0c0b0b0b0b0b0c0b0b0c0c0b0c0c0c0a0a;
    encBuf[1883] = 256'h0a09080008020405030603030603040403030403020402030303040304020302;
    encBuf[1884] = 256'h020203020303020202010008090a0a09090a0b0c0d0b0b0c0a0b0c0a0a0a0909;
    encBuf[1885] = 256'h0a09090908090c0b0f0b0a0c0b0a0e0b0c0c0b0c0b0c0b0c0c0a0c0b0c0b0c0b;
    encBuf[1886] = 256'h0c0b0c0b0b0b0b0b0b0c0a090a0a0a0a09090808010001030304030303020304;
    encBuf[1887] = 256'h03040100090b0c0a0a0808010205040404020101000102030203040306040404;
    encBuf[1888] = 256'h040303050303050304030303030303030303030302030200080e0d0c0c0b0b0c;
    encBuf[1889] = 256'h0b0b0c0b0a0c0b0a0c0b0b0b0c0a0a0b0a0d0b0b0c0b0b090a08000801010101;
    encBuf[1890] = 256'h000a0a0d0c0a0b0b0b0e0c0c0c0b0b0c0a0b0b0b0b0b0b0b0b0b0a0b08020101;
    encBuf[1891] = 256'h0302030603040402010303060503040402020301020402040303050303030302;
    encBuf[1892] = 256'h0100090801080100090a00090205010104020505030404020203030402020202;
    encBuf[1893] = 256'h0101010808090b0c0b0c0a0a090a0c0e0b0d0a09010605040404030304030204;
    encBuf[1894] = 256'h0202040304040303030302030102030204030403040102000808090909090a0a;
    encBuf[1895] = 256'h0a0e0b0b0d0a0a0901040405040303040302030204020304020202020000090a;
    encBuf[1896] = 256'h0b0d0c0b0d0b0c0d0b0c0c0b0c0b0b0c0b0c0a0b0a0c0a0b0b0b0b0b0a0a0a0a;
    encBuf[1897] = 256'h0a0a0a0a0909080000020303030200080a0a0b0b0e0b0c0c0b0b0b0c0c0c0c0b;
    encBuf[1898] = 256'h0c0b0b0a09090102040404050305030503030503030502030403030403040303;
    encBuf[1899] = 256'h030403030402030202020201010101010000000800000000080809090b0e0c0c;
    encBuf[1900] = 256'h0c0a0a09090a0b0b0c0b0b0a0c0b0e0c0a0c0b0c0b0b0c0c0b0a0c0c0a0b0c0b;
    encBuf[1901] = 256'h0c0b0b0c0a0b0b0c0b0a0b0a0b0c0c0b0b0b0b0a0b0c0b0b0b0a0b0909090800;
    encBuf[1902] = 256'h0100010000010101030305030404020304040403050303030304030403030403;
    encBuf[1903] = 256'h06040403040304020402030303020302030302020202010202010201080a0b0f;
    encBuf[1904] = 256'h0c0c0b0b0b0c0c0b0b0c0a0b0c0b0b0c0a0b0c0b0d0b0c0b0b0b0c0b0a0b0b0a;
    encBuf[1905] = 256'h0b0a090a0a090c0b0c0c0c0b0b0c0b0d0b0b0c0b0a0b0a090900010100080b0a;
    encBuf[1906] = 256'h0a0a09000a0a090b09000b0e0b0c090103070402040404030602030403040303;
    encBuf[1907] = 256'h0203020204020403030503020202010103030504030203020000090a0b0c0a09;
    encBuf[1908] = 256'h09090a0b0d0d0c0b0b0c0a0a0908090102030604040405040503050303030303;
    encBuf[1909] = 256'h0403030304030403030402030101010101020102020000090b0d0d0c0b0b0a08;
    encBuf[1910] = 256'h0800010008080800040405050304040303040202020203030402020108090b0e;
    encBuf[1911] = 256'h0b0d0b0c0b0c0b0c0b0d0b0c0b0d0a0b0b0c0a0b0a0b0b0b0c0b0a0b0b0b0a0b;
    encBuf[1912] = 256'h09090808000001020302030302030202080c0d0d0c0b0c0c0a0c0a0b0b0c0b0b;
    encBuf[1913] = 256'h0b0c0a0a0b0a0a08010205030604040404030502040203040203040303030403;
    encBuf[1914] = 256'h04020303030303030202010100000809080b0a0c0b0b0c0a0b0a0b0a0b0a0a0a;
    encBuf[1915] = 256'h0b0b0a09010404050302040102020808090d0b0c0d0c0c0c0c0b0d0b0c0c0b0c;
    encBuf[1916] = 256'h0b0c0b0c0c0b0b0b0b0c0b0b0c0a0a0b0a0a0a0a090908080001010202040304;
    encBuf[1917] = 256'h040303030304030303030100090a0a0b0c0c0c0b0c0c0a0b0c0c0b0b0a0a0801;
    encBuf[1918] = 256'h0205040503040402040203030404030403030304030303040302030301010008;
    encBuf[1919] = 256'h0b0c0c0c0b0c0b0b0b0c0a0b0b0b0c0c0b0b0c0a0b0b0a0b0b0b0b0b0a0a0802;
    encBuf[1920] = 256'h03050403020201000809090a0b0c090c0c0c0d0c0b0c0b0c0a0b0b0c0b0a0c0b;
    encBuf[1921] = 256'h0a0c0a0b0a0a0a0a0a0809080001020603040503030502030203030304030403;
    encBuf[1922] = 256'h0302010000080000080000090002000305030505030404020304020101000008;
    encBuf[1923] = 256'h0908000802000002080902020706040304030306030405040403050304030402;
    encBuf[1924] = 256'h02030303040303040402020302010101010101020301020108080c0d0b0b0b0a;
    encBuf[1925] = 256'h090a09090a09090902050506040403040303030304030304020202020201090a;
    encBuf[1926] = 256'h0b0f0b0d0c0b0c0c0b0b0d0b0b0d0b0b0b0c0b0b0c0a0b0b0b0c0b0a0b0b0a0a;
    encBuf[1927] = 256'h0a090808000800000808000001020203020201080a0d0c0c0c0a0b0c0b0c0b0c;
    encBuf[1928] = 256'h0b0b0b0a0a080203050604030603040305030305030304030304030402030402;
    encBuf[1929] = 256'h03030403030304020203010101010100000800090909090a0a0b0b0b0c0a0a0b;
    encBuf[1930] = 256'h0c0b0e0b0c0c0c0a0b0a0a0a0a0a0a0c0a0b0c0b0d0b0b0c0b0c0c0c0b0d0b0c;
    encBuf[1931] = 256'h0c0b0b0c0b0c0b0b0b0d0b0b0b0b0c0b0a0b0b0b0b0c0a0b0b0a0a0909000001;
    encBuf[1932] = 256'h000008090a090a00010404050304030204020304040304030302020201020104;
    encBuf[1933] = 256'h0404040403040303040303040303050304030303030304020302030302020301;
    encBuf[1934] = 256'h00090c0c0c0d0b0b0b0d0a0b0a0b0d0b0b0c0c0a0b0b0a0b0b0c0b0c0b0b0b0b;
    encBuf[1935] = 256'h0b0a090808010808080b0d0b0c0c090a0b0b0c0c0b0e0b0b0c0b0b0c0b0a0b0c;
    encBuf[1936] = 256'h0a0c0a0a0b0b0a0a09000002040202030808000a090202070603040403030401;
    encBuf[1937] = 256'h02030104030306030304030202030305030304030203010008090b0a0a0a0000;
    encBuf[1938] = 256'h0800090c0a0c0b08080307070404030304030306030405030403040303030402;
    encBuf[1939] = 256'h030304030304030203010201000001000201000100090a0a0e0a090b08080908;
    encBuf[1940] = 256'h080c090a0b090103070705040203030203020302040302030200090b0e0b0e0b;
    encBuf[1941] = 256'h0b0d0b0b0d0b0c0c0c0a0c0b0b0c0b0b0b0b0b0c0b0b0c0a0a0b0a0a0a0a0909;
    encBuf[1942] = 256'h090908000001010202020202020101080009090909090a090b0b0b0f0d0c0c0c;
    encBuf[1943] = 256'h0a0b0a0808020505040404040404030403040304020304020402030304030304;
    encBuf[1944] = 256'h020402020302030202010202010100000009090b0c0b0d0b0c0c0b0b0b0c0a0b;
    encBuf[1945] = 256'h0a0b0c0b0b0c0b0a0b0a0a0b0c0a0c0c0a0b0b0c0b0b0c0d0b0b0d0c0b0b0c0c;
    encBuf[1946] = 256'h0b0b0c0c0a0b0c0b0b0c0a0b0b0b0b0b0c0c0a0b0a0b0a0a0a09080800000000;
    encBuf[1947] = 256'h0808000800030306050204030303050203040304030302020101020102030103;
    encBuf[1948] = 256'h0303060403050303050304020402020303030403040502040303020302020101;
    encBuf[1949] = 256'h01000000000b0c0c0d0c0a0b0c0b0c0c0b0b0d0b0b0b0b0b0a0a0a0b0a0c0a0a;
    encBuf[1950] = 256'h0b0a080801020303050202030100010a0a000a0a0b0f0f0c0b0c0b0c0b0b0c0a;
    encBuf[1951] = 256'h0a0b0a0b0c0c0a0b0c0a0b0a090a090000020402040402030503040503050203;
    encBuf[1952] = 256'h0203030304040304030302010108090a0a0a09090b0a0c0d0b0d0c0a0b090900;
    encBuf[1953] = 256'h0205040403030404040306030404030304020303040204020303040202010101;
    encBuf[1954] = 256'h00000800080008080a0c0b0c0d0a0a0a09080001010002010104040405040304;
    encBuf[1955] = 256'h040203020203020203040204010108090b0d0c0c0b0c0b0b0d0c0b0c0c0b0b0c;
    encBuf[1956] = 256'h0b0b0c0a0b0b0c0a0b0b0b0a0b0a0b0a0a090908080100010102020302030302;
    encBuf[1957] = 256'h030301090c0f0c0b0d0b0c0c0b0b0b0b0b0c0b0b0c0a0a080801040404040303;
    encBuf[1958] = 256'h0503050305030403040303030403020403030303040302030202010201010101;
    encBuf[1959] = 256'h02010201010808090c0b0c0c0a0b0c0b0b0d0a0a0b0a0b0b090a0a090a0a0808;
    encBuf[1960] = 256'h0002080a0c0f0c0a0c0a0a0c0c0b0f0c0b0c0b0c0b0b0b0d0b0c0c0b0b0c0b0b;
    encBuf[1961] = 256'h0c0a0b0b0a0b0c0a0a0a0a090908000102030203030304030503040403030302;
    encBuf[1962] = 256'h010100080808090809090a0b0d0c0c0b09080003040202010800000004040306;
    encBuf[1963] = 256'h040204030403040203030304030404030402030102020001010008080c0d0c0d;
    encBuf[1964] = 256'h0c0c0b0b0c0c0b0b0b0b0b0b0b0a0b0c0b0b0b0b0a0a00080103010103020407;
    encBuf[1965] = 256'h0404040304020100000909090b0a0c0c0b0c0c0b0b0b0c0a0c0b0a0b0b090a0a;
    encBuf[1966] = 256'h0009010202040503030502020201020403040502030401020201020302020209;
    encBuf[1967] = 256'h0a0c0d0b0a0901040203010c0d0e0c0b0a090800010100010203050704050403;
    encBuf[1968] = 256'h050303030402030203040305030304020301020201010101010101080a0c0c0b;
    encBuf[1969] = 256'h0b09090800010800090c0a090a02070405030403030203030404030403030302;
    encBuf[1970] = 256'h0009090d0b0d0b0b0c0b0b0d0b0d0b0c0b0c0b0b0b0b0c0b0c0b0c0b0c0a0a0a;
    encBuf[1971] = 256'h090a09090a090a0a0909000001010201000001010202020301090b0f0e0c0b0d;
    encBuf[1972] = 256'h0b0b0b0b0c0b0c0b0a0b0b090a08010306040404030403050304040304030304;
    encBuf[1973] = 256'h030204030304020303020101000000080809090a0c0b0c0b0c0a0b0a0a0a0a0a;
    encBuf[1974] = 256'h0a0a0b0b0909010001040405040404030203020201000a0b0c0d0b0c0b0d0a0b;
    encBuf[1975] = 256'h0c0a0c0c0b0d0c0a0b0b0b0b0c0b0c0b0c0b0a0b0a0909090909090808000103;
    encBuf[1976] = 256'h050403030402020202020303030402030200090b0e0d0b0d0b0b0c0a0b0b0b0a;
    encBuf[1977] = 256'h0b0b0a0a08010203050204040405040304030304030303030304040203030101;
    encBuf[1978] = 256'h080b0c0c0c0b0c0a0b0b0b0c0b0c0b0a0a0a0909080909090809080809000204;
    encBuf[1979] = 256'h07030503030303040303040302020000090b0c0b0c0b090b0b0b0d0c0c0c0c0a;
    encBuf[1980] = 256'h0b0c0b0c0c0b0b0c0a0a09080101020008090a0a000205070304030303020201;
    encBuf[1981] = 256'h0403040403020300080a0e0b0d0b0c0a0a090a0b0c0b0d0b0c0a0a0909080008;
    encBuf[1982] = 256'h0808090001040604050305020402030304030403040302030303030403030402;
    encBuf[1983] = 256'h0303030202010101010001010008090a090b0802040703040304030304030504;
    encBuf[1984] = 256'h040403040303020302020303030403020208090b0c0d0a0c0b0b0d0c0b0e0b0c;
    encBuf[1985] = 256'h0b0c0b0b0c0a0b0b0a0b0c0a0b0b0b0b0a090a0a090b0a0b0c0a0b0a0a090809;
    encBuf[1986] = 256'h090b0e0b0d0b0c0b0c0a0b0a0b0c0c0c0b0b0b0b0a0a0a090808000801010307;
    encBuf[1987] = 256'h0503040203040304040304040304030402030303040402030303030303040302;
    encBuf[1988] = 256'h04020302030302020100000808000008090a0f0c0c0c0b0a0909080808000909;
    encBuf[1989] = 256'h0a0b0d0a090a000801030302040008010909090f0f0c0c0c0b0c0b0b0c0b0b0c;
    encBuf[1990] = 256'h0b0a0b0b0b0b0c0a0b0c0a0c0b0a0c0b0b0a0909000001020202030302010200;
    encBuf[1991] = 256'h090a0d0d0c0b0c0b0a09090908000a0b0e0d0c0b0b0a0a0b0b0a0d0a09090800;
    encBuf[1992] = 256'h0808010001040000010909000a09090e0d0b0e0b0b0c0a090908080b0c0c0d0b;
    encBuf[1993] = 256'h0b0d0a0b0d0b0a0b0b090a090808080001020503050502020402030404040303;
    encBuf[1994] = 256'h020301010202010300090b0f0c0c0c0b0c0b0b0a0b0909090801000102010103;
    encBuf[1995] = 256'h00030403040403040303040403050402030202010201010108090a0f0c0a0c0b;
    encBuf[1996] = 256'h0a0b0a080a0a0a0e0b0d0b0d0b0b0c0a0b090908000002040405040304030304;
    encBuf[1997] = 256'h0403040403030503030404030303040303020402020302020202010100000808;
    encBuf[1998] = 256'h0800090000080001090003010605040504040403030403020304020403030303;
    encBuf[1999] = 256'h0101080a0b0c0c0b0c0c0b0b0d0c0b0c0b0d0a0b0b0a0b0c0b0a0c0b0b0d0a0b;
    encBuf[2000] = 256'h0a0b0a0a0a090a0a0909090808080009080a0b0d0c0c0c0b0c0a0a0a0a0a0c0c;
    encBuf[2001] = 256'h0b0d0b0b0c0b0b0c0b0c0a0b0a0a090908010103040405040305020303030403;
    encBuf[2002] = 256'h040203040304030404020303030202010101000102010000090b0c0b0b0a0901;
    encBuf[2003] = 256'h02040303020000090b0c0c0c0c0b0b0c0b0c0c0c0a0a080002040201080a0e0c;
    encBuf[2004] = 256'h0c0b0c0a0909080000010100000808080001000a0d0f0d0c0c0c0b0a0b0a0908;
    encBuf[2005] = 256'h080000010108090b0d0c0b0c0b0a090900000000000001030504040302010100;
    encBuf[2006] = 256'h080a0c0d0b0b0b0b0900020404040108090a0b090909080b0a00080306020307;
    encBuf[2007] = 256'h030504030402010100090a0b0e0b0c0b0b0b0b0a0a0a08010105040402030100;
    encBuf[2008] = 256'h090c0c0c0b0c090a0900000000090909090106030503020000090b0b0e0a0900;
    encBuf[2009] = 256'h020604040403020208090b0c0d0a0c0a0a0a0a0a0a0909080802010304020203;
    encBuf[2010] = 256'h080a090e0b090b090800020604030501010009000101030301090c0f0b0d0b0c;
    encBuf[2011] = 256'h0b0b0a0b0a0a0800010303040304060404050305030403040304030303040303;
    encBuf[2012] = 256'h0304030303030303030302040302030402020201010009090a0b080808020401;
    encBuf[2013] = 256'h040403060403050403030402020201020404040304030202010009090c0d0b0c;
    encBuf[2014] = 256'h0c0a0c0c0b0b0c0b0c0b0b0a0c090b0a0b0b0d0b0c0b0a0b0a0a0a0a09090a0a;
    encBuf[2015] = 256'h090a08000001010001090a0b0f0b0b0b0a090808090d0d0c0d0c0b0b0c0b0b0b;
    encBuf[2016] = 256'h0a09080800000001030505040403030503040303040303040203030403030304;
    encBuf[2017] = 256'h0303030203020100000a0b0d0c0b0b0b0b0b0c0b0a0b0c0b0d0c0a0a09080100;
    encBuf[2018] = 256'h080a0b0d0b0b0a080204060504030403020200000809090a0a0909090a09090a;
    encBuf[2019] = 256'h090a0b0c0e0d0d0b0d0b0c0b0b0c0a0a0b090a0a090a09080101030303020202;
    encBuf[2020] = 256'h05040404020202010100080a0a0b0b0a0909080d0e0d0d0d0b0c0b0b090a0808;
    encBuf[2021] = 256'h090a0b0b0b0b0a09080900010002080b0d0e0b09080104040403000000090900;
    encBuf[2022] = 256'h0002010809080d0b0d0d0a090a08000809080b0c0c0e0c0a0b09000001020202;
    encBuf[2023] = 256'h0504040502030402030303030303040304040403030303020100090a0e0c0c0c;
    encBuf[2024] = 256'h0b0c0c0a0b0a0b0a0a0900080102000100080808090803060505030503020303;
    encBuf[2025] = 256'h0101000809080809090b0d0c0b0c0b0b0d0b0b0a0a0900010304030403040304;
    encBuf[2026] = 256'h0403040305040404040302040202020202040203040304030303040202010008;
    encBuf[2027] = 256'h0000010202030302020402030200080909020504050304030402030303040304;
    encBuf[2028] = 256'h040303050303030402020008090b0e0c0b0d0b0c0b0c0b0c0c0b0b0b0c0b0b0b;
    encBuf[2029] = 256'h0b0a0c0a0a0a0a0a0b0b0b0d0a0a0a09090b0b0b0c0a0a0b0a0a0b0d0b0d0b0b;
    encBuf[2030] = 256'h0c0b0a0b0a0b0b0b0b0c0b0b0c0d0b0c0a090102040302020101020202020306;
    encBuf[2031] = 256'h0406030502020201010103050404040304020101000808080808010002020302;
    encBuf[2032] = 256'h02010008090a0d0d0b0a0c090a09080001030503040202010000020407040503;
    encBuf[2033] = 256'h02020108090a0c0a0c0b0c0b0b0a090908090a0b0d0b0b0b0c0b0b0a0a0a0001;
    encBuf[2034] = 256'h030404030302020101020306030201090e0c0d0c0c0b0d0a0b0909080001080a;
    encBuf[2035] = 256'h0b0e0b0b0c0b0c0b0c0b0a0a08000801000008090b0c0d0b0b0b0b0909000103;
    encBuf[2036] = 256'h0304080c0d0d0b09090002010202000800090801010406020203090a0d0d0c0a;
    encBuf[2037] = 256'h0b0a0002060404040202020008090a0a09010306050305040303020100000908;
    encBuf[2038] = 256'h090a0a0a0a08000205030302010a0d0c0d0a0900020403040303040201080a0b;
    encBuf[2039] = 256'h0900040704020301080a0c0b0b0a08010203020100080000090b0f0d0c0a0900;
    encBuf[2040] = 256'h01020403030202020008080a0c0c0b0a02060704040302030101000000000103;
    encBuf[2041] = 256'h0306040403050303040202020201030203040203020100000900020306030202;
    encBuf[2042] = 256'h02020203030504040405030503030402000008090a0a0a08080003030203010a;
    encBuf[2043] = 256'h0d0d0d0a0c0a0a0b0a0a0b0d0b0d0c0a0b0b0a09090008090a0c0f0b0e0b0b0b;
    encBuf[2044] = 256'h0b0a0a09000000010109090b0f0b0d0b0b0c0a090a08080008000009080a0b09;
    encBuf[2045] = 256'h0a0909090a0a0b0e0b0e0c0b0b0b0a0800030405030402030202020304030403;
    encBuf[2046] = 256'h03040102000102020404040203030200090e0e0c0b0c0b0a0b0a0a0901020504;
    encBuf[2047] = 256'h040304030301000a0d0c0c0b0b0a0b090800000102020103020201000a0c0d0d;
    encBuf[2048] = 256'h0b0c0c0b0a0908010305040302020109090d0b0d0b0d0a0c0a090a0808080101;
    encBuf[2049] = 256'h000101080a0c0f0c0b0b0c0b0b0b0a0b0a0a090a09090001010201090a0c0d0c;
    encBuf[2050] = 256'h0b0b0a09010406020303010201020306020403030303000a0b0d0b0908020403;
    encBuf[2051] = 256'h03030102040205030303010a0b0d0b0a01050705040404020302020101000001;
    encBuf[2052] = 256'h0101030303030102010306050305020202000009090908000002010101020204;
    encBuf[2053] = 256'h0404030403020100090a0a0a09000102040504030100090b0a08030704030201;
    encBuf[2054] = 256'h090c0e0c0c0b0a090a090a0c0a0b090800010102030604040402020201010009;
    encBuf[2055] = 256'h0a090802070404040203040102010008080b0909080104030603020201000100;
    encBuf[2056] = 256'h0001030104030306040203030100080801050405040303040203030203030103;
    encBuf[2057] = 256'h0403060303040301030101000109000801040402040208090d0e0b0c0b090a08;
    encBuf[2058] = 256'h000808000908000a0f0d0d0d0a0c0a0a0a09090908000808090a0b0c0d0c0c0b;
    encBuf[2059] = 256'h0b0b0a090908090a0b0d0b0b0b09090001080a0b0f0b0c0c0c0a0b0a09000103;
    encBuf[2060] = 256'h040302000a0e0d0c0b0a0a090909090909090908000000010001080008090909;
    encBuf[2061] = 256'h0e0d0b0b0a010306030202020100000a0b080901050303030000080f0b0b0e09;
    encBuf[2062] = 256'h0909000202040301090d0f0c0a0a080202040303030402050403030302000a0d;
    encBuf[2063] = 256'h0d0a0b09080203040301010a0d0d0c0c0a0a090001010200090b0f0b0c0a0a08;
    encBuf[2064] = 256'h0001030302010008000003040302040103050303040202030008080d0c0c0d0b;
    encBuf[2065] = 256'h0a0a09080102030200080c0d0b0e0a0909010203050303020200010102040503;
    encBuf[2066] = 256'h0303020304030604040304020302010101010202010202020203020304050404;
    encBuf[2067] = 256'h030403020100080800000404040403020208000002050505040302020109090a;
    encBuf[2068] = 256'h0b080204050304020008090b0d0b0d0b0b0a0908080100000008080000000101;
    encBuf[2069] = 256'h0109080909020606050303030301030101090c0f0b0d0b0a0a0a000203070302;
    encBuf[2070] = 256'h03020000090b0a0a0b0801000202010504040604020403020301000008090001;
    encBuf[2071] = 256'h0206040404040303030201010808090908010205030305030204020101090b0d;
    encBuf[2072] = 256'h0c0c0a0a0a09090908080802020304010800090a08090b0a0f0f0b0d0c0a0c0a;
    encBuf[2073] = 256'h0a0a0b0c0b0c0b0c0b0a0b0b0b0c0b0a0b0b09090800080b0d0e0c0b0c0b0b0a;
    encBuf[2074] = 256'h0a09080809090c0c0d0c0c0c0b0a0b0b0908080101020102030100080c0d0c0c;
    encBuf[2075] = 256'h0c0a0a09080000020100080b0e0b0d0b0b0a09000103040403030200080a0c09;
    encBuf[2076] = 256'h0900040405040203010000080808000800000101040304030100080a0a090902;
    encBuf[2077] = 256'h07060404030403010100080a0b0d09090802040303040202020808090b0a0909;
    encBuf[2078] = 256'h0003050505040304020100090c0d0c0c0a0a0a090800000000080008080a0a0d;
    encBuf[2079] = 256'h0c0c0a0b090001040403040203010108000808080102020402030300000b0f0c;
    encBuf[2080] = 256'h0c0b0b0c0b0c0b0c0a0900010402030100080800020704050303020101020204;
    encBuf[2081] = 256'h0303030303030603040402010000090a0a0a0800030605040304030101080a0d;
    encBuf[2082] = 256'h0c0b0a0800030305020302010101000800080002040504040304030402020302;
    encBuf[2083] = 256'h020304020100090a0b0c0a090a090801020401090c0f0c0a0a08000104040403;
    encBuf[2084] = 256'h0303020302020201080a0b080407060403040202010108090b0b0c0b0a0a0000;
    encBuf[2085] = 256'h040403040101080a0b0c0c0b0b090803060404030101090c0b0b0a0003060403;
    encBuf[2086] = 256'h03020000090a0b09000207030404020201080a0c0c0b0c0a0a0a0a0a0a0a0a0a;
    encBuf[2087] = 256'h0c0b0c0b0d0a0b0b0b0d0b0b0b0c0a09080203040401000a0d0e0b0d0b0a0a09;
    encBuf[2088] = 256'h0800000108080b0e0c0c0b0b0c0a0a09080801010101000a0c0e0b0d0a0a0909;
    encBuf[2089] = 256'h000801000808090b0b0c0c0a0a09000204030602020200080a0c0c0a0b0a0908;
    encBuf[2090] = 256'h0002020202090a0b0f0a09000205040403020302020203020403040504020303;
    encBuf[2091] = 256'h0201020103050404030303020102010205030403030302020001000a0b0c0c0a;
    encBuf[2092] = 256'h0002050502030208080b0c0c0b0b0b0a0b080207060403040201000809090909;
    encBuf[2093] = 256'h0a0a0a0b090a010304040200090b0f0c0b0c0a0908010000000808090a0b0c0a;
    encBuf[2094] = 256'h0a0000020202010102040504040504030503030203010108080808000100080a;
    encBuf[2095] = 256'h0c0d0c0c0b090902040504020302000008090901030705040403030201010101;
    encBuf[2096] = 256'h01020403020208090b0b0a0204050301090c0e0d0b0b0a090001020202020108;
    encBuf[2097] = 256'h0a0d0d0b0b0a08010204030303030000090900010405030403030202080c0e0b;
    encBuf[2098] = 256'h0d090908090a0d0c0c0c0b0b09080002030300080b0d0b0b0804060404030301;
    encBuf[2099] = 256'h00080a090b080801050304030202000809090b0b0b0b0b090a0c0c0d0d0b0b0a;
    encBuf[2100] = 256'h080305050402020109090b0b0800040505030403020100080809000205040404;
    encBuf[2101] = 256'h02020108090b0d0b0b0a0a09090000010201080b0f0f0b0d0a09090801020302;
    encBuf[2102] = 256'h0201080a0c0b0c0b0a0909000002040203040100080b0e0c0c0b0d0b0b0b0c0b;
    encBuf[2103] = 256'h0b0c0b0b0c0b0b0b0b0908000000090b0e0b0d0a0a0808010000080a0c0b0c0a;
    encBuf[2104] = 256'h09080203050302090c0d0d0b0c0a0900010304030201080c0c0d0b0c0a0a0800;
    encBuf[2105] = 256'h010203030302010200000008000102050503040202010100010302030300090b;
    encBuf[2106] = 256'h0f0d0a0a08000001000809090c0d0b0d0b0a0901040304030100090b0c0b0a08;
    encBuf[2107] = 256'h01020304080a0b0e0a0103070404020200090a0d0c0a0a080203060403030301;
    encBuf[2108] = 256'h00090b0c0a0a000403060304020302010108090a0b0b0a0b0a0b0b0a00010604;
    encBuf[2109] = 256'h0404040304030202010102030405050306030403020301000909090a09090800;
    encBuf[2110] = 256'h0102040303020100090a0a0000090c0f0d0b0b09010605040403030201010008;
    encBuf[2111] = 256'h090800080008000002050504040203020101000809090b0b0b0c0a090a000101;
    encBuf[2112] = 256'h01090c0b0c0901020302000a08090107030605040305030201080b0c0d0c0a0b;
    encBuf[2113] = 256'h0908000100090c0b0e0b0a0b0a0b0b0d0b0c0b0b0c0a0a0b0a0a0a0800010204;
    encBuf[2114] = 256'h03040302020200000102030604030302010a0d0f0b0d0b0b0c09090908080008;
    encBuf[2115] = 256'h00010001090a0a0b080307060304020202010101010302030202010202040405;
    encBuf[2116] = 256'h030302000808090001000303040504040305030403020100090b0c0d0a0b0b08;
    encBuf[2117] = 256'h010405040303030000090a0b0a0909090a0a0a08020503020b0f0f0e0b0c0a0b;
    encBuf[2118] = 256'h0b0b0b0b0b0a0a0908000808080b0b0e0c0c0b0c0a0a09000205040402020100;
    encBuf[2119] = 256'h090b0d0c0d0b0a0b09090000010008090c0c0b0b0a0900010202040403040402;
    encBuf[2120] = 256'h020201080a0b0a080103060201090b0d0b0b080106050403020100090b0a0b09;
    encBuf[2121] = 256'h0002040505030303010101010403050303020100090c0d0b0b0a080203050403;
    encBuf[2122] = 256'h0202080b0c0d0b0b0909000203040301090c0d0d0b0b0c0a0908000102020201;
    encBuf[2123] = 256'h0001090a0c0d0a09010407030304010100090a0a0a0908000108080a08080104;
    encBuf[2124] = 256'h020100080c0d0d0c0c0b0b0a0001050404040202020008090a0900000302010b;
    encBuf[2125] = 256'h0f0c0c0b0b0a08090808080a0c0d0c0b0a0a0103060403030101090909080205;
    encBuf[2126] = 256'h040302020008090a0a0a0b0b0b080307060303020108090b0b0c090801050405;
    encBuf[2127] = 256'h020100090c0b0b0a0801030302080b0f0c0a0a0901020201080c0c0c09010405;
    encBuf[2128] = 256'h04030201080a0d0c0b0b0a0a0800020202030100090b0d0c0b09010406040202;
    encBuf[2129] = 256'h00080a0a090a00010305030201090c0c0c0a090800020100000c0c0c0a080104;
    encBuf[2130] = 256'h0404020000090900030606040304030203020202020303010201000404040403;
    encBuf[2131] = 256'h0203020008080908080103030202080d0c0c0b09080102020001080001020407;
    encBuf[2132] = 256'h050403040201080a0a0a0c0b0e0c0b0d0b0a0a0900080009090c0d0c0c0b0b0b;
    encBuf[2133] = 256'h0c0a0b0b0a0a09000203040201090b0d0d0b0a090002040403020108090b0c0b;
    encBuf[2134] = 256'h0b0b0c0c0c0b0c0c0a0a0a0a0a0a0b0c0b0b0a0902030502010a0d0d0b090801;
    encBuf[2135] = 256'h0305040302030201010203050304020000090000030404040404030402020109;
    encBuf[2136] = 256'h0a0c0c0c0b0b0b0002060404020100080a0b0a09010206030402010108080808;
    encBuf[2137] = 256'h08000800000008090a0a0c0d0c0c0c0b0a0a080103050304020008090c0a0a00;
    encBuf[2138] = 256'h030503030201090a0a0b080008090d0f0d0b0a090103050301080b0f0b0c0b0a;
    encBuf[2139] = 256'h0908020306030201090b0c0b0b0908000303050302080d0e0c0c0a0800020305;
    encBuf[2140] = 256'h0201080a0d0c0b0b080204050303020809090b0a09090808090a0b0c0a080406;
    encBuf[2141] = 256'h04040200090c0d0b0b0900010404030200090b0c0c0a0a08010203040201080b;
    encBuf[2142] = 256'h0d0d0b0c0a09080002020303030108090c0b0a0803050503020008090a090001;
    encBuf[2143] = 256'h0103020200090d0e0d0b0b090002040305020303020108090a09000203040404;
    encBuf[2144] = 256'h0405030401080b0e0c0b0a090801020504030401080b0d0b0c0a080103070403;
    encBuf[2145] = 256'h020200090c0c0b0a0901020503040108090c0c0b0a08010305020300000a0a0c;
    encBuf[2146] = 256'h0a0a0800030403030008090b0b0b0a0a0b0a080205040302080d0d0d0b0b0908;
    encBuf[2147] = 256'h010304030208080b09080103000a0f0f0a0a08010306030301000b0e0c0c0a09;
    encBuf[2148] = 256'h00020305030100090b0b0c0908020305030201090a0c0b0a0900000203030303;
    encBuf[2149] = 256'h01000b0e0c0b0c090901030703040301080b0d0b0a0802050404030200080a0b;
    encBuf[2150] = 256'h0d0b0908020504020200090b0c0a0a09090800000202050404030200090c0e0b;
    encBuf[2151] = 256'h0c090801030403020108090b0e0b0c0a0900020304030200090b0c0c0b0b0802;
    encBuf[2152] = 256'h0404040201080a0c0b0b0b090102050303080b0f0b0b08000305020200090b0b;
    encBuf[2153] = 256'h0c0a09020505030301090a0b0b0901030300090d0d0b0c0a0908020405030302;
    encBuf[2154] = 256'h080b0f0c0b0b0900040404030200090a0c0b0a0900020504030200090c0d0b0a;
    encBuf[2155] = 256'h080104040302010a0c0c0b0a000205040301000a0b0d0a0a0801020303030208;
    encBuf[2156] = 256'h0a0c0c0b0b09090101030302010103040303080d0d0c0b090901010102030303;
    encBuf[2157] = 256'h03090d0d0c0b0908000000000204060303080a0e0b0b0a000001020303050302;
    encBuf[2158] = 256'h0201080a0c0e0b0c0a0800030303010101010201090a0c0a0001090f0f0d0a0a;
    encBuf[2159] = 256'h08010204030306030400090c0e0b0a09010303030402020200090d0c0b0a0800;
    encBuf[2160] = 256'h020202020008090c0c0c0b09010405030201090b0d0b0a0a0800020303020809;
    encBuf[2161] = 256'h0b0b0a080307040303080b0f0d0a09000205030202000009090a0b0c0a080205;
    encBuf[2162] = 256'h0303080b0e0a09000204030201020201090d0e0c0b08020604040200080b0b0d;
    encBuf[2163] = 256'h090908010202020202080a0d0d0b0a09000103030108090b0c0b0b0b0a000405;
    encBuf[2164] = 256'h040201080a0a0a08080908080105040202080900020603010b0f0c0a09000203;
    encBuf[2165] = 256'h0200080808010202030202000a0e0e0c0b0a0a0801040604040201090d0c0b08;
    encBuf[2166] = 256'h01040302080a0c0a0900080809000207040301080b0d0b0b0a08010305040301;
    encBuf[2167] = 256'h080b0d0b09000205020201080b0b0d0a0a010306030301080a0b0a0801020201;
    encBuf[2168] = 256'h08090b0a0a0908010102010b0f0f0c0b0a000204040300090d0c0c0a00020504;
    encBuf[2169] = 256'h0302000b0d0b0a0902030501000a0b0b0b0a090a08010407040202090b0d0b09;
    encBuf[2170] = 256'h0002030302010009080900000202010a0f0c0c0a09080000090a0b0a08030705;
    encBuf[2171] = 256'h040201000a0c0b0c09080202030402010100080a0d0c0c0b0b0a000206040402;
    encBuf[2172] = 256'h0108090a0c0b0b0a0901040603030200080a0b0b0c0b0b08010202080b0b0805;
    encBuf[2173] = 256'h070402000a0d0c0a090001030402030100090c0c0a0a0a080000000203050200;
    encBuf[2174] = 256'h0a0d0c0a0a0900020304020108090a0104060401080a0d0b0a08010305030301;
    encBuf[2175] = 256'h000a0c0b0a08000201000a0b0e0b0c0a0a010407030301080a0b090800080c0c;
    encBuf[2176] = 256'h0c0801040402010008010001090b0e0c0a0a080103050503040108090c0b0b0a;
    encBuf[2177] = 256'h0901030703030201090a0c0a0808000108090908020404030200080801020303;
    encBuf[2178] = 256'h080d0f0d0a09000306040301000a0c0c0a0a0908010100000800010203010a0d;
    encBuf[2179] = 256'h0d0a0901010100080105060402080a0e0b0909010201020103040402080c0d0c;
    encBuf[2180] = 256'h0b0a08000202030303020200080c0c0d0c0a080104050301090b0d0b0a080204;
    encBuf[2181] = 256'h05020200090c0b0c0a080000000100020405030201090c0c0c0b090002030403;
    encBuf[2182] = 256'h0101090b0c0b0c090802030302000a0b0803070601000b0e0b0a080203040203;
    encBuf[2183] = 256'h020303000b0f0f0b0a0901020304020200090a0c0c0a09010204020201080a0a;
    encBuf[2184] = 256'h0b0b0b000306040201080a0a0a0a0a0c0a0901050402000a0b0b080306020009;
    encBuf[2185] = 256'h0b0b0a000203040401010b0e0d0b0c0900030504020200090d0c0b0a0a000204;
    encBuf[2186] = 256'h04030301080b0c0c0a090800020100000800010101000b0c0c09010404040100;
    encBuf[2187] = 256'h090b0a090a080a09090307040402080a0c0c0b0801040402010a0d0b0c090001;
    encBuf[2188] = 256'h0203030301080d0b0b01040602000a0d0c09080202010009090801020202000a;
    encBuf[2189] = 256'h0c0c0a0903060401090e0c0a09020403030109090a090900000002010a0f0e0b;
    encBuf[2190] = 256'h0a010406030301000a0b0e0b0c09080104040202080a0b0c0a08000304020109;
    encBuf[2191] = 256'h0b0d0a0001030101090a0900000809080105060302090c0e0b0a000103030300;
    encBuf[2192] = 256'h0a0c0b09000102000a0a090003010a0d0c08040603010a0c0d0a090002020202;
    encBuf[2193] = 256'h01090d0c0c0900020303000a0c0b09010305030303090c0f0c0b090002030302;
    encBuf[2194] = 256'h02030403090d0f0b0b080304040300000a0909080809080a0a0b0a0803070403;
    encBuf[2195] = 256'h020000000808090d0d0b0b0a00010203030305030200080b0c09010405030108;
    encBuf[2196] = 256'h0c0e0b0b0801030302090d0d0a08030704020200090a0b0c0a0a090002050302;
    encBuf[2197] = 256'h00090b0a01040502000a0c0d0a0a0808020306040202080a0d0b090801010109;
    encBuf[2198] = 256'h0a0a000405040208090c0b0b0900000101000102050303000a0e0c0b0b000104;
    encBuf[2199] = 256'h0304020101090c0b0b0a01050301080c0b0a0001020009090107060202080909;
    encBuf[2200] = 256'h000202000b0f0c0b08000304020101000808080909080008090d0c0a00040603;
    encBuf[2201] = 256'h030200080a0b0e0b0c0a010406020208090c0a0a08020203030000090a0a0801;
    encBuf[2202] = 256'h00080b0c0c0a0802050403040202000a0d0d0a090104040201080b0c0a090103;
    encBuf[2203] = 256'h040208090b0a0a08010306040404030200080a0c0e0c0d0a0b08020603030200;
    encBuf[2204] = 256'h090a08000001090b0c0a08020301090d0c0a000405030201080908080000090b;
    encBuf[2205] = 256'h0d0b09020302000c0d0c080205050302080a0c0b0b0908010202030100080800;
    encBuf[2206] = 256'h02040401080c0c0a000303080f0e0c09010405040100090a0c0a0a0800000000;
    encBuf[2207] = 256'h000000020203010101000001080a0f0d0b0b0b000205040300090d0c0b080205;
    encBuf[2208] = 256'h040200090b0a0a09080a0a0b0803060302090c0c0900030402080a0c0c0b0b08;
    encBuf[2209] = 256'h0105050301000b0c0a09000200080a0b0b0901020204040302080d0c0c090001;
    encBuf[2210] = 256'h01080a0d0a080306040201080b0c0c0a0a01020402010b0d0b09010603030109;
    encBuf[2211] = 256'h0c0b0b0a0800000000010202030403010a0f0c0b0b08020303010a0e0b0a0001;
    encBuf[2212] = 256'h0403030201010108090c0c0b0a0a0a0b0c0a0804060401080b0f0c0a09080103;
    encBuf[2213] = 256'h050302000a0c0c0a0901030401080a0d0a0a000204030301080d0c0b0a090102;
    encBuf[2214] = 256'h0201090b0b0803060401080b0d0b0c090801030505030201080c0d0b0b0a0002;
    encBuf[2215] = 256'h020301010009080b0b0c090104050302000a0c0d0a0a080205040301080c0d0b;
    encBuf[2216] = 256'h0b0a00010202030304030400090b0f0b0b0a0a00010405030200080a0a080103;
    encBuf[2217] = 256'h0401090e0c0c0b09000204040201090b0b0b0902030302010801020306030201;
    encBuf[2218] = 256'h080a0e0d0c0a0a080203050302010200090c0d0c0b08010404030200090a0b09;
    encBuf[2219] = 256'h0102040201080b0e0b0b08010505030301080a0c0b0b0a090801010202020201;
    encBuf[2220] = 256'h000002040502000a0e0d0b09080305040200090c0c0c0a090808000104040403;
    encBuf[2221] = 256'h0401080a0c0c0a0b09000205040202080a0c0c0a090801020100000808000103;
    encBuf[2222] = 256'h040200090b0b0b08030704030101090b0b0c0b0a090800000205040302010008;
    encBuf[2223] = 256'h090a0c0e0c0d0a09080304040302010101000008080809090c0e0d0c09080105;
    encBuf[2224] = 256'h0304010009090a09000104040302020109090b0b0d0a0b090808000000030706;
    encBuf[2225] = 256'h03040200090a0b0a0a0a090803070703040101090c0b0b0b0800040303030009;
    encBuf[2226] = 256'h0908000202000b0f0c0b0a0002040404020201080a0b0b0c0908030504020200;
    encBuf[2227] = 256'h0b0c0c0a090003040200080b0b0a00010203020304040302000a0e0c0b0a0a08;
    encBuf[2228] = 256'h0102040208090d0b0a0104050201090a0b09000000080b000307060200090b0b;
    encBuf[2229] = 256'h09020304010a0c0a0a0102080e0e0c0c090801030503030200090c0b0a090104;
    encBuf[2230] = 256'h0303000a0b0b08030502080a0c0a0908090c0d0c090804030402010800000108;
    encBuf[2231] = 256'h090d0b0b0903050302080d0c0c0b09000203040304020108090c0d0c0a080003;
    encBuf[2232] = 256'h040300090d0b0b00020503030108080800090b0f0e0b090002040302000a0b0c;
    encBuf[2233] = 256'h0908010202020304030301080b0c0b0802040303080c0e0d0b0c090002050402;
    encBuf[2234] = 256'h0108090b0a090909000001040202080c0d0c09000404040301080a0c0c0b0a08;
    encBuf[2235] = 256'h0800000101010100090a0e0d0b0a000506030401090a0b0b090808080a0c0b08;
    encBuf[2236] = 256'h0207040200080b0d0a0a08010304030301000a0c0b0b09010201080a0c0a0002;
    encBuf[2237] = 256'h0402010008020402080e0e0c0b0900030504020108080b0b0c0a0b0800040305;
    encBuf[2238] = 256'h03010109090b0b0b0c0c0a090803050301080c0d0b09090103040201080a0b0a;
    encBuf[2239] = 256'h09010504030201080b0f0d0c0b0a080105030302080b0d0b0b0a090101020101;
    encBuf[2240] = 256'h0000020405030200090c0b0c0b0c0a0a000204040300090b0e0b0b0900040505;
    encBuf[2241] = 256'h0201080b0c0a0a00010201010000010100080b0c0b0a090a0b0a00040503080c;
    encBuf[2242] = 256'h0e0b0a010405040202000a0b0e0c0a09080203040100090a0a080808090b0c0c;
    encBuf[2243] = 256'h0a0a080002030603030302080a0c0c0c0a0a080204060302080a0c0d0a090102;
    encBuf[2244] = 256'h0203000a0d0b0c09010305030201090b0b0c09000203040304010100080b0d0d;
    encBuf[2245] = 256'h0c0b0b09020604030200090b0c0a0a090809080801040405040202080b0e0b0c;
    encBuf[2246] = 256'h0908010100000008080000010101000000080800090a0c0f0b0b0a0802020009;
    encBuf[2247] = 256'h0c0b080305050302020201090f0d0b0d0908010304040201000a0b0c0b000205;
    encBuf[2248] = 256'h0303080b0e0b0a08020503040200080b0c0a0900010301080a0b080307040201;
    encBuf[2249] = 256'h08090a0b0b0d0b0a0802060403030008090a0c0a0a090003060402000a0c0c0a;
    encBuf[2250] = 256'h0901010200090a0a0002050403030200080b0c0c0a0900030401080b0e0b0a00;
    encBuf[2251] = 256'h020404020200010800010000080c0e0c0c0a0a0003060302010a0b0c09000306;
    encBuf[2252] = 256'h03020108080a090a0d0c0b0b0902060304020009090b0b0c0a08020504020108;
    encBuf[2253] = 256'h0a0909010101080b0b0a0206040300090d0b0c0909000203040403040202080b;
    encBuf[2254] = 256'h0c0c0900020301090c0a0805060301080b0d0b0901020302080a0c0b0b090005;
    encBuf[2255] = 256'h050503030100090a0b0a09010305040301090b0d0b0a080305040200080a0a0a;
    encBuf[2256] = 256'h09010305030302010000090b0d0a090507040302080a0b0b0802040201090a09;
    encBuf[2257] = 256'h0003050301090d0c0a0a01040305030102000a0b0f0c0b0a0004040402010800;
    encBuf[2258] = 256'h090809090b0a0b09000108090a0903070504020000000800080a0a0a09010201;
    encBuf[2259] = 256'h080c0c0a020504010a0e0c0a01030603020000080808090a0b0b080505030208;
    encBuf[2260] = 256'h0a0a0900030400090c0c0a080205020100090a0b0b0a0a090a01030704030008;
    encBuf[2261] = 256'h0c0b08000306020108090a090a0c0c0b0c0a090a0908020706030302090b0d0b;
    encBuf[2262] = 256'h0a08010205020401000b0d0c0b090104050301080b0c0c0a000104020300090a;
    encBuf[2263] = 256'h0c0a0a090203040402000a0c0c09000306030208090c0b0b0a08080002020201;
    encBuf[2264] = 256'h080a0c0c0b0909010405030400080c0c0c0b09080203050302000a0e0b0c0900;
    encBuf[2265] = 256'h02040201000a0a0c0c0a0909000104040303000b0f0e0a09080203030208090c;
    encBuf[2266] = 256'h0a0a09090809000204050201080b0c0c0b0a0a0908010504030201090a0d0a0b;
    encBuf[2267] = 256'h0a0a0909010203010a0f0e0b09080204040201090a0d0a0b0800020403030208;
    encBuf[2268] = 256'h0b0d0c0b0a0908000000080a0b0d0a090000020108090c0b0a09020704040208;
    encBuf[2269] = 256'h090d0c0b0a0901030402000a0d0d0b0a0002040301080a0d0b0a090800010203;
    encBuf[2270] = 256'h04030108090b0b090a0a0c0e0c0a090002030401090b0d0b0b09080204020201;
    encBuf[2271] = 256'h090a0b0c0b090b0b090b0b0a0c0a0102070501090c0f0d0a0a09010305040201;
    encBuf[2272] = 256'h080a0c0b0a08010303030101080a0c0c0c0c0a090002030502010a0e0c0c0a09;
    encBuf[2273] = 256'h01030503030100090a0a0a0b0a000307040301080b0c0b0909000a0c0b0b0803;
    encBuf[2274] = 256'h040302080908010303090d0d0b0a0105040403010100000008080a0e0b0c0a09;
    encBuf[2275] = 256'h00020303000a0d0d0a080105050201000a0a090a090000000303050401010809;
    encBuf[2276] = 256'h080809090a0b0a0204060300090b0e0a00020504020100080802010201090b0c;
    encBuf[2277] = 256'h0d0b0b0e0a0a010506030301090b0a0a08010101010103050303010809080800;
    encBuf[2278] = 256'h01080802030502090c0d0d0b0c0c0b0a010706030300090c0b09010404020208;
    encBuf[2279] = 256'h0809080001020302000b0e0c0909010303020102010301080e0d0c0a08030604;
    encBuf[2280] = 256'h020108090b0a000404040100080900010302090c0e0b080105030301080b0a0a;
    encBuf[2281] = 256'h090101000009000104040302080a08020706030200000001020401080c0d0b0a;
    encBuf[2282] = 256'h00030705020200090c0b0b09000305030108080908080001020205020100090a;
    encBuf[2283] = 256'h01040403080d0d0b09000404030201010000080009090a0a080808020200080d;
    encBuf[2284] = 256'h0e0b0b08030705030200080a0c0a0b0c09090003050603040200080b0a0b0900;
    encBuf[2285] = 256'h0000090b0d0a0901040301090c0d0a080205040200080a0a0908000101020203;
    encBuf[2286] = 256'h0502080b0c0c08020402090e0c0b0a00020403010008090b0c0c0b0900030602;
    encBuf[2287] = 256'h02010808080809090c0b080306050300000a0b0b0b0c0b0b0b00020304000a0c;
    encBuf[2288] = 256'h0b0803070302000908090a0a0d0d0a0802050301080b0d0a010406030302090c;
    encBuf[2289] = 256'h0d0c0a090001030301080a0d0a090001010100080a0800020602080b0f0c0b09;
    encBuf[2290] = 256'h0803040402020100080809090b0c0a0a080101010c0f0d0c0a09000205020201;
    encBuf[2291] = 256'h0009090a0b0a0b0a000102050202010108080c0f0c0b0b0002050401080a0d0b;
    encBuf[2292] = 256'h0908010101000a0a09080002000a0f0c0c0a0803050303010a0c0c0b09080000;
    encBuf[2293] = 256'h080b0b0b0004050401080a0d0c0a08080101010000080000000a0f0c0c0c0908;
    encBuf[2294] = 256'h02030303000b0c0b0a080203040301090b0e0b0c0a090800080102050303000c;
    encBuf[2295] = 256'h0e0d0b0a0808010101010008090a090002030400090d0a0803070300090d0d0b;
    encBuf[2296] = 256'h0a0900010100080a0d0b0b0a01010301080909000307030201000000080d0d0d;
    encBuf[2297] = 256'h0b0801050402080a0d0b0b0a0b090a08020704040200090b0c0b0b0a08020404;
    encBuf[2298] = 256'h030301090a0a090901080b0c0d0a0002040302090c0f0b0a0900020304040101;
    encBuf[2299] = 256'h00090b0b0e0b0a0908030405030301000a0b0b0a09080c0d0c0b090205050401;
    encBuf[2300] = 256'h08090c0b09090102020202030302080b0f0c0b09000204040200080a0c0b0a08;
    encBuf[2301] = 256'h03060303010a0c0b0b090004030301080a0b090004040302000a0b0c0b0d0c0c;
    encBuf[2302] = 256'h0a09030604030200090b0b0a08010305020301080a0c0c0900010202090b0e0b;
    encBuf[2303] = 256'h080104040201090b0c0b080004040302020108090a0b0a0a0107040403010009;
    encBuf[2304] = 256'h0c0c0b0a0a00000202030303020303000c0f0d0b0a0804050402020008080909;
    encBuf[2305] = 256'h0909000102040301080b0d0a0908000808010704040300090b0d0a0909000103;
    encBuf[2306] = 256'h04050402030000090a0b0a090102030100080004050401090c0a080505040108;
    encBuf[2307] = 256'h0b0a0901040402000b0d0b0900040403030201020201080b0f0c0a0900020304;
    encBuf[2308] = 256'h030202030201090b0e0c0908010304020302010100090a0b0c09000204030202;
    encBuf[2309] = 256'h020405040202080a0b0e0b0a09010605040303000a0c0c0b0800020201080802;
    encBuf[2310] = 256'h050403010a0d0b0901030302080b0d090002030503030201090c0d0b09000103;
    encBuf[2311] = 256'h01020103040300090d0d0a0908020403040100090b0b090003050200080a0901;
    encBuf[2312] = 256'h020201080903060403010a0d0c0c0a090801020201090b0b0804070502010000;
    encBuf[2313] = 256'h01020101090d0b0a0901040204010100090c0c0b0b0901020301090108000208;
    encBuf[2314] = 256'h0d0a0b0807070602020108090a0900010202000b0e0d0b0a0a08010305040202;
    encBuf[2315] = 256'h000a0c0c0b0a09080203040404040202080a0c0d0a0a0a080000020404040201;
    encBuf[2316] = 256'h090c0d0b0a090103040401080a0b0c0a0800000008080205060302090c0e0a09;
    encBuf[2317] = 256'h08010202030100090b0f0a0a09020304030109090a0b09090b0b0e0a09080204;
    encBuf[2318] = 256'h040302000b0d0c0b0a0801030200080909000000010809080b0f0f0b0b0b0801;
    encBuf[2319] = 256'h03050200090b0d0b0c0a090003050303010a0f0c0b0b080104030201080b0b0b;
    encBuf[2320] = 256'h0b090801020200080d0c0c0a0a080808000101000c0f0c0b08030503020a0d0d;
    encBuf[2321] = 256'h0a0a00010203020100080a0c0d0c0a09090001010101010108090a0a0b0b0e0f;
    encBuf[2322] = 256'h0c0d0a090104040301090c0d0a0a080102020202020301000c0e0c0b0a080101;
    encBuf[2323] = 256'h020108090b0c0a090800020102000000090c0e0d0c0a09080304030301090b0e;
    encBuf[2324] = 256'h0a0b090800000001010101090b0f0d0c0b0b0a0808010204030302090b0e0c09;
    encBuf[2325] = 256'h08010301000c0e0b0b0802050302000b0e0b0b09000001010100020100080c0e;
    encBuf[2326] = 256'h0b0d0a08080205040202090c0c0c0a080103050100080a0b0a09090008000008;
    encBuf[2327] = 256'h08000908000808080908020206050101000c0d0d0c0b0a090003040302080a0c;
    encBuf[2328] = 256'h0c090801030403030200090c0e0c0a0a08030405020008090c0b0a0900030403;
    encBuf[2329] = 256'h0200090a0c0b090b090103050502010200020301080b0f0b0908010401020504;
    encBuf[2330] = 256'h0304000a0d0d0a0908000100010103030502000009090a0a0800010504020100;
    encBuf[2331] = 256'h08010301000b0f0f09080204030201080a0b0c0c090a0104050302000a0b0d09;
    encBuf[2332] = 256'h010306040200080a0c0a09080202010008000306040300090d0c0c0908010404;
    encBuf[2333] = 256'h0202000a0c0c09080205030301080a0a0b0b08080101020203030200000a0901;
    encBuf[2334] = 256'h05060303000a0e0d0a0b080103050403030201000a0c0d0b0a00030604020100;
    encBuf[2335] = 256'h0a0a0c0a09000102040402020008090a08080000000802060404030108080908;
    encBuf[2336] = 256'h010000090c0c090105050402020009090a09010305030303010108090a0c0a08;
    encBuf[2337] = 256'h02060304030203050202000b0c0c0a080002030204050403030201090a0a0a08;
    encBuf[2338] = 256'h0104060305030100090b0b0a0802060304020008090a09000204020800090805;
    encBuf[2339] = 256'h060503040100090a0b0b0c08020405030201090b0908020502010a0c0d0a0901;
    encBuf[2340] = 256'h05030401080a0b0c09000203050303020100000a0a09090a0a0c0d0b0b0a0205;
    encBuf[2341] = 256'h0503030200090b0a0a0a01010203030106030305010b0e0c0c09010206020201;
    encBuf[2342] = 256'h090b0a0b0a00030302080d0b0b0904040301090a00010404080d0c0b09020603;
    encBuf[2343] = 256'h0302090b0d0b0b0a0900000003030203010c0c0d0b080204050200090b0c0908;
    encBuf[2344] = 256'h0001080b0c0b0c080908000103070302010a0d0c0c0a0908080202020301090c;
    encBuf[2345] = 256'h0e0b09080102020100000802090e0c0d0b09000203000b0f0b0a00030303080c;
    encBuf[2346] = 256'h0d0c0a000002020809090a09010208090f0e0b0c0a0002030302090d0d0c0a09;
    encBuf[2347] = 256'h01030301000c0b0c0a0a0808090809000001080809080001090d0f0d0b0a0901;
    encBuf[2348] = 256'h0101090b0e0b09000101090a0e0b0c090001040302080b0f0c0a0a0003050301;
    encBuf[2349] = 256'h090d0c0b0a08010201080b0c0909010100090a0b080201010a0e0b0b0908090d;
    encBuf[2350] = 256'h0e0c0b090104040300090e0b0b0a00010301080b0d0c0a0908010008090a0a00;
    encBuf[2351] = 256'h0406040201090d0c0b0a09000101000808090a090c0b0b0a00060303000b0f0b;
    encBuf[2352] = 256'h0b0803040302090c0c0b09010102000a0c0a09010301080a0e0b080901000a0e;
    encBuf[2353] = 256'h0c0b0b0802040401080a0e0a080004050100090c0b0a0802040200090d0c0b0b;
    encBuf[2354] = 256'h0908000203030404010101090a0a0d0b0a0b0a00000204030303090b0c0d0902;
    encBuf[2355] = 256'h03050400090c0d0b0b0900040202020a0a090904050302000b0c0c0a0a010103;
    encBuf[2356] = 256'h0302030208090a0f0a090a0000090c0c0c090406050301000b0e0b0a08030503;
    encBuf[2357] = 256'h0300080a090a09000a0809090102030504020202090b0b0b00060303010c0d0b;
    encBuf[2358] = 256'h0a02070404030108090b0b0b0b09010306030301080b0b0a090307040202000a;
    encBuf[2359] = 256'h0a0c09000203050108090b0901040704020208090b0b0a090800000202040402;
    encBuf[2360] = 256'h0008090106060303000a0c0c0a08010403040202080a0a0c0901030503030100;
    encBuf[2361] = 256'h0808080a090809020304040101020405040402000009090a0909000104030203;
    encBuf[2362] = 256'h030706040302090e0c0b0a0802050303020008090a0808010102030101000909;
    encBuf[2363] = 256'h0909080200090f0d0a010706050201000b0b0c0a080101020100000101020303;
    encBuf[2364] = 256'h03020000090c0c0c0a080103060304030201000a0d0b0a080206030402000909;
    encBuf[2365] = 256'h0b0a0a0901020504030302010a0a0c090002040302080b0d0c09020605040101;
    encBuf[2366] = 256'h090b0b0a09010101010809000001060303040200090b0d0b090804050302000a;
    encBuf[2367] = 256'h0c0b0b0802040503030300090c0d0c0a0800040303010009090802040301090d;
    encBuf[2368] = 256'h0d0b090802030403030100000909090c0b0d0b08010305020808080901000c0d;
    encBuf[2369] = 256'h0d0b000406050201080a0d0a0a090801020201000008090008010100090c0e0c;
    encBuf[2370] = 256'h0a09000305040202080a0b0e0a0800010200000808010202080d0e0a0a080205;
    encBuf[2371] = 256'h0302010a0d0d0b0a090802030404020008090b0b0901030501090c0e0a0a0801;
    encBuf[2372] = 256'h0102020100080a0d0c0b0b00010303010b0b0c08020402000b0e090801030301;
    encBuf[2373] = 256'h080c0d0c0c0b0a09080101000108090909000404000b0f0f0d09080203030401;
    encBuf[2374] = 256'h080a0a0a0b0909000100090e0c0b0a00020401000b0e0a080004040200080b0c;
    encBuf[2375] = 256'h0b0b0a0a0a09080307040201090c0b0b0a000008090d0c0a0902040303000a0c;
    encBuf[2376] = 256'h0c0a09080801030302080c0e0c0a0a00010303030200090c0f0b0c0a09080102;
    encBuf[2377] = 256'h0201080b0b0b0a0808010104070404010a0f0c0b0a0003050300090b0d0a0900;
    encBuf[2378] = 256'h0101000808090a0a0b0a0801060502000a0d0c0a090003040202080a0c0c0b0b;
    encBuf[2379] = 256'h090900080808080002040502010a0d0e0c0a0a08020304040200080a0c0c0b0a;
    encBuf[2380] = 256'h09000102010000000100080c0d0d0c0a0908020403030108090c0c0b0a0a0801;
    encBuf[2381] = 256'h020300090b0d09010303010d0f0c0b0a000203030200080a0c0b0d0c0b0a0803;
    encBuf[2382] = 256'h04040308090a0b0800080a0f0d0b090803060302010a0b0d0b0b090800020303;
    encBuf[2383] = 256'h0400080b0e0b0908010402020109090a0a0b0b0c0a090002040201000b0b0a0c;
    encBuf[2384] = 256'h0a090a090304050400090b0d0a000800000b0c080107070201090b0e0a0a0802;
    encBuf[2385] = 256'h02010201000300000a0f0b0a0802040301000a0801020404000a0d0e0b090104;
    encBuf[2386] = 256'h06030201080c0c0b0a080003030304020200080b0c0b0a080304050200080809;
    encBuf[2387] = 256'h00020101000a0a00010605020201080a090a0a00080206030504010000000001;
    encBuf[2388] = 256'h00080a0c0b000307060303030008090c0a090801040302030001000102050201;
    encBuf[2389] = 256'h080c0c0900050604020301010009090b0b0b09020705030301000a0b0b090004;
    encBuf[2390] = 256'h05030201000a08080204040100090b090207040502020108090a0b0a09010305;
    encBuf[2391] = 256'h0402020100080a0a0b0903070405020108090a09000204040201080808000103;
    encBuf[2392] = 256'h0403020208080a0a0900030703040403030301080a0c000407040201090c0b0a;
    encBuf[2393] = 256'h080205040304010000090b0a0a0900030404020100080908000001000a000107;
    encBuf[2394] = 256'h0704040200090b0d0a0900010402030201000108090a0c0c0b09000404020300;
    encBuf[2395] = 256'h080002020302090a0a0907040302080b0b0a090101090908020707060201080a;
    encBuf[2396] = 256'h0b0c09080001020101000901010406030101090b0908020503090c0e0c0a0001;
    encBuf[2397] = 256'h05030101080a08080001010a090a0a040403020a0f0c0a08010403040108080a;
    encBuf[2398] = 256'h0b0a0a0908000808090a020604050202080a0e0b0c0b08000103030101090a00;
    encBuf[2399] = 256'h00020302090a0d0d09080a080a0d0b0b0d090a0a0101030706020301090b0f0c;
    encBuf[2400] = 256'h0b0a080102030300090b0b0a00010202000a0a0c0d0c0c0b09080103020a0d0d;
    encBuf[2401] = 256'h0a0802050402080a0e0b0a0909010201010008090a0c090909010200090e0f0b;
    encBuf[2402] = 256'h0a0a0101020301000100090b0f0d0a09020403000a0f0c0b090003040200090a;
    encBuf[2403] = 256'h0b09000101080a0c0d0a0909080908000102020208090c0b090b0d0c0d0b0b09;
    encBuf[2404] = 256'h000201090c0e0a08020403010a0e0c0b0a0800000a0a0a0902060303000a0e0b;
    encBuf[2405] = 256'h0b0a09080808080808080c0f0c0c09080305030301090b0c0c0a0c0a0a090102;
    encBuf[2406] = 256'h04030300090c0c0c0b0b090002060303000a0d0d0b0a09000101020201010008;
    encBuf[2407] = 256'h0a0d0c0c0a0b0801030301090b0c0b000201000e0e0b0c0901020303000a0d0c;
    encBuf[2408] = 256'h0a090002030100090a0b090a0d0d0c0c0a09000403040201090b0d0b0a090801;
    encBuf[2409] = 256'h010102090c0d0c0a080102040108090b0a010203000f0d0b0b09010304020009;
    encBuf[2410] = 256'h0c0b0a090908080901030304020b0f0b0d09080801030101010a0c0c0d0b0a09;
    encBuf[2411] = 256'h0004030403000a0d0d0a080802030201000b0b0b0a080300090b0f0e09010406;
    encBuf[2412] = 256'h0201080b0d0a0a08010102010000010203030a0e0c0c090203050300090b0c0b;
    encBuf[2413] = 256'h080802020201020001020101020b0e0c0d0b08010505020300090a0a0b080101;
    encBuf[2414] = 256'h02020808010002040009080b00070504020008080a00020000000c0a01040706;
    encBuf[2415] = 256'h030202080b0c0d0a08010404030301090a0c0a090103050401010109090a0a0a;
    encBuf[2416] = 256'h000205050201000909000205040201080b0b0908020602010009090102050402;
    encBuf[2417] = 256'h02020002020100080d0c0a08040703040200080b0c0a0901040504020208090b;
    encBuf[2418] = 256'h0c0a09010304040101000001020403010a0d0c0b0901050503030100090a0a09;
    encBuf[2419] = 256'h0909090802040603040101090a0a0a08010406030301000a0a0b0a0801020101;
    encBuf[2420] = 256'h020407040303000b0c0c090104040301090a0a0900010203020205050302010a;
    encBuf[2421] = 256'h0d0a0902030402090b0b0106060302090b0d0a080306030200090b0c09090102;
    encBuf[2422] = 256'h0202010204040302080c0d0b0a080304050100090a0a080104040300080b0d0a;
    encBuf[2423] = 256'h0801030302000a0b08010505020009090a01030303090f0b0a0903040302090b;
    encBuf[2424] = 256'h0a09000704020300090a0c0c090a08020504040200090c0c0a0001040302080c;
    encBuf[2425] = 256'h0d0a0800040301000a0d0a080104040201090b0c0a0a09000900000105040302;
    encBuf[2426] = 256'h000b0d0c0b08080103030100080c0a0c0b0808000201010403040502090c0e0c;
    encBuf[2427] = 256'h0b0a08020304030300080a0b0c0c0b090001040301080a0e0a0900010100090a;
    encBuf[2428] = 256'h0901040502000b0f0b0c09000103020001090909090b090c0d090a0902010101;
    encBuf[2429] = 256'h0a0e0b0c0a000303050209090d0a090808080c0f0b0b090104040300090b0d0b;
    encBuf[2430] = 256'h080000020009090a0a00090b0c0e0b090003060202080a0b0c0b0b0b0b0c0a09;
    encBuf[2431] = 256'h0104030202000a090a0c0c0f0b0b0a0804050201090e0b0c0a0802030402080b;
    encBuf[2432] = 256'h0c0c0a0900020100080b0c0b0b0a08000002000100090b0f0d0b0c0a0a000000;
    encBuf[2433] = 256'h010108090b0c0b0c0c0b0d0b0b0908020402000a0e0b0c0a090b0b0b0a010605;
    encBuf[2434] = 256'h03010a0e0d0c090801020301080b0c0a09000100080c0c0c0909000202010009;
    encBuf[2435] = 256'h0a0a0c0b0b0d0a0a0801030300090f0d0b0c0a090002020200090d0c0b0b0900;
    encBuf[2436] = 256'h010102000a0b0f0b0c0b0a090001040302000a0f0c0b0c090900020102020009;
    encBuf[2437] = 256'h0a0e0c0b0c090800000202020201000a0f0d0b0c0a000102040100090a0c0a0a;
    encBuf[2438] = 256'h09080809000a09010001010c0e0b0c09080808080a0a080902050201000f0c0b;
    encBuf[2439] = 256'h0e0a080801010101010008080b0d0b0d0a080900030001020a0a090c0a090c09;
    encBuf[2440] = 256'h020003050a0b0d0e0a0001020500080a0f0b09090204030302090a0a0e0a0909;
    encBuf[2441] = 256'h08000102040203030808090f0a0a0c09080900040305040108090c0b0a090003;
    encBuf[2442] = 256'h0305030101000b0b0b0d09000003070202020001010801010909010b00020801;
    encBuf[2443] = 256'h0601070502030501000008090809000203060402020300010100020401020502;
    encBuf[2444] = 256'h0504020201080900010405020202010205030403010000080205040303000101;
    encBuf[2445] = 256'h0105060303020108090a09020406040402020100000808000003040405030303;
    encBuf[2446] = 256'h0100000908010205040304030403030202000008010205050303030101020204;
    encBuf[2447] = 256'h0503030404020200000808010307030502010100080000020305030502030101;
    encBuf[2448] = 256'h01080a0801010506020402020100090000000404030401080100010404020300;
    encBuf[2449] = 256'h0808000004050204020103020002000801020207040203010002020105030103;
    encBuf[2450] = 256'h020001000a03060307040102080a080909040303050200010108020109020000;
    encBuf[2451] = 256'h07030204010900080903020806010803030004010a02010807030003090c0008;
    encBuf[2452] = 256'h0b04020805020106020003080b0a0d0c00010106030102080a0a0b0d08000804;
    encBuf[2453] = 256'h030003010902000c000a0f09090904030204080d0a0a0c01010103010b080c0d;
    encBuf[2454] = 256'h08090a00090a02000a020a0f0a0b0e090808030300010b0f0e0b0a0808000301;
    encBuf[2455] = 256'h00080b0f0a0a0b09090a010009000b0e090b0b090a0b080d0c0a0a0d090a0b08;
    encBuf[2456] = 256'h090a000a0e0a0d0c0a0a0a08080a090b0d0a090a000b0d0d0c0c0a0908010100;
    encBuf[2457] = 256'h080a0e0b0d0a0a0a08080808080a0c0b0d0b0b0b0b090a09080b0e0b0d0b0b0a;
    encBuf[2458] = 256'h0909090b0b0d0c0b0c0a0a0a0a0a0b0a0b0c0c0c0c0b0b0c0b0a0b0909080008;
    encBuf[2459] = 256'h0b0f0d0c0a0b0909000008080a0b0c0c0b0c0b0c0a0a080800000a0d0c0c0b0a;
    encBuf[2460] = 256'h0a0909090a090c0b0a0c0a0a0c0b0b0c0a090a090b0e0c0b0b0c09090800090b;
    encBuf[2461] = 256'h0b0f0c090a0a000909080a0b0a0c0c0b0d0b0a0a09000800000d0c0a0d0b0909;
    encBuf[2462] = 256'h09080908080c0b0b0f0a090900020909090f0b0b0b0a000801030808000f0b0a;
    encBuf[2463] = 256'h0e0a090a08020100010b0c0b0e0a080a08010909010b09030b0a080f0f090b09;
    encBuf[2464] = 256'h02010204090a0b0e0a0000020408090a0d0b000902030808000d09010900030b;
    encBuf[2465] = 256'h0a000c01060002020a0a090e09010901040002040002040a0a080e0901000405;
    encBuf[2466] = 256'h0001020908010a00030003070801020901050002040001030901020901070002;
    encBuf[2467] = 256'h060102020800080a010601030500020201030401010209080300050602040301;
    encBuf[2468] = 256'h0102080102010307010304010102000205010403020202000303020604020204;
    encBuf[2469] = 256'h0103030104030102040102040205040203030102010001030306050303040202;
    encBuf[2470] = 256'h0100000101040503030402020202030502020100010303070403030201010001;
    encBuf[2471] = 256'h0404040202000000030605030301010809080103050402030203020402020200;
    encBuf[2472] = 256'h0102030703030402020103020305020302020304030405020202010203020504;
    encBuf[2473] = 256'h0203020100010105050305020101080900010205040204020101000801010004;
    encBuf[2474] = 256'h0302050301030302040300020200030401060202040302050100010808020304;
    encBuf[2475] = 256'h06030002000902030207020101080a00000807020204020801080a0101080501;
    encBuf[2476] = 256'h0004010103020002080b01010907030004010903010905010a02080c01000b05;
    encBuf[2477] = 256'h010005020802090c08090c02000a03020b07010802080e090a0b00080a04000a;
    encBuf[2478] = 256'h02000a04000e080c0d09090902010803090c0a0c0c08080a01090e09090c0008;
    encBuf[2479] = 256'h0a010a0d080b0c00090b080a0e090a0b080a0d080b0b090a0b090c0f090a0b08;
    encBuf[2480] = 256'h080a080b0e0a0d0b0a090b08080a080a0d0a0c0d0a0a0b09090a0a0b0d0a0b0d;
    encBuf[2481] = 256'h09090a090b0d0b0c0c0a090a00080a0a0d0d0a0b0b090a0a0a0a0c0a0b0b0b0c;
    encBuf[2482] = 256'h0e0a0c0b0a0a0a090a0b0b0d0b0a0b0d0a0b0d0a0a0a0a0a0b0c0c0c0a0b0a0a;
    encBuf[2483] = 256'h0a0b0b0b0d0a0b0d0a0b0b0c0b0b0c0b0b0a0b0a0b0d0c0b0c0a0a0a0a0a0b0d;
    encBuf[2484] = 256'h0c0b0c0a0a090a090a0b0c0c0c0b0a0a0a0b0b0c0b0c0b0a0b0a0b0c0c0b0c0b;
    encBuf[2485] = 256'h0b0a0b0b0c0b0c0c0a090b0b0c0b0d0b0b0a0909090a0b0d0c0c0b090a09080a;
    encBuf[2486] = 256'h0c0b0e0b09090800080a0b0f0b090a0801090a0a0d0b0a0b0a000a0b0a0c0b09;
    encBuf[2487] = 256'h0b0a000d0a090e09010809000d0c0a0c0900000203090b0b0f0a00000104090a;
    encBuf[2488] = 256'h0a0d0902000304080a0a0e09080802050000020900020a09080e0a0108030701;
    encBuf[2489] = 256'h01010a0a000a08030103050900020901060102030a08020c0106000204090003;
    encBuf[2490] = 256'h0902060000020b00030803070000010802060103040009090d09020106040101;
    encBuf[2491] = 256'h010a0a000801040102040800020908020a00050003070201010a0a0009020703;
    encBuf[2492] = 256'h03030809090d0900080406010102080808090003010204090901090107010403;
    encBuf[2493] = 256'h0800010909020103070303050808080b0a010106040203010909000a00050305;
    encBuf[2494] = 256'h040202000b0c0909020703040200090a09080303050301080008000403030400;
    encBuf[2495] = 256'h00000a0105030504010100000002010102020307020205020001080000020505;
    encBuf[2496] = 256'h020200090a090803070404020108000909010103040203040101020008000205;
    encBuf[2497] = 256'h0603020300000808010404040201000800010306030303010200020403050401;
    encBuf[2498] = 256'h010202010301000102030705030302080a0908030605030301080a0b09010405;
    encBuf[2499] = 256'h0402020200080000020202030301030602010402030303040302020401010302;
    encBuf[2500] = 256'h0305030403020001010307030404020000080801020404020303080900000207;
    encBuf[2501] = 256'h0403050200080909000204040202010009010102070202030300020100030003;
    encBuf[2502] = 256'h05020205020001010804020406020102010a01000005040204010809090a0404;
    encBuf[2503] = 256'h0405020108090b09000206010101000801010102020103020207020802080a09;
    encBuf[2504] = 256'h0909070301040109080909030502050108090a0c000800040108020109030109;
    encBuf[2505] = 256'h03090c01000903000003090b01080a02000c09090a03000805010b000b0f0809;
    encBuf[2506] = 256'h0a000108040009010c0f090809020208010b0f0a090a01010801080c090a0c08;
    encBuf[2507] = 256'h080b090a0b01090c080b0f090c0a08000801010a0a0e0c09090801000b0b0f0d;
    encBuf[2508] = 256'h090908010208000b0e0b0a09010100010a0d0b0d0b08080901080b090b0d0809;
    encBuf[2509] = 256'h0b080b0e09090900080b0b0f0c0a0908030200090f0c0b0a08020301010a0f0b;
    encBuf[2510] = 256'h0b0900010101080a0c0c0a09000800090a090c0e09080901080a090c09000800;
    encBuf[2511] = 256'h01090c0a0c0a090800020a0f0b0b0a0002060401080b0d0c090901020302080a;
    encBuf[2512] = 256'h0d0b0b0902040201080b0c0b0902040200080e0c0a0900020301080b0a0b0002;
    encBuf[2513] = 256'h0201090d0d0a0808020204080a0c0b0a08030503000c0c0d0b0901020402000b;
    encBuf[2514] = 256'h0e0b090800030302090a0d0b0a08000801080b0e0b0a0900030209090b0b0b08;
    encBuf[2515] = 256'h08080a090c0d0a0a080102000a0c0d0c0909020301000c0c0b0c09000001000a;
    encBuf[2516] = 256'h0e0b0c090801010200090b0f0c0a0a09010100080b0c0a0a080200090c0b0e0b;
    encBuf[2517] = 256'h09080808090c0c0a09080002010a0c0e0b0a0a08010008080b0f0b0b0a000001;
    encBuf[2518] = 256'h000a0d0c0c0900020201090c0d0d0a0908080200000a0b0b0b0b09080b09080c;
    encBuf[2519] = 256'h0a0a0a0a090b0b090b0c090a0b08090b0c0b0b08090801090c0b0f0c09090001;
    encBuf[2520] = 256'h0108080a0e0a0a0a000800080c0c0b0d0908000103080b0b0f0c090900010809;
    encBuf[2521] = 256'h090c0c090a09000a09090d09080808000c0c0b0e09000800020a0d0b0d0b0800;
    encBuf[2522] = 256'h010208090a0e0b090a09010909090e0b0a0a09020a08010d0c0b0c0900090002;
    encBuf[2523] = 256'h090b000f0b090b09080a00000b0a000c0a0a0e0b0a0a08020900000f0b090b0a;
    encBuf[2524] = 256'h01000305090b0c0f0a080800020008080d0a090a0003000a080d0a080c000408;
    encBuf[2525] = 256'h09080c0a090b08030801030a09010c09030b0b010c08020900030808080e0901;
    encBuf[2526] = 256'h0802060001000c0b000a00050201040808080a08040001040800020801060000;
    encBuf[2527] = 256'h0208090208040600020208000200050400000209010301050401020208020601;
    encBuf[2528] = 256'h0105010103000002080004040405010102080000000306030304010002000103;
    encBuf[2529] = 256'h0204030104040304040101020002030104050101020102060303040101020002;
    encBuf[2530] = 256'h0302040501020301040301030502020303040402010201020403040502010001;
    encBuf[2531] = 256'h0104020404030203000002040304030102020303050402020203030405020203;
    encBuf[2532] = 256'h0100020304040403030101020304020603030202010102000604020302000800;
    encBuf[2533] = 256'h0104030504030201010901020203040203030604020100010101040203020502;
    encBuf[2534] = 256'h0000020001060302050100080000030403050300010809020305040301010008;
    encBuf[2535] = 256'h0102040603020200090100080403010503000301010205010200010300030602;
    encBuf[2536] = 256'h0100080900010307020201000b08000006030304000b08090a01060204010908;
    encBuf[2537] = 256'h0908020402040109080a0a03030102000b00000004020002080c090809020400;
    encBuf[2538] = 256'h03080a090a0b01020204010c090a0c080101050208090b0f090800010201000a;
    encBuf[2539] = 256'h0f090800010109080a0e0a090801010102090d090a0b00000901090c0a090903;
    encBuf[2540] = 256'h0009080d0c0a0b08030202030a0f090a0b01010001080c0b0d0b00000003020b;
    encBuf[2541] = 256'h0b0b0c08000802000b090d0a090000030208090c0e080808010008000a0b0909;
    encBuf[2542] = 256'h0003090a00090d090900040108080b0e090900020100020a0d090a0902020202;
    encBuf[2543] = 256'h090d090c0a000100020109090a0b080008080809090b0b02010001010b0a0d09;
    encBuf[2544] = 256'h08080801000a0a0b0c0002030100090a0f0b0908000302000a0e0a0a0a000402;
    encBuf[2545] = 256'h08090c0c0c0a08020201000a0e0b0b08080009000b0e080909010000090d0c0a;
    encBuf[2546] = 256'h0b09000001000c0c0a0c09000809080c0c090b0c09080000080b0c0d0b0a0a08;
    encBuf[2547] = 256'h00080b0b0c0b0a0c09000a0c0b0d0b0b0b080008080a0d0c0b0a090909080c0d;
    encBuf[2548] = 256'h0b0b0b080108090a0d0c0b0b09000a090a0e0b0b0a09000809090c0d0b0b0b0b;
    encBuf[2549] = 256'h000809090a0c0d0a0a0a00090a0a0c0d0a0a00000800090f0b0a0b0900090808;
    encBuf[2550] = 256'h0c0b090c09010909080d0c090b0a080000000a0b0a0c0b080009080b0c0b0c0a;
    encBuf[2551] = 256'h01010102080c0c0b0c08090802000a090c0a08080102080b0b0c0b0b0a020301;
    encBuf[2552] = 256'h08080b0a0b0c00020908000c0b090800030201080b0c0a0a00010801010a0a01;
    encBuf[2553] = 256'h0901010100000d0a090900040201020008090909010801010b09000800020205;
    encBuf[2554] = 256'h030800080b0a010002040201010908080005020002020a090000020602020108;
    encBuf[2555] = 256'h0001000203020300080102010503030402090000080105030403000000010206;
    encBuf[2556] = 256'h0202020008010102060304020101010000030403050200020102040504020301;
    encBuf[2557] = 256'h0000080102050403020102040203060202010008000104050304020101000102;
    encBuf[2558] = 256'h0305030202010103050403040102080801020305030304020102030404040101;
    encBuf[2559] = 256'h0001080003060302030301000100010405010100000102020702010108080000;
    encBuf[2560] = 256'h0804040202010001020302000101080909080003050203000000080900000100;
    encBuf[2561] = 256'h0100000a09080204030109080a0a08000102000808090a00000800090a0a0a09;
    encBuf[2562] = 256'h01080803010908080b090b08090a0a080b0a080001000a09080c0c080a090009;
    encBuf[2563] = 256'h0a080a0d0a080909080a0a0b0b0c0a0b0a08080808090c0c0b0a0a0b09090c0b;
    encBuf[2564] = 256'h090b0800080a0c0b0c0b0b0c0b0a090a08080b0a090a0a0b0d0a0a0b0a0b0b0c;
    encBuf[2565] = 256'h08090a0b0c0b0c09090908090b0c0b0a0a080a0b0a0b0c0b0a0c0a0a09090908;
    encBuf[2566] = 256'h090a08090b0d0a0b090a0b09090a09090a0a080b0a090a0b090a0b0a0809090a;
    encBuf[2567] = 256'h090a090c090a09090a0b0a0909000008090c0c090808090908090c0908090001;
    encBuf[2568] = 256'h0009090b0a0b0c09000100080909090808090a000008090a0a08010000000908;
    encBuf[2569] = 256'h090a09000008080908010008000101080808090b000109000200080008080808;
    encBuf[2570] = 256'h04020808000b09090802040001000909080900010101010808080a0004010008;
    encBuf[2571] = 256'h0909080a0802030301090a000800000101010b0a000909020200010800090a08;
    encBuf[2572] = 256'h010801030908080b080101000100080b0a08000802030008080a090108000801;
    encBuf[2573] = 256'h00090a0800000001000808000808090202000008090a090002020101080a0001;
    encBuf[2574] = 256'h0808010001080801090a01010002030900080909010203030800080b0a000103;
    encBuf[2575] = 256'h020008080900080203030908000008080000010000080900090802040100000a;
    encBuf[2576] = 256'h09000801010203080b0a08080103010100090900000802010101000908000800;
    encBuf[2577] = 256'h00000201090808000102030001000b0a00010202030808080000010102010308;
    encBuf[2578] = 256'h0801010900030100010008000100010202040108080008020401010001090900;
    encBuf[2579] = 256'h0302020201000100020302010200000801010202020102010008010101030402;
    encBuf[2580] = 256'h0100080001030302020300090108010304020202010001010202030202000002;
    encBuf[2581] = 256'h0101010304020202020001010002040101000102030103030201030000020403;
    encBuf[2582] = 256'h0202020100020101030201030101020203040303020100010900020103040202;
    encBuf[2583] = 256'h0300090304030101010200000301020302010102000202010202000201000202;
    encBuf[2584] = 256'h0103020802000902010002020202080002000103020901000801080801010202;
    encBuf[2585] = 256'h080002000908010101010008080900000201000900080a08000002020a000008;
    encBuf[2586] = 256'h08090902080b090909080800020000000b0b080809010908010a0d0908080808;
    encBuf[2587] = 256'h08000b0b090809080809080a0a0a0b0a080909080b09080b0a09080900090b0a;
    encBuf[2588] = 256'h0b0b0a0b0a000a0b0a0b0c000009000a0b0a0e0b00090a09090a0a0d0a000a09;
    encBuf[2589] = 256'h000a0c090b0d090908090a0b0b0b0c0b0a0a090b0a0a0b0d0a0808080a0a0c0b;
    encBuf[2590] = 256'h0a0b0b0a0a0c0a0b0e09090909080a0a0b0b0b0b0c09080a0a0c0b0b0b0d0a09;
    encBuf[2591] = 256'h09080a0b0a0a0d0a080a0a090b0b0b0c0a0a0b0a0a0c0a090a09090b0a0d0a09;
    encBuf[2592] = 256'h0a0b0a0a0b08090a0b0b0a090c0a080b0b0b0a090b0c09080b0a080b0a0a0c0a;
    encBuf[2593] = 256'h00090b090a0b090b0a08090b080b0b09090c090908090908000a0b090a0a090a;
    encBuf[2594] = 256'h0908090a080a0a000a09000b09000000080b09090a09000908080b08000b0001;
    encBuf[2595] = 256'h0b0903080900000800080a00080800090908080800080201090001090a020009;
    encBuf[2596] = 256'h000800020808000800020800020800020900030801030a000308080308080200;
    encBuf[2597] = 256'h0103000102010101080001010102080002020304010002010103010302000302;
    encBuf[2598] = 256'h0808020104030002030802060101020001050000020103040003020802060001;
    encBuf[2599] = 256'h0302010401020301030302020201000402030303030302040102040202010203;
    encBuf[2600] = 256'h0302030301020402010102010303020502000203000204010103080103020302;
    encBuf[2601] = 256'h0103040201020103010801030101030301000203020202010000010202010103;
    encBuf[2602] = 256'h0102010101020101000101020202000201010102000000000001020200020201;
    encBuf[2603] = 256'h0801010001020100020100000800020008020109020200080101000001000101;
    encBuf[2604] = 256'h010908010109000800020108000109010009020008000009080800010008080a;
    encBuf[2605] = 256'h0800080800010801090a09000808090800000909000909090808080a09080908;
    encBuf[2606] = 256'h080908080a0a080908000909080a08090a08000a09090a08080a00090a09080a;
    encBuf[2607] = 256'h08090a080a0a08000a08090908090909090a000b0a080009000809090a0a090a;
    encBuf[2608] = 256'h0800080908090a09080a09090900000b09080908000b08080a090a0b01000a09;
    encBuf[2609] = 256'h0809080b0900080a08090a080a09080908090808080900090a090809090b0901;
    encBuf[2610] = 256'h080a0008090809090a08080900000809080a080800000908000a0b0000090908;
    encBuf[2611] = 256'h01020900010909080000080808090908080001010901080a0002000100010009;
    encBuf[2612] = 256'h0a08020009000200080000080101080000090101010908000101000008000001;
    encBuf[2613] = 256'h0100000808000201080801030808000809010008010200080101000008000101;
    encBuf[2614] = 256'h09000801090101000002010a0800000002000001090800090102000900000808;
    encBuf[2615] = 256'h0001000001080800000800020809000800000901010100000801000909000802;
    encBuf[2616] = 256'h080a080008000301080808000001090800080000000809000008000908000108;
    encBuf[2617] = 256'h0008090000000808080909000000000108090808090800080009000000080909;
    encBuf[2618] = 256'h0008080809000808080008090801090a0801080a00090800000808090901000a;
    encBuf[2619] = 256'h0900000800080b090009080808080000000909000901080908000a09080a0900;
    encBuf[2620] = 256'h0a09020909000800080a00010a09080808090b080009090909090808090a0101;
    encBuf[2621] = 256'h0809090909080909080b0a00080b09000809080a08000809080009080a0b0908;
    encBuf[2622] = 256'h000009090909080a08080809080009080800000a09000909000a090108080009;
    encBuf[2623] = 256'h090808000101080a0008080a0908000808080100080800000001000908000808;
    encBuf[2624] = 256'h01090b0002000009080001080801080001080800000908080800000001080800;
    encBuf[2625] = 256'h0801010909010000000008090801010900010201080800080802000900020801;
    encBuf[2626] = 256'h0009010300090001000100010200080201090002000800000102020102000002;
    encBuf[2627] = 256'h0000000202000000000001020101020201020000010100020009020200000301;
    encBuf[2628] = 256'h0101000000020001010201010801010100000000000800010202000800020001;
    encBuf[2629] = 256'h0100080808090202090901030008080001000908000900020108000000080808;
    encBuf[2630] = 256'h0a01010a0801090101080102000a080908080908000100090808080002010009;
    encBuf[2631] = 256'h09080801000000000001080900000908000908000802010001010001090a0101;
    encBuf[2632] = 256'h0900080001000800000800000000010908000000000008000809080808020809;
    encBuf[2633] = 256'h000800010001080808000a0a090800020900080a080009090808000a0a090108;
    encBuf[2634] = 256'h00090902080909090900090b09090a09080800000008080a0a0a0b0801090900;
    encBuf[2635] = 256'h0809080908000800080a090a0a00080808080909000101000900090a080a0c00;
    encBuf[2636] = 256'h000101010908010808080a000109090809080302090908080800080000080009;
    encBuf[2637] = 256'h0a08010100080001080908000908000900080000080900000809080908000909;
    encBuf[2638] = 256'h000001000008000909080008000800090a090a09090109010100010908000808;
    encBuf[2639] = 256'h0008090800080000090a08080908000001000801080808000901000808000000;
    encBuf[2640] = 256'h0802010808010800080800080901080901010800010100010100010800000800;
    encBuf[2641] = 256'h0301080801080908080000020301080101000008080009000208000301000200;
    encBuf[2642] = 256'h0a00000900000001010800000000000008080000000100080101080800000900;
    encBuf[2643] = 256'h010009080001000901010200000808080908010001080800080b080000020000;
    encBuf[2644] = 256'h020201010a080109080809000100020300080100080109090000080000000000;
    encBuf[2645] = 256'h0108010201020108010201080001000809080101080802000900000002000203;
    encBuf[2646] = 256'h0100010000000000010909010101000800020108090808080001000800010101;
    encBuf[2647] = 256'h0003010908000a08080900000001010800000808000908000008080801080908;
    encBuf[2648] = 256'h0100090801080108090808000800080908080800080808000800010109000100;
    encBuf[2649] = 256'h08090a08000900090b0801000000000100080008000900000000010808080909;
    encBuf[2650] = 256'h0809090001000808090800010008080002000a08000908000100000101080808;
    encBuf[2651] = 256'h080b090a090a0900000001020200010100090908090a0a090808090008000108;
    encBuf[2652] = 256'h0001020908090a090a090008080900000a08080a0002080801080b09090a0008;
    encBuf[2653] = 256'h0000010000090b0a0a08080a000108000809090a0a0a08090801000809010000;
    encBuf[2654] = 256'h0808000909090a0800090900090900090b090808000100010008000809090b08;
    encBuf[2655] = 256'h080909000900010900010008000a0a090a09080001000001010809080a090808;
    encBuf[2656] = 256'h000800090009090800080001000809080a0909080801000001020a0800090908;
    encBuf[2657] = 256'h090a080809090001000102000800080a010a0900000900000a09090809080908;
    encBuf[2658] = 256'h0800080002010101000008090908090a080000000100080b0909080908000101;
    encBuf[2659] = 256'h0100090009080200000301080008090908090801020008000809090909000009;
    encBuf[2660] = 256'h0202010303020302010100090b0c090a090801030203040201010008090a0900;
    encBuf[2661] = 256'h0000010302020302000008090b0a0a090a010304030201030200000808090009;
    encBuf[2662] = 256'h0909080801020203010108090b0c0a0a090003040403020202000a0b0b0c0909;
    encBuf[2663] = 256'h0800010204010000080a0b0a0a090801010402030303010101080a0a0a0b090a;
    encBuf[2664] = 256'h0a09010103040403030100090c0b0c0a0a010103040303030200080909080800;
    encBuf[2665] = 256'h0203040201000a0c0b0c0b0b0902030604040302010008090b0c0c0a0a090800;
    encBuf[2666] = 256'h010104040204030203020808090d0b0c0a0a090901040202020100080a080002;
    encBuf[2667] = 256'h030404040200000a0c0d0b0d0b090901040305030301000a0c0b0c0a08080002;
    encBuf[2668] = 256'h0103030000090909080901010100080a0a0c0b0b08010403040301080a0b0b0c;
    encBuf[2669] = 256'h0b0908000003030201000a0c0b0c0a00030703040201090c0d0d0a0a0a000103;
    encBuf[2670] = 256'h050402030100090a0c0d0a0b0909080001020202020203020301000a0d0c0b0b;
    encBuf[2671] = 256'h0c0a08080908080a0a0a0b0c0a0903050506040202000a0c0d0c0c0a0a080001;
    encBuf[2672] = 256'h030403030201000a0b0b0d0a0a0808010008090b0c0c0b090002040502030200;
    encBuf[2673] = 256'h090a0b0d0b0c0a090a0908080a08090802060503050201080b0e0c0c0a0a0800;
    encBuf[2674] = 256'h01040304020100090b0d0c0a0a08000204040201000a0a0c0b0b0a0800010203;
    encBuf[2675] = 256'h030208090b0b09080205030303090e0c0d0b0b0b090002030502020100080808;
    encBuf[2676] = 256'h000207020303000a0f0d0c0c0a0a08000205030402010008080a090000020201;
    encBuf[2677] = 256'h080d0f0b0d0b0a080004040503030201080a0b0c0c0a0a090800000001020202;
    encBuf[2678] = 256'h04030404020201000b0c0d0c0b0a090001030502030101080a09080802050403;
    encBuf[2679] = 256'h0201080c0d0c0b0b0a0900040404030402020100090a0b0d0a0a0a0800020304;
    encBuf[2680] = 256'h0303020108080a0a0a0a0801030704040503030301000b0f0c0c0a0b09080205;
    encBuf[2681] = 256'h040303030208090c0b0a0a08020504040200080a0e0b0c0b0908010306040302;
    encBuf[2682] = 256'h030108080a0c0b0b0b0b0b0a0a000003050504040303020200090c0c0c0c0a0a;
    encBuf[2683] = 256'h09080102030403030201000808000101020300090d0e0c0c0b0a0a0801030504;
    encBuf[2684] = 256'h04020202010108080a0a0c0b0d0b0c0b0a0900030505030502010108090b0c0b;
    encBuf[2685] = 256'h0b0b0a0800010203030402030302030202080a0d0e0b0c0b0a09000204030302;
    encBuf[2686] = 256'h0208090b0c0b0a0a09020306040303030200090b0d0d0c0b0c0b0c0a09080001;
    encBuf[2687] = 256'h0304030503040303030201090c0c0d0c0b0c0b0b0c0a0a080002040505030403;
    encBuf[2688] = 256'h020208090c0d0c0b0b0a0a0900020403040202020008080a0a0b0a0b0b0b0a0b;
    encBuf[2689] = 256'h0b0a0a0a00020605040403030201000a0c0d0d0c0b0c0b0b0908010405040403;
    encBuf[2690] = 256'h020301000a0b0e0b0d0a0a0a0900010103030304010101080908090001020302;
    encBuf[2691] = 256'h01090d0e0c0c0b0b0b090001040304030201080a0a0c0a0a0003050504030101;
    encBuf[2692] = 256'h080b0e0c0b0c0b0b0a080002050304030302010008090a0b0b0a0a0908010100;
    encBuf[2693] = 256'h080c0d0e0b0c0b0a0800030405040303030201090b0d0c0b0a09080204040402;
    encBuf[2694] = 256'h01000a0c0e0c0b0b0b090802040603050203010108090b0c0c0c0a0a09080001;
    encBuf[2695] = 256'h02030303020000090a0a090908010206040303040100080a0c0c0c0b0b0a0b0a;
    encBuf[2696] = 256'h09080001020303020304030504040503030403020200090c0e0c0d0b0c0b0a0b;
    encBuf[2697] = 256'h09080203070305030303030100090c0c0c0b0b0c0a0808000103030303020108;
    encBuf[2698] = 256'h0a0b0a0a000406040404020200090c0c0c0c0b0a0a0901010404030302020009;
    encBuf[2699] = 256'h0a0b0c0a0a080103060402030208090c0c0d0b0b0b0a08010205030403020100;
    encBuf[2700] = 256'h08090a0a0a080001040304030201090c0d0d0b0c0c0a0a0a0800010404040404;
    encBuf[2701] = 256'h0203020200090a0c0d0b0c0a0b09090000020303040202000008090800020505;
    encBuf[2702] = 256'h04030202010a0d0d0c0c0b0b0b090802030604030302020109090c0b0c0b0a08;
    encBuf[2703] = 256'h00020305030202080a0e0c0c0b0a0a0900030604030402020108090b0c0c0b0b;
    encBuf[2704] = 256'h0a090001030304030200080b0d0c0b0a0a00020504040402030100090b0d0c0b;
    encBuf[2705] = 256'h0c0a09080002030503020101090a0c0b0c0a08000204040403020200080b0c0c;
    encBuf[2706] = 256'h0c0b0a0b090900020305030402020100090a0a0b0b0908020404040202000a0d;
    encBuf[2707] = 256'h0c0d0b0b0b0a000103060304030303020101080a0b0e0c0c0b0b0c0a09080104;
    encBuf[2708] = 256'h04030503020108080b0b0d0a0908000305030301000a0d0d0c0c0a0a08000205;
    encBuf[2709] = 256'h040304020200080a0c0c0b0c0a0908010204040303020108090c0c0c0b0b0a09;
    encBuf[2710] = 256'h000205040304020000090b0c0c0a0a090001040403040201000a0c0c0c0b0c09;
    encBuf[2711] = 256'h0900010305030403020108090a0c0c0b0b0a09080202050303030208090d0b0d;
    encBuf[2712] = 256'h0a0a09010204040402020009090c0c0b0a0b090801020503040302010108080a;
    encBuf[2713] = 256'h0c0b0b0c0b0b0b0909000104040305020202000809090b090908010103020208;
    encBuf[2714] = 256'h0b0f0c0c0c0b0b0a090002040505030402020208090c0d0b0d0a0b0a09000304;
    encBuf[2715] = 256'h06030403020108090c0c0c0b0a0a09080203040304020108090b0b0b0b090803;
    encBuf[2716] = 256'h04050402030100090a0d0b0d0b0a0b0908000304040403020200080b0c0c0a0b;
    encBuf[2717] = 256'h09080104030502020008090b0d0a0b090900030305030200090b0d0c0c0a0909;
    encBuf[2718] = 256'h00010303040403040303030201000a0c0e0c0c0b0b0b0b090001040403040303;
    encBuf[2719] = 256'h02010008090b0b0d0a0b0b0a0a000103060304020201080a0c0b0c0b0a080102;
    
    encBuf[2720] = 256'h040302000a0d0c0c0b0a09080102040504030503020200080a0c0c0b0b0b0b0b;
    encBuf[2721] = 256'h0a0a0900010403030302000a0c0d0a0a00050506040304020208090d0c0c0b0b;
    encBuf[2722] = 256'h0b09080204040403020200080b0d0b0c0b090900020304040203030202010809;
    encBuf[2723] = 256'h0b0f0b0c0b0b090900010302030202000809090b09000406050403030201090b;
    encBuf[2724] = 256'h0f0c0b0c0b0a08000305040402020208090b0c0c0c0a0a0a0808010304040403;
    encBuf[2725] = 256'h03030100090a0c0c0c0a0b09090801020403040200080a0c0c0b0b0a09000206;
    encBuf[2726] = 256'h04040303030108090d0c0b0c0b0a09080203050403040101080a0d0c0b0b0b0a;
    encBuf[2727] = 256'h00010306040303020208090b0d0b0c0a0a0801030403030301090b0d0d0b0b0b;
    encBuf[2728] = 256'h0908010504040304020108090a0c0c0b0c0a0908000304040402020108090b0c;
    encBuf[2729] = 256'h0c0a0b0908000102040202010009090b0a09080305050403020201080a0d0d0b;
    encBuf[2730] = 256'h0c0c0a0a09080002030504030303020201090a0d0d0b0b0c0909010103050303;
    encBuf[2731] = 256'h020201090a0d0b0d0a0a09090001020202020304020303020101080a0c0c0d0b;
    encBuf[2732] = 256'h0b0b0a09010304030301080a0c0c0a0800030703030200090d0d0c0a0b090802;
    encBuf[2733] = 256'h04050503030201080a0d0c0c0b0a09080003040304030200080a0c0d0c0a0b09;
    encBuf[2734] = 256'h00010404040402030100090b0c0d0b0a0b080801010303020201080909090900;
    encBuf[2735] = 256'h02050503040301080a0c0d0c0b0a0a0001030404020200080a0b0c0c0b0a0908;
    encBuf[2736] = 256'h010504030403020100090b0c0c0c0a0b09080102040203010101000000000809;
    encBuf[2737] = 256'h0b0a0c090a080a0c0c0d0b0b0a01040704040402010008090c0b0b0c0a090808;
    encBuf[2738] = 256'h00010102020203030402020100090b0e0c0c0a0b080003050503030401010808;
    encBuf[2739] = 256'h0b0c0c0c0a0b0a0909090908080003060505030304020108090c0b0c0b0b0a08;
    encBuf[2740] = 256'h000103020200090b0d0c0a090103070404030201080a0c0c0c0a0b0908010305;
    encBuf[2741] = 256'h0304020108090c0b0b0b090002040304020100090a0c0d0b0a0a090002050304;
    encBuf[2742] = 256'h040202020000090b0d0d0b0b0a0b09080203050503030302080a0d0c0b0b0a09;
    encBuf[2743] = 256'h0003050403020208090b0b0c0a09090909090a08000204050303020100080909;
    encBuf[2744] = 256'h0a090801030503000b0f0f0d0b0b0a08020405040403020200090c0c0c0c0a0a;
    encBuf[2745] = 256'h09080001030304030203010201010100080b0c0e0b0c0b0a090a090909080801;
    encBuf[2746] = 256'h0404050304030303030200080b0e0d0c0b0b0b09090102030503030302010808;
    encBuf[2747] = 256'h0909000800090d0e0d0b0c0a09000306040303030100090b0d0b0c0a0a090900;
    encBuf[2748] = 256'h0001010202010809090004060504030301080a0d0c0c0b0b0a0a080002030403;
    encBuf[2749] = 256'h0402030303030301090d0d0c0c0b0a09080101020301010008080a0908010407;
    encBuf[2750] = 256'h050404020301000b0f0c0c0b0b0b09000203060303030302010000090a0c0c0b;
    encBuf[2751] = 256'h0b0c0a0a0a0900010204030303030202020200080a0c0d0b0b09000204020009;
    encBuf[2752] = 256'h0b0e0b0a00020405030300090b0e0b0b0a080801020304050404030302080a0d;
    encBuf[2753] = 256'h0e0b0c0b0b09000204050402030100080a0b0a0a0a09080a0a0c0c0b0b090801;
    encBuf[2754] = 256'h040504050303040101090b0d0c0b0b08080303050202080a0c0d0b0a0a000104;
    encBuf[2755] = 256'h040403030100080a0c0b0c0a0a08080103030504020301090b0f0c0c0a0a0900;
    encBuf[2756] = 256'h02030504020302010100080a0c0d0b0b0b0a0a08000102030402030302030203;
    encBuf[2757] = 256'h0304030201000b0f0d0c0b0b0c0a09080801030404040303020108090a0b0901;
    encBuf[2758] = 256'h020403010a0f0d0c0b0a0a09000001020304030504030203020100080a0b0e0c;
    encBuf[2759] = 256'h0c0c0a0b090900000202030503030303030108090a0b0a0b0a0b0b0c0b0b0a00;
    encBuf[2760] = 256'h04050402010b0e0d0b0c090900020203040305040304030200090c0c0c0c0b0a;
    encBuf[2761] = 256'h0b0909000103040403030100080809000102030402020101080a0f0d0d0c0c0a;
    encBuf[2762] = 256'h0b0900010304030503020303020201080a0c0d0b0c0b0c0a0b0b0a0908010406;
    encBuf[2763] = 256'h0403030401010008090a0c0b0c0b0a0a0900020204030302020100090b0e0c0b;
    encBuf[2764] = 256'h0c09000104040302020201000108080a0e0c0d0b0b0b0a080001040305030304;
    encBuf[2765] = 256'h0302020108090c0d0b0c0b0b0b0a0a08010405040304020100080a0b0c0b0c0b;
    encBuf[2766] = 256'h0a090003060403030301090a0c0c0b0c0b0b0a0a090104050404020301010809;
    encBuf[2767] = 256'h0a0b0b0c0a0b0a0b0a090a080801020604040402030100090b0b0b0a09000000;
    encBuf[2768] = 256'h090d0c0c0b090003050403030108090c0b0c0b0b0a00030704040202000a0b0c;
    encBuf[2769] = 256'h0c0b090900020202030100090a0b0b09020705040202010a0c0d0c0a0a080001;
    encBuf[2770] = 256'h0203030402010200080a0c0c0d0a0b0908030504040301010a0b0d0c0b0a0900;
    encBuf[2771] = 256'h0104030502020109090c0b0a0a090000020302010100080a0909080405050302;
    encBuf[2772] = 256'h000c0d0d0c0a09080103050403020100090b0c0c0a0b09090001010203040303;
    encBuf[2773] = 256'h03030100090a0c0c0b0a0b0b0a0a0a0c0a0b0a080407050503040201080a0c0c;
    encBuf[2774] = 256'h0c0b0a0a090002030405020302020000090a0c0c0c0b0b0b0908000204040403;
    encBuf[2775] = 256'h0203030101090a0c0d0b0c0b0b0a090800030505030403030100080b0d0d0c0b;
    encBuf[2776] = 256'h0b0a09000205040403030101080a0b0c0b0c0a0a0a0900000202040203010202;
    encBuf[2777] = 256'h010304030401080b0e0d0c0b0b0a080103060304020100090c0b0b0c09080102;
    encBuf[2778] = 256'h030203030202020302000a0f0c0c0c0a0a090808010203040403040303020108;
    encBuf[2779] = 256'h080a0c0d0c0c0b0c0a09080203050403030200080b0c0b0c0a09000204050303;
    encBuf[2780] = 256'h00080b0d0d0b0a0908000303030303010000010101000108090a0a0b0b0d0b0a;
    encBuf[2781] = 256'h0b0b0c0c0d0d0c0b0a09020507030403030108090c0b0c0b0a0b090900000204;
    encBuf[2782] = 256'h03040304010100090a0c0c0b0d0b0b09080306040502030201080a0b0c0d0b0c;
    encBuf[2783] = 256'h0b0a090801030405030203020100080a0b0d0b0b0a090001030201080c0c0b0c;
    encBuf[2784] = 256'h09000205030403020100080a0a0c0b0a08080101020108090a0b0a0800000a0f;
    encBuf[2785] = 256'h0f0e0b0a08010406040303030300000a0c0d0c0c0b0c0a0a0808020306040304;
    encBuf[2786] = 256'h03020100090c0c0c0b0b0b09090101040304030302020008090a0c0b0c0a0b0a;
    encBuf[2787] = 256'h09090000020305040303030101080a0b0c0c0b0b0c0a0b0b0900010504040402;
    encBuf[2788] = 256'h02020108090a0b0b0b0a090008090d0d0d0b0c09000206030502020100090b0b;
    encBuf[2789] = 256'h0b0b0b0a0800020403020201090b0e0c0b0b0a09000206040403040201000a0b;
    encBuf[2790] = 256'h0d0b0c0a0a0809000000010204030404030202010100090c0e0c0d0b0c090900;
    encBuf[2791] = 256'h0204040403030101080a0a0d0b0b0b0b0a080801020203030403030303020202;
    encBuf[2792] = 256'h0305040302000c0f0e0c0b0b0a09000203060303040102000008080a0a0c0c0b;
    encBuf[2793] = 256'h0c0b0a0a0800020306040303020200080a0a0b0b0c0b0b0c0b0b0a0900030504;
    encBuf[2794] = 256'h04040303030201080b0f0b0c0b0a0a0808010203020402040303040200080b0e;
    encBuf[2795] = 256'h0b0d0b0a0908010304030401010809090a090001020302000b0e0d0b0a0a0908;
    encBuf[2796] = 256'h0002020306040403040301080b0e0c0c0a0b0908000305040402020108090c0c;
    encBuf[2797] = 256'h0b0b0b090801030403030303010200000808090a0a0c0d0d0c0c0a0a09010306;
    encBuf[2798] = 256'h03030302010008090b0b0c0b0a0b0b090802060403030208090b0d0b0c0b0a09;
    encBuf[2799] = 256'h01030504030201080b0c0a0a00040603040100090b0d0b0d0b0a0b0a08010505;
    encBuf[2800] = 256'h03040302010000090a0c0b0d0b0b0c09090101030403040303030302000a0c0d;
    encBuf[2801] = 256'h0c0c0b0a0a0908010303040304030303020200090b0d0c0b0c0b0c0b0b0a0801;
    encBuf[2802] = 256'h040504030203020201080a0c0d0c0b0b0a0a000102050304030202020100090c;
    encBuf[2803] = 256'h0c0c0c0b0b0a0a09090101040405040305020201080a0b0e0b0b0b0a0a080001;
    encBuf[2804] = 256'h020302020101010305050305020108090c0c0b0b0b0b0a090900020404040402;
    encBuf[2805] = 256'h020208080a0b0a0a090a0b0d0c0b0a0a000104050304030503030302000c0d0d;
    encBuf[2806] = 256'h0b0c0b0b0a0908020405050203020108080a090b0a0c0a0c0a0c0a0a09000306;
    encBuf[2807] = 256'h04040303010108090c0b0d0b0a0b090800010303040303030302020108090b0c;
    encBuf[2808] = 256'h0b0b0c0a0b0b0d0c0b0b0a000306030303010103050202080b0e0a0a08000102;
    encBuf[2809] = 256'h010301080c0f0c0b0b080002020403030201080a0b0b0901030504030402000b;
    encBuf[2810] = 256'h0e0c0b09000101080b0d0a08000301000a0900030704030304030201090b0e0b;
    encBuf[2811] = 256'h0c0a0b0c0b0b0a0901040305030403030301090a0b0d0c0a0a0908020303000a;
    encBuf[2812] = 256'h0c0d0a0a08000304040302000009000000080c0d0b09010403010b0f0c0b0a09;
    encBuf[2813] = 256'h09000106050403020108090a0a0b0c0b0c0a0b09080808010303040203030404;
    encBuf[2814] = 256'h0303010103070502010c0e0d0b0a090800010202030402020000090909090909;
    encBuf[2815] = 256'h0001020300080b0d0c0b0b0c0a09020504030108090a0b0c0b0c0b0902050502;
    encBuf[2816] = 256'h03010203050303020a0d0d0e0b0b0c09080102040302010203040201080b0d0b;
    encBuf[2817] = 256'h0c0b0b0b0c090104060305020201000a0c0d0b0c0b0a09000103050403030202;
    encBuf[2818] = 256'h0100090b0d0c0b0a090909090a08010505040203010009090c0b0c0b0a090800;
    encBuf[2819] = 256'h01030503040301010800080b0d0c0d0a09080102020304030401080c0c0b0a00;
    encBuf[2820] = 256'h0102010201030302090f0c0b0b090001030505050202080a0c0c0a0b09090a08;
    encBuf[2821] = 256'h0104050303020101010008090c0c0c0a09080809080000010000080800030505;
    encBuf[2822] = 256'h0304030302000b0d0c0a080100090d0c0b0b000102020103060504030301000a;
    encBuf[2823] = 256'h0c0d0c0b0a0a0900010304040303020009090a0909080808010304010b0f0d0a;
    encBuf[2824] = 256'h080001000a0a09020505030202030101080c0d0a090801010a0c0c0a09000108;
    encBuf[2825] = 256'h090902060504030202000008090a0b0c0b0b0d0b0c0908020403030303030402;
    encBuf[2826] = 256'h02080a0a0d0c0c0e0b0b0a0004050303030203030302080c0f0b0c0b0b0b0900;
    encBuf[2827] = 256'h010304040305020202080a0c0c0a0909090908010504040201080a0a0b0c0d0b;
    encBuf[2828] = 256'h0b08010504030301010100000a0c0b0d0a0a0a0a090003060303020100010108;
    encBuf[2829] = 256'h0b0f0b0b090102030301020200090c0e0b0a090103030503050302080b0d0b0a;
    encBuf[2830] = 256'h0900000909080102010b0f0e09010304030009080003050202080908090a0f0c;
    encBuf[2831] = 256'h0c0b0a080801030505040301000a0c0b0b0a090b090901060403020008090000;
    encBuf[2832] = 256'h00090a0b0a08000a0f0d0b0b0103070202010000000008090b0c0a090a0a0a0a;
    encBuf[2833] = 256'h09000304040304030303000b0e0d0c0b0b0908010304040404030401010a0c0c;
    encBuf[2834] = 256'h0c0b0b0a0a090801030504030303030301080b0d0d0b0b0c0a09090102020302;
    encBuf[2835] = 256'h030403050201000a0a0a090b0e0c0d0b0908010303030303060302000b0e0d0b;
    encBuf[2836] = 256'h0a0a080002040404030100090a0c0b0a0a0a0908010101010101020304010000;
    encBuf[2837] = 256'h00030402080f0c0b0b0a0a0c0c0b0a08030504030403030100090c0a0b0a0b0d;
    encBuf[2838] = 256'h0d0a090103060200080809090a0b0c080106040301000b0b0d0b0c0b0a090003;
    encBuf[2839] = 256'h0504020102030301000a0d0c0a0a0b0c0b0c090103050201000000020202090b;
    encBuf[2840] = 256'h0c0a090808090b0a0801020b0f0d0a090205030301080009090c0b0b08040703;
    encBuf[2841] = 256'h02000909090a0d0d0b0c090800010000000206040303020201000a0d0d0b0b0b;
    encBuf[2842] = 256'h0b0c0b0b0a01060503040203010200090a0e0b0c0a0b09080808010203040402;
    encBuf[2843] = 256'h020008080001080008000102010b0f0f0b0a0909090800040405020000000203;
    encBuf[2844] = 256'h02000b0f0c0a080000080a0900010301090b0b010706040200000909090b0b0c;
    encBuf[2845] = 256'h0c0909010202030101010203030302020102000a0f0e0b0c0a0a090a0a0a0006;
    encBuf[2846] = 256'h060404010100090808090b0c0c0a090002020201020204030300090b0b0b0b0e;
    encBuf[2847] = 256'h0c0b08020504020008000101080c0d0b09020603020008000101000c0f0b0b00;
    encBuf[2848] = 256'h0305030200080808090a0d0b0a00030603020200000a0c0c0a0a000101010103;
    encBuf[2849] = 256'h0704040108090b0a090a0e0d0b09020504030101020101090c0f0b0a08000200;
    encBuf[2850] = 256'h010103070201090c0c0a080002010002030603010a0b0e0a0908080900000305;
    encBuf[2851] = 256'h03020109080800000a0d0c0b09000203020102030404010a0c0d0a0801020108;
    encBuf[2852] = 256'h090104050400090c0b0a080201080a0a00050402000b0c090204030200000000;
    encBuf[2853] = 256'h080c0f0c0a0900010201010205030401080a09080101000b0d0d0b0b0a0a0900;
    encBuf[2854] = 256'h0205050404030200080b0b0b0b0b0b0c0a090002030303030305030202010001;
    encBuf[2855] = 256'h080c0c0c0a00030502000a0c0c0d0b0c0a09010305040303030302080c0c0c0a;
    encBuf[2856] = 256'h080809090b0900030602080b0b0804060401080b0b08040402090d0d0a090102;
    encBuf[2857] = 256'h0100090801050401080a0a0a080108090a090002040201010201090f0f0a0a00;
    encBuf[2858] = 256'h030403010008000100080c0d0b0a08020303010a0b0a000502080d0d0a080404;
    encBuf[2859] = 256'h040200010001000a0f0f0b0a08010202020202040402000b0c0c09080008090a;
    encBuf[2860] = 256'h09030504010a0c0c0a00010108080105060302080a0c0a0008080b0e0b090001;
    encBuf[2861] = 256'h0202010205040302080a0b0b0a0a0a0b0a00030503000a0e0c0a090000010100;
    encBuf[2862] = 256'h010506040302000a0b0b0a0a0c0e0c0b0900020304020304050201090c0c0b0b;
    encBuf[2863] = 256'h0a0908020405030301090b0c0b0b0a0b0a080206040302000809000201080d0e;
    encBuf[2864] = 256'h0b0a08010000080004050402080a0a0b090900090909010303000b0b0a01010a;
    encBuf[2865] = 256'h0f0f0a010505030208090a09090a0c0e0a0a00030303010008020403000c0d0b;
    encBuf[2866] = 256'h090001000b0902070703080b0d0b0901000a0d0b0005060302080a090801000a;
    encBuf[2867] = 256'h0f0b0b00020402080908020403000d0c0a08010301080908020602080c0b0a08;
    encBuf[2868] = 256'h0200090d0b00040502000909000204000c0c0b080203020a0c0a00050400090c;
    encBuf[2869] = 256'h0b08010301090b0903070401090b0a080100080d0c0a00030401080900020403;
    encBuf[2870] = 256'h080b0c0b0800090b0c0b02060402000909080000090d0b0a010503010a0b0a01;
    encBuf[2871] = 256'h0504000a0c0b080102010a0a0903060301090b0a0102010a0f0d090002020009;
    encBuf[2872] = 256'h0800020401090b0b000502000b0d0a02050401090b0b0a08080b0e0b0a000504;
    encBuf[2873] = 256'h030303020302080d0d0c0a09090808000002040202080800010203000c0e0b09;
    encBuf[2874] = 256'h0802040202020201080c0e0c0b0b0a09000204060402010009080809090b0c0a;
    encBuf[2875] = 256'h08020303090d0b09010303080a0b0007040201080900030501090d0d0b0a0808;
    encBuf[2876] = 256'h0100010306040201080a0c0b0b090001040502030100080b0d0c0b0909000202;
    encBuf[2877] = 256'h020305040402080a0c0c0a0808000909000406040201090b0c09090008090800;
    encBuf[2878] = 256'h0307030100090b0b0a09090a09090206050303020100090a0c0c0c0a0a080102;
    encBuf[2879] = 256'h030304030302080b0c0c090001020304030403000a0d0d0a0900000008080104;
    encBuf[2880] = 256'h060201090b0a0803060201090a000102000a0c0a010504010a0e0b0a01020402;
    encBuf[2881] = 256'h0102020202080b0c0b08030503030301000b0f0f0c0908010201020103050402;
    encBuf[2882] = 256'h01090b0b0b0908080b0b0901050504020200080b0d0c0b0b0901020505040304;
    encBuf[2883] = 256'h02080a0c0d0a0a08080000020305040208090a0b08010100090c0a0001040201;
    encBuf[2884] = 256'h0801020502000c0c0b0b0a08000104040403020009080008090b0f0a09010302;
    encBuf[2885] = 256'h080a080207060301080a0c0c0b0a0b09000306040303020100090b0e0c0a0a08;
    encBuf[2886] = 256'h000203020302030100090c0c0a08090a0a0b01070503030009080801080d0d0d;
    encBuf[2887] = 256'h0a0901030301000101040302080c0d0a0a0800000000020305040201090c0c0c;
    encBuf[2888] = 256'h0b0a090002050304020108090b0b0c0a0a08020305030108080a080a0b0d0d0a;
    encBuf[2889] = 256'h08010202000002070403020a0c0c0a09090a0b0b080605040208090b0b0b090b;
    encBuf[2890] = 256'h0c09000407030301090a0a0a0b0c0b0b09010306020100080808090a0a0a0a09;
    encBuf[2891] = 256'h090a0b0b010707040201090b0c0c0b0b0b0908040504030208090a0b0b0b0d0b;
    encBuf[2892] = 256'h0900020603030009090a0909090a0c0c0a0900010304030201080a0b0c0d0c0b;
    encBuf[2893] = 256'h0b09020704030200090b0a0c0b0d0c0b0a080105040303020208090c0c0c0a0b;
    encBuf[2894] = 256'h0a090900020504040201080a0b0c0c0a0b090800040404030201090b0c0d0b0a;
    encBuf[2895] = 256'h0a080802020403040200080c0b0b0b0900000008000103040300090e0c0c0b0a;
    encBuf[2896] = 256'h080103040303020000090c0d0b0d0a08080808080103060303080c0b0b090809;
    encBuf[2897] = 256'h0b0c09010603010b0d0b000305010b0e0b0902030400080a000202000d0f0b09;
    encBuf[2898] = 256'h080102010100020302000a0e0c0a090909080002040303000a090002000c0f0f;
    encBuf[2899] = 256'h0a090102020101010102000a0f0d0908020301080a0b0a0102080b0c0a030705;
    encBuf[2900] = 256'h01000a0b0908090a0e0a090106030301000909090b0d0c0a0801030302000801;
    encBuf[2901] = 256'h0101000b0d0b09000108080801060302090c0c090101010a0e0b000307050008;
    encBuf[2902] = 256'h090a090800090a0b0903070502000a0a0b0b090000010103030403040201090d;
    encBuf[2903] = 256'h0d0c0a080204020200000800000a0c0c090005050200090a09000101080b0a08;
    encBuf[2904] = 256'h010503000a0a08050503010a0b0b01050302090c0a01050402080a0e0a080802;
    encBuf[2905] = 256'h0201030404040201080a0b0c0a0b090a090802040605030302010909090b0a0c;
    encBuf[2906] = 256'h0b090005040301000001040401090d0c0a0801030101020405040200090a0b09;
    encBuf[2907] = 256'h0809090b0a0105060303030100080a0b0b0a000406030401010000080b0d0c0b;
    encBuf[2908] = 256'h0a01050503030101000009090a0c0a0802050402010008000800000a0b0b0903;
    encBuf[2909] = 256'h07070303020100090a0b0d0b0a0900030505040202000809090b0a090a080004;
    encBuf[2910] = 256'h050602030108090a090808090800010304010100090206040402000008090808;
    encBuf[2911] = 256'h0b09080105030101080805050303010a080102060209090b0904050302000b0a;
    encBuf[2912] = 256'h0a0a030404040303050208090c0e0a0908030403030201030201000d0e0b0908;
    encBuf[2913] = 256'h01020000080006040303000a08000103080f0d0c0b0800020203040404030208;
    encBuf[2914] = 256'h0c0d0c0a09080801020306030202080b0d0b0b0b0a0b08000406040202010800;
    encBuf[2915] = 256'h0a0b0d0c0c09090001030303040302000b0e0c0a0a090801000203050203000a;
    encBuf[2916] = 256'h0b0d0c090a0900080101020102010800090b08080a090d0d0a0a0a080b0b0909;
    encBuf[2917] = 256'h00050108090a09040402080c0f0a0a0a0a0b0d090001040100090b0c090a0b0a;
    encBuf[2918] = 256'h0c0b080000020008080809080e0e0c0c0c0a0a090908010203040401080b0e0c;
    encBuf[2919] = 256'h0a0a090a090a0a09020202080b0f0a0a08090a0c0b0a0900000909080802020c;
    encBuf[2920] = 256'h0f0f0b0c0a0b090908010305030308090a0e0b0b0d0a0a09000200080a0c0c0a;
    encBuf[2921] = 256'h09080100020202010a0f0d0b0b090909090b0b0a00010302080a0e0b0b0d0c0b;
    encBuf[2922] = 256'h0c0b0a0a0003030503000b0d0c0c0a0a0c0a0b08010202010b0e0a0908000809;
    encBuf[2923] = 256'h00010704010a0e0d0b0b0a08000800030404040200090c0c0a0b0b0a0a080802;
    encBuf[2924] = 256'h0404030302000a0a0e0c0b0c0a090800030303030202000b0d0b0b0a08090c0c;
    encBuf[2925] = 256'h0d0a000204030009090908080b0e0b0b0005030302000000000a0e0f0c0a0900;
    encBuf[2926] = 256'h010101020202040201080a0a0b0c0a0a0a0b0b0f0a090903070403030101080a;
    encBuf[2927] = 256'h0c0c0d0b0a09000304040302020100090a0d0c0a0b0a00000203030405020303;
    encBuf[2928] = 256'h00090a0e0a0a0a09000801010101040103040202030203040009090d0b0a0c0c;
    encBuf[2929] = 256'h0b0b08060405030201010908080b0b0a0a01070203030000000a0a0b0e090002;
    encBuf[2930] = 256'h0604020202010302080a0d0d0a09090102040405030302080a0c0c0a09080001;
    encBuf[2931] = 256'h0203070303030100090a0a0909080a0b0a090004070304040204020100090b0b;
    encBuf[2932] = 256'h0808010108090808060404020200010303030400000800020200000909010503;
    encBuf[2933] = 256'h0403040605030302000001010101090c0c0a0104040403040404020208090a0a;
    encBuf[2934] = 256'h0a0a08080103070504020301000008090a0a0a08010305030403020203030402;
    encBuf[2935] = 256'h02010101040402010a0d0c090804060402030001000000010001000800010800;
    encBuf[2936] = 256'h010802050407030203020203030302080c0a0908040300010800070602040301;
    encBuf[2937] = 256'h01010001010a08090c09080005060204020101010000000b0908000503010000;
    encBuf[2938] = 256'h0006040202000900020205020908090901080c0a08000707020203010302080a;
    encBuf[2939] = 256'h0e0d0a0908020203030301010009010102070300080b0f0a0a09080100030404;
    encBuf[2940] = 256'h040200000a0a090808030100020a0f0b0d0c08000104030304030001000a0b0c;
    encBuf[2941] = 256'h0e0a0a0b090801040203030201020109000b0e0b0d0d0a090902020204020102;
    encBuf[2942] = 256'h000a0a0c0d0a0a0b080809010109080b0e000304070100090a0c0b0b0d0a0a09;
    encBuf[2943] = 256'h010100010809010303070109000a0d0a0c0d0b0b0a0808000303030601080a0c;
    encBuf[2944] = 256'h0c090909080a0c0a0909000009090c0c090a0a01010204000d0c0d0c090a0a09;
    encBuf[2945] = 256'h0a0a09000005020101090b0a0d0e0c0c0b0b090801020001010203010a0d0e0c;
    encBuf[2946] = 256'h0b0a0908090b0a0c0b09000103040101080b0d0c0c0c0b0b0a0a09090a0b0b0a;
    encBuf[2947] = 256'h0a010104060302000d0e0d0b0c0a0a0900010204030200090b0c0d0b0c0b0a0a;
    encBuf[2948] = 256'h080103040201000b0c0d0b0b0b090909090800000201000a0e0d0c0c0b0a0908;
    encBuf[2949] = 256'h0103040200080b0f0b0c0b0b0a0a080103040301000b0e0b0c0a090909090909;
    encBuf[2950] = 256'h080808080a0c0b0d0b0a0c0a08090002010102090d0d0e0c0c0a0a0800010201;
    encBuf[2951] = 256'h02030100090e0d0b0c0a0a090908010205030301080b0c0d0b0a0b0b0b0b0900;
    encBuf[2952] = 256'h01020702030300080b0f0c0a0a0901000101000000090b0b0d0a090a08020003;
    encBuf[2953] = 256'h060101080d0c0a0a00030100000b0b090b0a000b08040003060808030b09080f;
    encBuf[2954] = 256'h0c080801040800010b01070100010c0b0a0a0901090806010405010001080001;
    encBuf[2955] = 256'h0a0a090f0b080a08020104060202010908000801030809010b000509090a0f0c;
    encBuf[2956] = 256'h08090307020403020101090b0b0e0b0b0b08020306050203030100080d0c0b0b;
    encBuf[2957] = 256'h0a080104040304020202000a0b0d0c0a0908010303040302030208090b0d0b08;
    encBuf[2958] = 256'h090205020404020101090b0b0e0a090900030307030402030000090b0d0a0b09;
    encBuf[2959] = 256'h01020504030101090908090a080a08060405030201000908090a0b0a0b080204;
    encBuf[2960] = 256'h04040203040304010008090908000800030506040302020008080a0b0d0b0a00;
    encBuf[2961] = 256'h010405040306020302010008090a0a0a0b090908030306040204030403040201;
    encBuf[2962] = 256'h000909090908020101030405040302020102010008090b080507050303030102;
    encBuf[2963] = 256'h0101000a0c0c0a00020503040302020101080801030504040203020202000809;
    encBuf[2964] = 256'h0b090801010101040606050303030101020100000a090a090403030302010306;
    encBuf[2965] = 256'h03050201030305050402030108090c0c0a0a0901040306040302030001080a0a;
    encBuf[2966] = 256'h090c090a09020503070303030100080a0c0a0a0b090102070402040201010108;
    encBuf[2967] = 256'h08090a0808080000090003050703020201010202010108080001080302000604;
    encBuf[2968] = 256'h0103030006040304010800000803020908090a05050307020203020000090c08;
    encBuf[2969] = 256'h090903040204020802010805030204030003020103020806030004020900090f;
    encBuf[2970] = 256'h09090a01030507030205020101080a0a0c0a08000003010103030204000b0800;
    encBuf[2971] = 256'h0207050102010803010801090d01010005010a080a0e09080a01020207040204;
    encBuf[2972] = 256'h030102000a0a0d0c0a0b0c09080902030405030001000901010801080d0a0b0c;
    encBuf[2973] = 256'h08090c090a0a02020204000a00080a03080b030208070408080c0f0a0c0c0a0a;
    encBuf[2974] = 256'h0a08000802030205020102010a080d0d0b0c0c0a090a08090a08080801080a00;
    encBuf[2975] = 256'h090902020004000b0c0f0f0b0c0c0a090a080800020100000a0b0b0b0c080909;
    encBuf[2976] = 256'h08090a0a0f0f0b0c0c0a0a0a09090800000103030200090d0c0d0c0c0a0b0b0a;
    encBuf[2977] = 256'h0908000800080a0a0b0e0b0c0b0b0a0909090808080a0b0f0d0c0c0b0b0c0b0a;
    encBuf[2978] = 256'h09080101030101080a0c0e0c0b0c0a0b090909090a090a0b0d0b0c0b0b0b0a09;
    encBuf[2979] = 256'h090908090c0c0b0c0b0c0c0c0c0c0a0a0a0a090908000002080a0e0d0d0a0b0a;
    encBuf[2980] = 256'h09090800000100080b0e0e0b0b0b0a09090001000102090b0d0f0b0b0b0b0908;
    encBuf[2981] = 256'h00010101000b0c0c0e0c0a0c0a090800010100010808080c0d0b0d0b09090800;
    encBuf[2982] = 256'h0808000a09000c0d0a0d0b080a08010808020808020b0c0a0e0b0a0c0b080b0a;
    encBuf[2983] = 256'h000c09080b0b000d09000a0105010104090a090f0b090d0b090b090102020500;
    encBuf[2984] = 256'h00010801020909010d09020a0a090f0b080b0801090206000205080001090105;
    encBuf[2985] = 256'h0001030800020d09090d0a080b08040105050102020102030001010b08040801;
    encBuf[2986] = 256'h04090a000d09020901070102050203060102020000010908010a09000c080208;
    encBuf[2987] = 256'h0207000304030406020202010102080001080a000c0901090004000307040404;
    encBuf[2988] = 256'h0201020101010001010801040102040008080a0a010804070404030304030202;
    encBuf[2989] = 256'h0208000008000108000200030702030401030702040302020200010201010201;
    encBuf[2990] = 256'h01040203040100000902060404050303040302020201000909090a0002040404;
    encBuf[2991] = 256'h0202050303040101010003040305030203040202000a0a090901040307040403;
    encBuf[2992] = 256'h0303020108080808000103070504030302010108090a0a0a0802070503040303;
    encBuf[2993] = 256'h020101090909090802050503030303020001090a080103070403040203030202;
    encBuf[2994] = 256'h0201000204040402000008090000000403030707020303020302000201010303;
    encBuf[2995] = 256'h0203020004030307030104040304040203030206020303040102020101000900;
    encBuf[2996] = 256'h080004040307030305020204020102010103010102010801080a000808040404;
    encBuf[2997] = 256'h07030205030203020101000801090b090b0d0008090100090703030603020402;
    encBuf[2998] = 256'h0204020102010800080b0a0b0f00090903040207040204030103020102010902;
    encBuf[2999] = 256'h000003030005010802020107020207030305030304030103010801090a08090a;
    encBuf[3000] = 256'h02030107050204030203020103030104030104030103010a000a0f08090a0103;
    encBuf[3001] = 256'h0107050104020002000808090b08090a01010902000b02090f00080b02010a04;
    encBuf[3002] = 256'h010a02080f080c0e0a0b0e0a0b0b0b0a0c09090900080900090c0a0e0c0b0d0c;
    encBuf[3003] = 256'h0a0b0c0a0a0a0a0b0c0b0b0d0b0b0c0b0b0b0a090a090a0b0c0d0c0c0c0b0c0b;
    encBuf[3004] = 256'h0c0a0b0a090a0a0a0a0a0b0b0d0b0b0c0b0b0a0b0b0a0a0b0c0b0d0b0d0c0b0b;
    encBuf[3005] = 256'h0c0a0b09090908010000010a0b0e0c0c0b0c0a0a0a09080908080a0b0c0d0c0a;
    encBuf[3006] = 256'h0c0b090a0a080808000a0d0b0e0d0a0c0b0b0b0b090a0a000909090d0b0c0d0c;
    encBuf[3007] = 256'h0a0c0a0a0b0a090b0a0b0c0d0a0c0b0b0b0c09090900080001090a0a0f0b0b0d;
    encBuf[3008] = 256'h0b0a0c0a090909080808010908000908020802060102050001010a0c090e0a0a;
    encBuf[3009] = 256'h0b09000901050202050102030101030001050003050101030800000c0b0a0f0a;
    encBuf[3010] = 256'h090a000201040502040401020208000008000100040503050403040402040302;
    encBuf[3011] = 256'h0403030403020402030304030503030603030503030403030403040203020402;
    encBuf[3012] = 256'h0202030204020304030305030304030305020303030403030303030303020101;
    encBuf[3013] = 256'h0800090a0a0a0a000000050302040108090e0e0b0d0c0b0c0b0a0b0b0b0b0c0b;
    encBuf[3014] = 256'h0b0d0b0c0c0b0b0c0b0a0c0a0a0b0b0c0c0b0d0b0b0c0a0b0a0a080908000809;
    encBuf[3015] = 256'h080b0c0d0b0d0b0b0b0b0a0a0909080008080800080000030405040304030303;
    encBuf[3016] = 256'h010009090c0b0b0a0802040605030304020100090a0b0e0c0a0b0b0a0b090809;
    encBuf[3017] = 256'h08000a0a0a0e0c0a0d0c0a0b0c0a0c0a0b0b0c0b0c0c0a0c0a0b0b0b0a0b0a0a;
    encBuf[3018] = 256'h0a0a090b0b0c0d0b0c0c0b0b0b0c090a08000001020103020101010908010903;
    encBuf[3019] = 256'h0704050503050403030503030403030303030401020200000008080809090008;
    encBuf[3020] = 256'h02040405050304040203030302030100080b0c0c0d0b0b0d0a0a0a0a08080800;
    encBuf[3021] = 256'h080a0a0e0b0d0b0c0b0a0a0908000201030202010809090b0a09080801000a0b;
    encBuf[3022] = 256'h0f0f0e0b0b090903070605040404030304030202010000080908090000020305;
    encBuf[3023] = 256'h0403030402030203040305030504030303040201020008080809080001020403;
    encBuf[3024] = 256'h04020100090d0c0c0c0b0a0b090801020204030200000a0d0c0c0c0b0c0b0a0c;
    encBuf[3025] = 256'h0b0b0c0c0b0c0b0c0b0b0b0a09090000030203030200000a0d0b0c0b0b0b0b0a;
    encBuf[3026] = 256'h0a0b0a0d0c0c0c0c0a0b0b090800040404050304030302030202020201030302;
    encBuf[3027] = 256'h0503030402020202000800090001020506030603030403030302020101010008;
    encBuf[3028] = 256'h08090b0c0d0c0d0b0c0c0b0b0b0b0a09000103040304020100090b0d0c0d0b0b;
    encBuf[3029] = 256'h0b0b0b0c0a0a0a0b0b0d0c0b0b0b0c0b0a090a0808000800080809090a080900;
    encBuf[3030] = 256'h020403050100090d0e0c0d0b0b0b0b0900010404050304030201010009090b0b;
    encBuf[3031] = 256'h0b0c0b0a0a0a090a0c0b0d0c0c0c0a0b0b0b090a0808000000080a0a0d0c0b0d;
    encBuf[3032] = 256'h0b0a0b0b0b0e0b0c0d0c0b0c0c0a0c0a0a09090900080101010008080a0c0b0b;
    encBuf[3033] = 256'h0d0a090a08010001020200020909000a00050306050305030302030000080a0a;
    encBuf[3034] = 256'h090b00020104060102030809080c0b080a00060206030202020a0d0c0e0c0b0b;
    encBuf[3035] = 256'h0c090a0900000103010101080a0c0c0c0b0b0b090a08010000000b0c0d0d0b0c;
    encBuf[3036] = 256'h0b0b0a0a090809080a0c0b0b0a02070707040404030503030303010200080a0a;
    encBuf[3037] = 256'h0b0b0a0a09010304050403040203030304030404030404020302030101080809;
    encBuf[3038] = 256'h0909080801020304030200090c0d0d0b0b0c0a08080203050402030201080b0d;
    encBuf[3039] = 256'h0c0d0b0c0b0c0a0b0a0b0b0c0b0b0c0b0b0a0b0a0a0808010101020100090a0d;
    encBuf[3040] = 256'h0c0c0c0b0c0b0b0b0d0b0b0c0b0c0b0b0a0a0900010504040404030304020201;
    encBuf[3041] = 256'h0101000800080808010002020304030403030403040403050304040304030402;
    encBuf[3042] = 256'h030302030102000809090b0d0b0b0d0a0b0b0a0b090900000203050304020301;
    encBuf[3043] = 256'h00090b0f0b0e0b0c0b0c0b0b0b0b0b0c0b0b0b0b0b0c0a0b0b090a0800000203;
    encBuf[3044] = 256'h030304020100090a0c0d0c0c0c0b0c0c0b0b0c0b0a0a0a080001040404040303;
    encBuf[3045] = 256'h03030302010000080909090809000000010108090a0d0b0c0c0b090900030605;
    encBuf[3046] = 256'h04040404030303020201080a0d0d0c0c0c0b0b0c0a0a0a0a0908080001000000;
    encBuf[3047] = 256'h0809090b0b0c0b0a0a0908080000080a0c0f0c0c0c0c0c0b0b0a0c0a08090002;
    encBuf[3048] = 256'h030406030404030303030303020102000008090a0a0c0c0b0d0b0b0c0a0a0900;
    encBuf[3049] = 256'h020305050304040202020001080909090b0b0b0c0c0b0d0b0c0d0a0b0c0a0a09;
    encBuf[3050] = 256'h09000001020202020108080a0b0d0b0d0b0b0b0d0b0c0c0b0b0d0a0b0a0a0a09;
    encBuf[3051] = 256'h090809090909000407070406040404030403040202020008080a0b0b0c0b0a09;
    encBuf[3052] = 256'h0801020404030402030201030204030404030303030200000a0b0c0c0c0a0909;
    encBuf[3053] = 256'h0801020303040200080a0b0d0b0b0a08010305040301000a0d0e0c0d0b0c0b0b;
    encBuf[3054] = 256'h0b0b0b0b0c0a0b0b0b0b0d0a0a0a0a08000002020102090a0e0d0c0c0c0b0b0b;
    encBuf[3055] = 256'h0b0b0a0a0a0a0a0a0a0b0a0a09010406050503050303030302020008090a0b0b;
    encBuf[3056] = 256'h0b0b0a0000030503050402030404020403040403030403020301010100080809;
    encBuf[3057] = 256'h0800000202030202010a0c0e0d0b0b0c0a09080103050304020208090c0d0c0c;
    encBuf[3058] = 256'h0b0c0b0b0a0a0a090a090a0a0b0c0b0b0b0a0a0801020402040101090a0e0c0c;
    encBuf[3059] = 256'h0b0c0b0a0b0b0a0a0b0b0b0c0b0b0a09010306050503030402020100090a0b0d;
    encBuf[3060] = 256'h0b0b0a0909000103030203020101010104060405040304030302020108080a0b;
    encBuf[3061] = 256'h0a0a0908080001080b0d0f0c0b0d0b0b0a0a09000104030304020100080b0d0b;
    encBuf[3062] = 256'h0d0a0b0a0a09090809090a0b0c0c0b0b090a0802030406020203030204030404;
    encBuf[3063] = 256'h04040303030200090b0f0d0b0c0c0a0a09090800010202040101010009090b0b;
    encBuf[3064] = 256'h0c0c0b0b0c0c0b0c0b0c0b0c0a0a0909080001010101080a0b0f0c0b0c0b0b0b;
    encBuf[3065] = 256'h0b0a0b0a0a0b0c0b0e0b0c0c0b0b0c0a0a090002070504050404040304030402;
    encBuf[3066] = 256'h0201010008090a0b0a0b09090003050405030303030402020203030305020402;
    encBuf[3067] = 256'h0302010108080a0b0d0b0a090002030504030303020000090b0a0c0b090b0a0a;
    encBuf[3068] = 256'h0c0c0d0d0d0b0c0c0b0c0a0b0a0a0a090a090a0a0b0b0c0b0b0b0b0b0b0a0b0c;
    encBuf[3069] = 256'h0b0d0d0b0d0c0b0c0b0b0b0c0a090a0909080808080000010203050404030404;
    encBuf[3070] = 256'h0202020101000809090a09080103060504050304040303040203030303040202;
    encBuf[3071] = 256'h020201010000080a0a0b0c0a0a0801060504050304040202020000090a0b0d0b;
    encBuf[3072] = 256'h0c0b0a0a0a0909090a090b0b0c0b0b0b0b0901010404030301080b0f0d0c0b0c;
    encBuf[3073] = 256'h0c0a0a0a09080908080808090a0a0b0a0a0a080101020300000b0f0c0d0b0d0a;
    encBuf[3074] = 256'h0b0a090a0909090a0c0b0c0b0c0a09000205050403040302020108090a0c0b0b;
    encBuf[3075] = 256'h0c0a0a090a09090a0b0c0b0c0a0a080803050404040302020100090b0c0b0d0b;
    encBuf[3076] = 256'h0b0c0a0b0b0c0a0d0a0b0b0b09090004040503050203010100090b0b0d0b0b0b;
    encBuf[3077] = 256'h0b08090101010202010001000103040604040303030302080a0a0e0b0b0d0b0a;
    encBuf[3078] = 256'h0b0a0a0c0b0b0c0c090b0a08080002010203090b0d0f0d0b0d0b0a0c090a0908;
    encBuf[3079] = 256'h00080808090a0b0c0c0b0b0a0a0a080909090a0c0c0b0d0a0909000101050303;
    encBuf[3080] = 256'h070404060405040503040304030302010108090b0c0a0b0b0800020504040403;
    encBuf[3081] = 256'h03040201020001010102020303040101080b0c0d0b0c0a0a0900010305030403;
    encBuf[3082] = 256'h0202010009090b0a0c0a0a0a0c0b0c0e0b0c0c0c0b0a0b0b090a080908080a0a;
    encBuf[3083] = 256'h0c0c0c0b0c0b0b090a080900080a0a0d0d0c0c0b0b0c0a0a0908000801000008;
    encBuf[3084] = 256'h09090b0a0a080205050504030303020201080809090900020405040304030302;
    encBuf[3085] = 256'h0304030404040403040402020202010008000000020304050303030201080b0c;
    encBuf[3086] = 256'h0c0c0b0b0a090002030403030200090c0d0b0d0b0b0b0b0a0c0b0b0d0c0c0b0c;
    encBuf[3087] = 256'h0b0a0b090900010103030200000b0e0c0c0b0b0b0b0a0a090a0a0c0b0d0c0b0c;
    encBuf[3088] = 256'h0a0a0a0001020403040302020008090b0b0b0a0a0800010001000a0b0d0c0909;
    encBuf[3089] = 256'h0005040604020304010000080a0a0b0a09090802020203000b0c0f0b0c0b0a08;
    encBuf[3090] = 256'h000203050202080a0e0d0d0b0c0b0b0b0b090a0a090b0c0b0c0b0c0a09080103;
    encBuf[3091] = 256'h06030502030100080a0b0e0a0b0a0a0808000101010108080809020704050503;
    encBuf[3092] = 256'h0503020101080a0b0e0b0b0c0a0a080801020203020100090b090b0a01020407;
    encBuf[3093] = 256'h020201090d0c0e0b0c0b0b0b09080002030403020108090b0c0b0b0a09080001;
    encBuf[3094] = 256'h080c0d0e0d0b0d0b0a0a08000204050304030202030304050404050304040203;
    encBuf[3095] = 256'h020000090a0c0b0c0a0a08020404050304030302020100080008080801010100;
    encBuf[3096] = 256'h01080a0b0d0c0a0b0a0003070403040402010108080a0a0c0a0b0c0a0a0b0c0b;
    encBuf[3097] = 256'h0d0b0b0d0a0a0a0808010203020301090c0e0c0d0b0c0a0b0a0a0a0908080908;
    encBuf[3098] = 256'h090a0a0a0b0a090808010100080b0f0d0b0d0b0b0a0908010305040303030302;
    encBuf[3099] = 256'h02010102040305040304030201010809090a0801030706030503040302020200;
    encBuf[3100] = 256'h01080808000102040504030403020100080b0c0c0c0a0b0a0808020404030402;
    encBuf[3101] = 256'h0201080a0d0c0b0d0a0b0b0a0a0a080900080808080809080a0909090a0c0c0c;
    encBuf[3102] = 256'h0c0c0c0b0c0b0c0a0b0b0a0b0b0b0a0a090001040604040303030300090c0d0d;
    encBuf[3103] = 256'h0b0d0a0b0a0a090801020304040303030303040201010008090c0d0b0d0b0c0b;
    encBuf[3104] = 256'h0a0a0a0000020305040303030402020302010100090c0c0d0c0c0b0c0b0a0a09;
    encBuf[3105] = 256'h080102050304030203010100090b0b0b0d0a0b0a0a0b0a0b0b0b0c0b0a080003;
    encBuf[3106] = 256'h06050403050203030202000108080a0a0b0c0b0c0b0b0c090908010404050403;
    encBuf[3107] = 256'h0304020100090a0b0e0b0b0c0a090908010000020800090b0b0c0c0a09090003;
    encBuf[3108] = 256'h0303050100080c0c0d0b0c0b0b0b090a09080a090a0b0c0b0b0a080005040504;
    encBuf[3109] = 256'h030305030505040404050304030403020100080a0c0b0c0a0a09010305060304;
    encBuf[3110] = 256'h030303020200000808080908080800000809080a090800040604050403030401;
    encBuf[3111] = 256'h020008090a0c0b0c0b0c0a0c0a0a0c0a0a0b0a0908000103040202000a0f0c0d;
    encBuf[3112] = 256'h0c0b0d0a0b0a0a0909080000000000080809090a0a0b0b0d0c0c0c0c0b0c0b0a;
    encBuf[3113] = 256'h0b0a0900010205040303030402010201000100000008090a0a0b0c0a08010705;
    encBuf[3114] = 256'h05040404030303040201020000000908090a09090a0908080104040505030404;
    encBuf[3115] = 256'h0203020100080a0b0d0b0c0b0b0a0a0a090909090a0a0a0b0b0b0b0a09090808;
    encBuf[3116] = 256'h0a0b0e0e0c0c0d0b0c0b0c0b0b0b0a0b0a09080002020403040201000a0c0e0c;
    encBuf[3117] = 256'h0c0b0c0a0a0a0808010304030403030201000809090b0b0b0c0b0a0a09090001;
    encBuf[3118] = 256'h050404040404020303020201010808080a09080a09090a0c0b0c0c0a0b0a0000;
    encBuf[3119] = 256'h0405040304020200090b0e0d0b0c0b0c0a0b0a0a0a0908000102030504020302;
    encBuf[3120] = 256'h0108090e0c0b0d0b0c0a0a09090801010203040404020304030203020101080a;
    encBuf[3121] = 256'h0a0c0c0b0b0b0909000303060403040303030304030303030301090a0f0e0b0d;
    encBuf[3122] = 256'h0c0b0b0b0a09080102040502030401010009090b0c0c0b0c0b0b0b0b0a090908;
    encBuf[3123] = 256'h0001010000080c0c0c0c0b0b0b00010605030504020303030304030603050304;
    encBuf[3124] = 256'h0302020108090c0b0c0b09080206040404030402010100080809080908000100;
    encBuf[3125] = 256'h020001000000010205050405030304020100080a0b0d0b0b0b0b0a0b0a090b0c;
    encBuf[3126] = 256'h0b0d0b0a0b090801020302000b0f0f0d0c0b0c0b0b0b090a0800000101010808;
    encBuf[3127] = 256'h0a0b0c0c0b0c0b0b0c0c0b0c0b0c0a0a0908010204040304020201000809090a;
    encBuf[3128] = 256'h0a09080102030304020202040405040603050303040202010000090909080001;
    encBuf[3129] = 256'h04050404030403040202010200000809090a0b0b0b0a0a090002040504030304;
    encBuf[3130] = 256'h0101000a0b0d0d0b0c0c0a0b0b0b0b0a0a0a090909080008000809090c0e0c0c;
    encBuf[3131] = 256'h0c0b0c0c0b0a0b0a09090908000001000008090a0b0e0b0d0c0b0b0c0b0a0a09;
    encBuf[3132] = 256'h0800020304030403020101010008000908090a0b0d0c0c0b0b0a080105060404;
    encBuf[3133] = 256'h04040203030302010100080a0a0d0b0c0b0b0b0a090001030405030304010200;
    encBuf[3134] = 256'h080a0c0c0c0c0b0b0b0b0a090001030404020200090b0e0c0b0c0b0b090a0808;
    encBuf[3135] = 256'h0000010102010102040204040203040202020008090d0b0d0b0d0a0a0a080002;
    encBuf[3136] = 256'h040404040203020108080a0c0b0d0b0a0a0a0800010304030403030401030303;
    encBuf[3137] = 256'h03050100090c0e0b0d0c0a0b09090000010101000b0c0d0c0c0b0a0a09080202;
    encBuf[3138] = 256'h05040304030304040204040305040404030402030101090a0c0c0b0a09000307;
    encBuf[3139] = 256'h0404040203020100080a0a0a0a0a090900020103040204030305030403030202;
    encBuf[3140] = 256'h00080a0b0d0c0a0a0a080001020102000a0b0f0b0c0b0a0a090808090a0d0e0d;
    encBuf[3141] = 256'h0c0c0c0b0b0a0b0909080000010100000a0b0c0d0c0b0c0b0c0b0c0a0b0a090a;
    encBuf[3142] = 256'h0001020404040203020008090c0c0c0b0b0a0900010305040304020302010201;
    encBuf[3143] = 256'h0202030303020303010304050505040403030403010100090809080002040603;
    encBuf[3144] = 256'h030402010009090b0c0a0a0a000003030403030101090a0e0b0e0b0c0b0c0b0c;
    encBuf[3145] = 256'h0a0a0a09080001010001090b0d0e0c0c0b0c0b0a0a0908080102010200090b0e;
    encBuf[3146] = 256'h0c0c0c0b0a0a0a0908000102030402020100090b0d0c0c0c0b0a0b0908010305;
    encBuf[3147] = 256'h04040303030201080a0b0c0b0b0a090103060404030304030102000008080a0a;
    encBuf[3148] = 256'h0a0a0a0800020504050303030300080b0d0d0b0b0b0909000204040402020108;
    encBuf[3149] = 256'h0b0c0e0b0c0b0b0b0a09000101030304020000080a0c0b0e0b0b0b0b0b0c0909;
    encBuf[3150] = 256'h080003050503050303020200090b0e0b0d0b0a0a08000205040303030200080b;
    encBuf[3151] = 256'h0c0c0c0a0a090800020303050303030303030401020008090b0d0c0c0b0b0a0a;
    encBuf[3152] = 256'h080801010201010109090c0d0b0d0c0b0c0c0b0a0a0901040504040303030201;
    encBuf[3153] = 256'h010305060504050304020200090a0d0c0a0b0908020505040303030101080a0a;
    encBuf[3154] = 256'h0c0b0a0a0908010203040304030403040303020200080a0c0c0b0c0909080202;
    encBuf[3155] = 256'h040304010100090a0a0c0b0b0b0a0a0a0b0b0d0c0c0c0c0b0c0c0a0a0b0a090a;
    encBuf[3156] = 256'h0809080809090b0d0c0c0c0c0b0c0b0b0c0a090a080800010201020100090c0c;
    encBuf[3157] = 256'h0d0c0b0c0a0a09080003040404030202010108090a090a080003050404030304;
    encBuf[3158] = 256'h0304030404030503040202020108080809090801030703050303040201000008;
    encBuf[3159] = 256'h080a0a090a0a0a08080002030404030301080b0f0d0b0d0a0b0a0a0800000100;
    encBuf[3160] = 256'h08090d0c0c0d0b0b0b0c0a0909080808080808090b0d0d0b0d0b0c0b0b0b0a09;
    encBuf[3161] = 256'h0800020304030202000a0d0e0b0d0b0a0b09080002030404030302010109090b;
    encBuf[3162] = 256'h0c0b0c0a0a08000307030603030303020008090b0c0b0b090802040504040303;
    encBuf[3163] = 256'h0402020108080a0b0d0b0b0b0a08010304050303030200090a0d0b0c0c0b0a0a;
    encBuf[3164] = 256'h09080102040305020201080a0c0d0c0b0c0a090800010203030402010100080a;
    encBuf[3165] = 256'h0a0c0b0b0d0a0a0a0900010404040402020100090b0e0c0b0b0b0a0800030603;
    encBuf[3166] = 256'h050302030100080b0a0c0b0a0a090900090809090a0909080306040402020009;
    encBuf[3167] = 256'h0c0c0d0b0c0a0b09090908080001020504040302020208080103070707040403;
    encBuf[3168] = 256'h030201080a0d0c0c0a0a0801040504040203010008090b0b0c0a0a0900010203;
    encBuf[3169] = 256'h04030403030303030201080a0c0c0c0b0a0901020603040303020109090c0b0c;
    encBuf[3170] = 256'h0b0a0a0908000002020100090d0d0c0d0b0c0b0b0b0909080000010000090c0c;
    encBuf[3171] = 256'h0d0c0c0b0b0c0b0a0a090908000001010008090b0e0c0b0d0b0c0a0a09090101;
    encBuf[3172] = 256'h03050402030100080a0c0c0a0b0a080104050403050304030203020108080a0b;
    encBuf[3173] = 256'h0c0b09080306050503040302020100090a0a0b0b0b0900020405040403020302;
    encBuf[3174] = 256'h00000a0b0d0b0c0a0a0a08080102030304020101090b0f0c0c0c0b0b0b0a0a08;
    encBuf[3175] = 256'h0002020202000a0d0d0c0c0b0c0a0a09090800080000000809090c0b0d0c0c0a;
    encBuf[3176] = 256'h0b0b0a09080001020303030100080c0c0c0c0b0a0a0801030603050302030101;
    encBuf[3177] = 256'h0808090a080002040504030404020303030303020109090b0c0b0a0004070404;
    encBuf[3178] = 256'h0403030200080a0b0d0b0c0a090900010203040202010008090c0d0b0d0c0a0b;
    encBuf[3179] = 256'h0b0b090900020403040201000a0c0c0d0b0c0a0a09080001020303030300000a;
    encBuf[3180] = 256'h0c0c0c0d0a0b0a0900010205030403010200090a0b0c0b090a08010305050403;
    encBuf[3181] = 256'h040303020101090b0c0b0d09090801030305040201010009090a0b0b0c0a0909;
    encBuf[3182] = 256'h00010103030205030304040404020301090c0d0c0a0105070505030403010109;
    encBuf[3183] = 256'h0c0c0c0c0a0900010405030403020000090b0c0b0b0a09080103030504020302;
    encBuf[3184] = 256'h0202010008090b0c0c0b0a090802050404040202010008090b0c0b0b0a0a0908;
    encBuf[3185] = 256'h00020403030301090b0f0d0c0c0b0b0b0a0900000202020208090d0d0c0c0b0b;
    encBuf[3186] = 256'h0b0b0a090908000801000808090b0d0c0c0b0c0c0a0b0a090801020403040302;
    encBuf[3187] = 256'h00080b0e0c0b0a0a080104050403040302030102010100010000080808010307;
    encBuf[3188] = 256'h060405040304020201080a0b0d0b0b090902040405030303020108090c0b0b0c;
    encBuf[3189] = 256'h0a0a0a08010103040403030302000a0d0d0c0b0c0b0b09080002030502010109;
    encBuf[3190] = 256'h0a0d0c0c0b0b0b0a0a0808000201020101090b0d0d0c0b0c0b0b0b0909000203;
    encBuf[3191] = 256'h0403030100090c0e0b0c0b0a0a080102040305030202000008090b0a0b0a0900;
    encBuf[3192] = 256'h030605040404030302020100080a0a0b0a090003070305030304020101010808;
    encBuf[3193] = 256'h080a0a0a0b0b0a08020505040403030201090a0d0c0c0b0c0a09090800010303;
    encBuf[3194] = 256'h030301080a0e0c0d0b0c0a0a090808000101010008080a0b0c0b0c0c0b0b0c0a;
    encBuf[3195] = 256'h0a09080001010200080c0d0c0c0a0a0900000204030202010809000908010908;
    encBuf[3196] = 256'h0809020604050403030400080b0e0b0b0b090104050404030202010008090b0c;
    encBuf[3197] = 256'h0b0d0b0b09080206040503040201010808000104060503030301080b0f0b0c0b;
    encBuf[3198] = 256'h09000306040403030200080b0b0d0b0b09080102040403040203010101080809;
    encBuf[3199] = 256'h0b0c0b0b0a0800030704030403020108090a0c0b0c0a09090801020303040101;
    encBuf[3200] = 256'h080a0d0d0c0b0c0b0c0a0908080102010201080a0c0e0c0b0c0b0b0a0a090808;
    encBuf[3201] = 256'h01010001080a0c0c0d0b0c0b0a0b0a0a09000000030303030300090c0d0d0c0b;
    encBuf[3202] = 256'h0b0b09010307040403030303020008090a0a0909000305060404030403040202;
    encBuf[3203] = 256'h010100080a0a0a0909000205050404030302020008090a0b0b0b090801040304;
    encBuf[3204] = 256'h03020201090a0b0c0c0b0b0b0c0b0b0b0b0b0a0b0b090c0c0d0e0c0c0b0c0b0c;
    encBuf[3205] = 256'h0a0909080808080a0b0c0d0b0c0b0b0b0a0a0909090a0b0c0b0c0c0a0b0a0a0a;
    encBuf[3206] = 256'h0a0a090a0909090001010108090c0d0c0c0b0b09080206040503030502020201;
    encBuf[3207] = 256'h0100010102020204040304040303040403030303020101000008090800020405;
    encBuf[3208] = 256'h0403030402030201000909090a0b0a0c0b0b0a0a080008000108080c0f0d0c0c;
    encBuf[3209] = 256'h0c0a0b0b0b0b0b0a0b09090a0a0b0e0c0d0c0c0c0b0a0a0a0001020304030108;
    encBuf[3210] = 256'h0b0f0b0d0b0b0a08080103040303020008080c0b0c0c0b0a0908010204040304;
    encBuf[3211] = 256'h030100090a0b0b0c090909000303060402030403040402020008090c0d0b0c0b;
    encBuf[3212] = 256'h0a08030605040402020100090a0c0a080106060404030202000a0b0f0b0b0909;
    encBuf[3213] = 256'h020406030403020108090b0c0c0a0908000304030502020200000808090a0b0a;
    encBuf[3214] = 256'h0a0a0801040405040304020000090a0c0b0c0a09090002020403020201080a0c;
    encBuf[3215] = 256'h0d0b0d0b0b0b0c0a0908080102020101080b0e0d0c0b0c0b0a0a090800000008;
    encBuf[3216] = 256'h090a0c0c0c0b0c0a0a0a0a08090808080909090a08090808090a0c0d0c0c0b0a;
    encBuf[3217] = 256'h090104060404030302020009090a0a0801050403040301020101030704060304;
    encBuf[3218] = 256'h03030100090c0c0b0b0a00020604040303030100080b0b0c0b0a090800010303;
    encBuf[3219] = 256'h06030303020200090b0e0d0b0c0b0a080001030503030200080c0c0d0b0b0b0b;
    encBuf[3220] = 256'h090808010202010008090b0d0c0b0d0b0b0c0a0b0b0a08080102020200090c0d;
    encBuf[3221] = 256'h0d0c0b0c0a090801010202020200090a0b0c0b09000101010101000102030605;
    encBuf[3222] = 256'h0405030303020101000800010105040503040202030202040303030203000a0c;
    encBuf[3223] = 256'h0e0b0a09020505040303030208090c0c0b0b0b09080001020403030302010000;
    encBuf[3224] = 256'h090b0f0e0c0c0b0b0a0a0800030504030201080a0d0c0c0c0a0b0a0900000202;
    encBuf[3225] = 256'h0303020100090b0d0b0c0b0b0c0b0a0b0a080002040504030101090b0d0c0b0b;
    encBuf[3226] = 256'h0a0a000103050302010009090a0b0c0b0b090000030404030603030401010009;
    encBuf[3227] = 256'h0808080000000101030606050604050403030201090b0e0c0b0b090802060404;
    encBuf[3228] = 256'h0402020000090b0c0b0b090901020503050202020008080a0b0b0b0a0a090103;
    encBuf[3229] = 256'h0505030403020101090a0c0c0b0c0909080002030403020200090b0c0d0c0b0b;
    encBuf[3230] = 256'h0c0a0a0a0900000102010200090d0c0d0b0c0b0b0a0a090808000008080a0c0b;
    encBuf[3231] = 256'h0d0b0b0b0b0b0a0b0b0c0c0b0a0a0a08000204030301000a0d0d0c0b0c0a0900;
    encBuf[3232] = 256'h030504050303040202010100080809080801050505040403030303020008090b;
    encBuf[3233] = 256'h0b0a09010504060304030203010009090a0b0a0a080003060403040302020008;
    encBuf[3234] = 256'h0a0b0d0c0a0b0a0909000102020201000a0d0d0d0c0b0c0b0b0a0a0908090808;
    encBuf[3235] = 256'h0a0b0d0d0c0b0c0b0b0a0a0a080808080a0b0d0c0d0b0b0c0a0a0a0909000801;
    encBuf[3236] = 256'h080100000100080a0b0d0c0c0a0b0a0a00010306030403030303030304020403;
    encBuf[3237] = 256'h0304030304030405030403040304020302030201020000080900010406050404;
    encBuf[3238] = 256'h030302020100090b0b0b0d0a0a0a08000204040403030201080b0f0c0b0c0b0b;
    encBuf[3239] = 256'h0a090800010303030200080a0c0c0d0d0b0c0b0b0c0a0909000101020201090a;
    encBuf[3240] = 256'h0d0d0b0c0b0c0a0b090909000102020302020008090c0c0c0c0c0b0b0c090a00;
    encBuf[3241] = 256'h010205030403020108090c0c0b0b0b080104050404020302010808080a090908;
    encBuf[3242] = 256'h010204060403050203010008090800040705040404020200080b0c0c0b0b0901;
    encBuf[3243] = 256'h0405050304020100080a0b0c0a0a0801020404040202000000090a0a090a0908;
    encBuf[3244] = 256'h0101030504030402030108090c0c0d0b0a0a080002040304020208090a0d0b0c;
    encBuf[3245] = 256'h0b0b0a0a0a090909090908080809090d0c0e0b0d0b0b0c090a0900000800080b;
    encBuf[3246] = 256'h0c0d0c0b0b0a0a0900000800090c0c0c0b0b0a08010204030302080a0d0c0c0a;
    encBuf[3247] = 256'h0a08000204050304030303040201020100080808090800040405050305030404;
    encBuf[3248] = 256'h030304030201000a0b0e0b0b0908020605040303030200080b0c0c0b0b0a0901;
    encBuf[3249] = 256'h020404040203010108090c0c0b0c0b0b090900020305030201080a0c0d0c0b0b;
    encBuf[3250] = 256'h0b0b090908080101010000090b0d0c0d0b0c0b0b0c0b0a0a0909000101020108;
    encBuf[3251] = 256'h0a0c0d0c0b0b0c0a09090801000201010100080808000302040302080a0c0a09;
    encBuf[3252] = 256'h0307070603030403020101080809080900020405040403030303030202020101;
    encBuf[3253] = 256'h00080908090103060505030403020100090b0b0d0a0a0a080001030302030200;
    encBuf[3254] = 256'h080a0b0e0b0d0c0b0d0b0b0b0a090808010009090e0d0b0d0b0b0a0b0a090a09;
    encBuf[3255] = 256'h0a0a0b0d0b0c0b0c0a0b0b0c0b0b0b0a0c0a0b0a0a0a0a08090801020303090d;
    encBuf[3256] = 256'h0e0e0c0b0b0a080104050404020200080a0b0d0b0a0a08030406030403020301;
    encBuf[3257] = 256'h08080a0b0c0908000305040403030303040304050403030201090b0e0c0c0909;
    encBuf[3258] = 256'h010504040403020100090b0d0b0a0a08010404030402020108090a0a0b0a0908;
    encBuf[3259] = 256'h0001030404040203030101080a0c0c0b0b0b0908020304040202000a0b0d0b0c;
    encBuf[3260] = 256'h0a0a0a0b0a0b0c0b0c0b0c09090908090b0d0c0d0b0b0c0a0b0a0908090a0a0c;
    encBuf[3261] = 256'h0c0b0c0c0a0b090a0908090a0b0e0c0b0b0b0a0a00020404030201090a0e0c0c;
    encBuf[3262] = 256'h0a0b090802040404030402020100080809090809000104050405040304020301;
    encBuf[3263] = 256'h010009090a090900030604040403020301000808090909080102030504030202;
    encBuf[3264] = 256'h0208080a0b0d0a0b090800010101090a0e0c0c0c0b0b0c0a0a0a0b0a0c0b0b0b;
    encBuf[3265] = 256'h0d0b0c0b0c0c0b0c0b0c0b0b0a0a090908090a0b0d0c0d0b0c0b0b0a09090808;
    encBuf[3266] = 256'h000808080a0b0b0c0b0c0a0a0a09090900080808000103050504030404030304;
    encBuf[3267] = 256'h0303030304030404030404030402030203020203020304040303050204020303;
    encBuf[3268] = 256'h0403040402030301010109080909080203050403030300090a0d0c0b0b0c090a;
    encBuf[3269] = 256'h0908090a0b0e0c0b0c0c0a0a0b0b0b0d0b0d0b0c0c0b0a0b0a0a090909080a0b;
    encBuf[3270] = 256'h0d0e0b0d0a0b0a0a080000010000090c0d0c0b0c0b0a09000102050304020108;
    encBuf[3271] = 256'h090b0e0b0b0b0a0801040404040303020100080a0a0a09080204050404030303;
    encBuf[3272] = 256'h030202020108090b0c0b0a080207050404040303020101080908080203070402;
    encBuf[3273] = 256'h0201080b0c0c0a000207040503030200000b0c0b0d0a08080204040304020101;
    encBuf[3274] = 256'h09090a0b0b0b09080002040403050203020100090b0c0c0c0a0a080001040304;
    encBuf[3275] = 256'h030201000a0b0e0b0b0b0b0a0a0908090a090b0b0b0b0c0b0c0c0c0c0d0b0c0b;
    encBuf[3276] = 256'h0b0a0a0a0808080008090b0d0c0c0b0b0c0a0a0b0b0b0d0c0a0b090800030504;
    encBuf[3277] = 256'h020200090c0d0c0b0b0a09000305040304020200000809090900010203050402;
    encBuf[3278] = 256'h0403040304030403030301010809090808010504050402030302010008080008;
    encBuf[3279] = 256'h00010008080a0a0c0a090103070303040100090c0c0c0c0a0b0b0b0b0b0b0b0b;
    encBuf[3280] = 256'h0b0a0c0a0b0c0c0b0f0b0d0b0c0b0b0b0b0b0b090a0908090a0a0d0c0d0c0b0d;
    encBuf[3281] = 256'h0a0b0a0a090808000000000008090909090a0b0d0b0c0b0a0908020505040403;
    encBuf[3282] = 256'h0303020100080909080901040505040305030304030202020001000801010104;
    encBuf[3283] = 256'h04040305030402030302020201000008090b0a0c0b0b0909000202050201000a;
    encBuf[3284] = 256'h0f0d0c0c0c0b0b0c0a0a090909080909090b0c0c0c0c0b0c0c0b0c0a0b0a0a08;
    encBuf[3285] = 256'h080101010101080c0d0d0d0b0b0c0a0a09000101030202020008090b0d0b0c0b;
    encBuf[3286] = 256'h0b0a080203060404030302010108080909080002040504040303030303040304;
    encBuf[3287] = 256'h0305020303020201000101010305030603050403030402030101010001030504;
    encBuf[3288] = 256'h050403020200090b0d0a0a080207040403030300080b0d0b0c0a080003040403;
    encBuf[3289] = 256'h03020100090a0c0a0a0a09080801030306030403030100090c0c0d0b0a0a0900;
    encBuf[3290] = 256'h020403030302080b0c0d0c0a0b0a0a0a0a0a0a0c0a0b0a090a08080a0b0e0e0b;
    encBuf[3291] = 256'h0d0c0b0a0b0a080800000108080c0c0c0b0c0b0b0a090a090a0b0b0d0b0a0a09;
    encBuf[3292] = 256'h010205030202080b0d0d0c0b0909000305040402030102010001020102030302;
    encBuf[3293] = 256'h020101040605050405030302030008090b0b0c09000205050403020302010808;
    encBuf[3294] = 256'h0a090a090808010102040303040302020200090b0e0b0d0a0a0a09000800080a;
    encBuf[3295] = 256'h0c0d0c0c0c0a0b0a0a0a0a0b0b0c0d0b0d0b0c0b0a0b0a090a09090b0b0e0c0b;
    encBuf[3296] = 256'h0d0b0b0b0b0b0b0a090908080808090a0a0b0d0c0c0b0c0b0a09080204050404;
    encBuf[3297] = 256'h0202010808090b0a080801050405040204020202020100010102020205030403;
    encBuf[3298] = 256'h04030302020201000101010404040403020200080a0b0c0b0a0b0a080909080a;
    encBuf[3299] = 256'h0b0b0f0b0c0c0b0d0c0c0b0c0b0b0b0a09090808090a0d0d0c0c0b0b0a0a0800;
    encBuf[3300] = 256'h000008090b0c0c0c0a0b0b0a0a0a0b0b0c0909080302030400080b0e0c0b0b09;
    encBuf[3301] = 256'h0103070303030200000908000307050403030202020101010202040403040303;
    encBuf[3302] = 256'h0503040403020302010102030404040404020101000009080002030604030303;
    encBuf[3303] = 256'h03020203060306030302000a0d0c0d0a09080306040403030100090c0c0b0c09;
    encBuf[3304] = 256'h09000203050303020100090a0b0c0b0a0a090901020405030304020108090c0c;
    encBuf[3305] = 256'h0b0c0b09080003030503020108090b0d0b0c0a0b0909090809090a0b0c0a0b0a;
    encBuf[3306] = 256'h0a090b0a0e0c0c0c0c0b0b0c090a09080800080a0a0b0d0b0c0b0a0b0b0b0c0c;
    encBuf[3307] = 256'h0b0b0c0a0900020503030301080b0f0c0b0c0a0a000105040304030301010008;
    encBuf[3308] = 256'h080a090908000102050603060304030303020108090b0b0c0908020505040403;
    encBuf[3309] = 256'h0302010108090a0a0a0a09090102040404030303010208090a0c0c0b0b0c0b0b;
    encBuf[3310] = 256'h0a0a0a0800000101090a0e0e0c0c0b0c0b0c0a0a0a090a0a0a0a0b0c0b0b0c0b;
    encBuf[3311] = 256'h0b0c0c0c0b0d0b0b0c0a0a0908080100010009090c0c0c0b0c0a0b0908080103;
    encBuf[3312] = 256'h0303040302020001010800000802030406040304040304040303040202020201;
    encBuf[3313] = 256'h010203040504030403030202020008090a0b0b0b0a080103070404020200090d;
    encBuf[3314] = 256'h0c0d0b0c0b0c0a0909080808000809090b0d0c0b0d0c0b0b0b0b0b0909080900;
    encBuf[3315] = 256'h000800080a0a0d0c0c0d0c0b0c0a0a090102050403020200090b0d0b0b0a0901;
    encBuf[3316] = 256'h030603050203010108000908000002030404050305020302010008090a090002;
    encBuf[3317] = 256'h0704040304010100080a0a09090103060304030301010809080908000008080a;
    encBuf[3318] = 256'h0a090107060503040301000a0b0d0a0a01030703040200090c0c0b0a09010406;
    encBuf[3319] = 256'h03040201090a0c0c0b0a0900020405020301010809090a0a0a08080800010203;
    encBuf[3320] = 256'h0504040303030200080b0d0b0b0a000104050304020000090b0c0b0b0a090808;
    encBuf[3321] = 256'h010100000a0b0c0d0b0c0b0b0c0b0b0b0d0b0b0d0b0c0a0a0a0b0a090b0b0c0d;
    encBuf[3322] = 256'h0c0c0b0c0a0b0b0a0a0a09090a0a0a0b0a0a090808090b0f0d0c0c0b0b090004;
    encBuf[3323] = 256'h06040304020000080a0a0a090002050503030202020100020304040503030201;
    encBuf[3324] = 256'h0108080801020504040402020200000000080000010102020101080008000102;
    encBuf[3325] = 256'h020401090b0f0f0b0c0b0b0b0a0a0a0a080a0b0b0e0c0b0d0b0d0c0c0b0b0b0b;
    encBuf[3326] = 256'h0a0a08090808090a0c0c0c0c0c0b0b0d0b0a0b0909000002020202080b0e0d0c;
    encBuf[3327] = 256'h0b0a0a08000102020301010008080003060403030108090b0d0a090803060504;
    encBuf[3328] = 256'h0403030302020201010008000808080000020704050304030200090a0d0b0c0a;
    encBuf[3329] = 256'h08000104020301080b0d0d0b0b0b0a0800000101080b0c0d0d0a0c0a090a0908;
    encBuf[3330] = 256'h0908080809090c0c0b0d0c0a0b0a0a09090808080809080008010208090a0f0c;
    encBuf[3331] = 256'h0b0c090801050403030302010100020302040201020303050604050404030302;
    encBuf[3332] = 256'h0108080808080001020503040302020306050304020108090a0b0b0b0a010407;
    encBuf[3333] = 256'h03030302000009090a0b0a0a08040405030304030200090c0d0a0a0902030405;
    encBuf[3334] = 256'h020201090c0c0c0a0003050504020301000a0c0d0b0a09000204040304030101;
    encBuf[3335] = 256'h08090a09000001010302030402010002030704030200090a0b0b0a0a09020605;
    encBuf[3336] = 256'h04020109090b0b0a0b090b09080101000d0e0b0c0a09090a0b0d0a0a0a0b0c0d;
    encBuf[3337] = 256'h0b0b0a0b0a0c0c0b0b0a09090b0d0c0a0a0a0b0b0f0b0a0a0a0a090800040504;
    encBuf[3338] = 256'h0201080a0e0b0d0b0b0a08020505040202010009090a0c0a0900010303040303;
    encBuf[3339] = 256'h040303020302010100080a0b0c0901060505030402030101090b0c0b0a090002;
    encBuf[3340] = 256'h03050403040101080a0a0b0b0c0b0c0b0909010103020201000a0f0d0c0b0b0b;
    encBuf[3341] = 256'h0a0a0b0c0b0b0b0b0c0c0a0a0908080b0d0c0d0b0a0c0a0a0b0a080908090b0b;
    encBuf[3342] = 256'h0c0b09080808090a0b0d0e0c0c0b0a09080102040304030301000a0d0b0a0b08;
    encBuf[3343] = 256'h000204050403050203020201010009090a0a0808030704050304030301000009;
    encBuf[3344] = 256'h09080a09090800020305040202040204030302000a0c0e0c0c0b0a0900020304;
    encBuf[3345] = 256'h03020108090a0d0c0c0b0a0a08000000000008090c0e0c0c0a0a090808010104;
    encBuf[3346] = 256'h03050101090a0d0b0b0c0b0b080003060303030202020200090a0b0a090a0a0c;
    encBuf[3347] = 256'h09010507040402020202020201080809080001020202030303010b0d0b080706;
    encBuf[3348] = 256'h040303030201080a0d0c0c0b090900000102030604030402020100080a0e0d0b;
    encBuf[3349] = 256'h0b09080304050304020108090a0b0a080304050403020100090a0b0c09000204;
    encBuf[3350] = 256'h04040403030402010108090a0c0b0b0a0901050505030402020108090c0b0b0c;
    encBuf[3351] = 256'h0908000202020302010009090a0b0d0b0d0a0a090908080a09090a0a0e0d0c0b;
    encBuf[3352] = 256'h0c0a0a0a090a0909090a0c0d0d0b0b0b0a0b0a0b0a090808080c0c0d0b0b0b0b;
    encBuf[3353] = 256'h0c0a0908010202080b0d0d0c0a0a0900030505020201090a0c0b0a0a08020605;
    encBuf[3354] = 256'h0403030302010008000808080101020403030404040503040202010008080801;
    encBuf[3355] = 256'h030404030201080a0c0b0b080004040404030201090d0d0c0b0b0b0a0a0a0909;
    encBuf[3356] = 256'h000204040201080b0e0d0c0c0b0b0b0b0909000002010100090c0c0b0a0b0a0a;
    encBuf[3357] = 256'h0b0d0b0b0b0a0a0a0a0c0b0b0a080205050404020301000a0b0e0c0b0a0a0801;
    encBuf[3358] = 256'h030404040402030202000008090b0b0c0a00030705040302030108080a0a0b0b;
    encBuf[3359] = 256'h0a0900010404040402030200000009090a0c0b0a090801030403020201010103;
    encBuf[3360] = 256'h010a0f0f0e0b0b0c0909080001020304020300080b0c0d0b0b0c0b0b0c0b0c0b;
    encBuf[3361] = 256'h0a0803050504020201000a0b0e0c0b0b0b090801020403050303030200080a0b;
    encBuf[3362] = 256'h0c0c0b0b0a0900040504040203010009090b0c0b0a0900030604040304010100;
    encBuf[3363] = 256'h0a0b0c0b0b0b0900020406030403020108080a0b0c0b0b0b0a09020406040403;
    encBuf[3364] = 256'h02000009090a090a0909080001030304020100010204070403030301090b0d0b;
    encBuf[3365] = 256'h0a090103040502020303030303020202010108090b0d0b090800030604050303;
    encBuf[3366] = 256'h0201090b0d0c0b0a0a000203070402030201090b0f0b0d0b0c0a0a0808010304;
    encBuf[3367] = 256'h04020100080a0c0d0b0d0b0a0a09080801010203030201000a0b0e0c0d0c0b0c;
    encBuf[3368] = 256'h0b0a09000203040303020101090a0d0c0c0c0a0a080103050303010108090a0a;
    encBuf[3369] = 256'h0a09000204050302020008090908000307040303020000000103040202010102;
    encBuf[3370] = 256'h00000b0e0c0b0a000204050304020200090c0c0c0b0b0a0a080001010101080b;
    encBuf[3371] = 256'h0d0d0d0c0c0a0b09090908090a09090808090b0e0d0c0b0b0a0a0a0a09090800;
    encBuf[3372] = 256'h01020201090d0e0c0c0a09000808080b0a080106040201080809000001080a0a;
    encBuf[3373] = 256'h00050704020201080a090a08020406040303020102020101080c0c0c09000206;
    encBuf[3374] = 256'h03040302010108090a0a0908020200090c0d0b090900030305030301080b0e0c;
    encBuf[3375] = 256'h0b0c0a0a0b090a0a0a0c0b0c0b0a090909080a0a01040405010a0e0e0c0b0b0b;
    encBuf[3376] = 256'h0800020404030201080a0c0c0a0b090800000101010102040604030208090b0b;
    encBuf[3377] = 256'h0a0908090b0c0a0007050503030300080a0d0b0b0a0802030503030303020301;
    encBuf[3378] = 256'h0202030202080e0d0c0c0a0a080204050503030201080a0a0a09000203040201;
    encBuf[3379] = 256'h00090a0b0a00020605040404030101080a0a0a09080800080003050404040202;
    encBuf[3380] = 256'h02020200080808080000000305050302090d0c0b08030704030101000008080a;
    encBuf[3381] = 256'h0a0b0d0a0a09080000020303070302040100090c0e0c0b0a090901010101080a;
    encBuf[3382] = 256'h0b0c0b0c0a0a09090a0a0a09090008080b0f0f0b0c0b0a090909080a0b0b0b08;
    encBuf[3383] = 256'h0105040201080b0d0c0b0b0b0b0a08010201080a0a080507050203010009090a;
    encBuf[3384] = 256'h0a0b0b090003050403030403040302000809080103060403030201080c0c0d0b;
    encBuf[3385] = 256'h0a000104050303010009090b0b080801080d0e0d0c0a0908020402020109090b;
    encBuf[3386] = 256'h0c0a0b0b0b0c0c0b0b0d0b0b0a0900020202080b0f0e0b0b0a0a090900010102;
    encBuf[3387] = 256'h01090a0e0c0b0c0a0a0909090908020204040201000b0d0c0b0c0a0a09000103;
    encBuf[3388] = 256'h050405040203010009090b0b0a09000205050403020108090908000304030203;
    encBuf[3389] = 256'h040404030200090900020504030301080a0b0d0b0c0a09010505040402020008;
    encBuf[3390] = 256'h0b0d0b0b0a090900000801020304030101090a0a0c0d0d0c0b0b0a0003040302;
    encBuf[3391] = 256'h010b0d0c0c0a0b0a08000204050201000b0d0b0c0a090000010100080a090900;
    encBuf[3392] = 256'h0306030100090b0a080800090c0c0c0a0a0802070604040303020008090b0b0c;
    encBuf[3393] = 256'h0b0b0a080204040404030403030301010809090a0b0a09000406040304030304;
    encBuf[3394] = 256'h020100080a0a0a0a0800040505040402010108090a0909010104030402020101;
    encBuf[3395] = 256'h000002030403040201000909090b00020506030401010a0b0c0b090103070302;
    encBuf[3396] = 256'h01090c0d0c0b0a090808000800090801020303080d0e0d0d0b0b0b0b0a080000;
    encBuf[3397] = 256'h00000809090a0c0c0d0c0b0a0a000100080a0e0c0c0b0a0a0800010202030101;
    encBuf[3398] = 256'h090c0c0c0d0a0a0a0800010202020204020201090b0e0a0a0808010102030404;
    encBuf[3399] = 256'h02020108000901020604030301080a0d0a09000202030403040201090d0d0c0a;
    encBuf[3400] = 256'h09080101010108090c0d0c0a09000002080c0c0d0b0c0a0b0a0a0a0908090909;
    encBuf[3401] = 256'h0908090c0e0e0d0b0b0a080008080b0d0b0c0a09090a08080003040302080c0d;
    encBuf[3402] = 256'h0d0b0c0b0a09000204040200080a0b0c0c0b0a09010405040101000909090809;
    encBuf[3403] = 256'h090900050403040009090a080203070303030208090b0c090103060301000809;
    encBuf[3404] = 256'h080001020705040502030008090c0c0a0a090802030304030303030403020200;
    encBuf[3405] = 256'h090b0e0c0c0909000304030301000908080203050302080a0e0c0c0a0b0a0900;
    encBuf[3406] = 256'h0306040304010100090a0c0c0c0b0a0909000202040403030302080b0e0c0c0b;
    encBuf[3407] = 256'h0a090002040303010100080000080a0b0b090105040200090c0b080106040403;
    encBuf[3408] = 256'h03040201000a0b0c0c0a090004050404030202020100010000080a0908010503;
    encBuf[3409] = 256'h03020101050504040402020201020100090b0d0a09080205050403030100080a;
    encBuf[3410] = 256'h09090800010102020201090a0a0a030703040108090b0e0a0c0c0a0b0a090809;
    encBuf[3411] = 256'h080809080a0b0d0d0d0b0c0b0a0909000108080b0f0b0d0b0b0a0a0908080000;
    encBuf[3412] = 256'h090b0d0e0b0d0b0a0a090002020402020008090a0d0b0d0b0a0a00000100090a;
    encBuf[3413] = 256'h090a000103030305040403020200080a0c0b0a080307040201080a0b0b080205;
    encBuf[3414] = 256'h0503030302000c0f0c0b0b0a0004040403030100080a0b0d0b0c0b0c0a090801;
    encBuf[3415] = 256'h0103030302080a0f0d0c0b0b0a00000203010108090a0c0c0b0c0a0b0c0b0b0a;
    encBuf[3416] = 256'h0a01020303000a0d0e0c0b0c0a0a0001040201080b0d0a080001020202000008;
    encBuf[3417] = 256'h090b0e0c0b0a090203020201090a000104060202020808000802040305030203;
    encBuf[3418] = 256'h020101010a0e0d0c0b09000407030503020101090c0b0d0a0800030502020202;
    encBuf[3419] = 256'h010201010109090b0d0a0909000100030404050503030302020201080a0f0c0b;
    encBuf[3420] = 256'h0a090103060402030302000a0b0d0c0b0b0a0901030604030302010009090b0d;
    encBuf[3421] = 256'h0b0c0b0909080100000001020405030200090b0d0c0b0b0b0a09000305030502;
    encBuf[3422] = 256'h010108080a0a0b0e0b0d0b0b0b0a0003060504040202020008090b0c0b0c0908;
    encBuf[3423] = 256'h0103050304020101010101010100080808090102050604050304020201000001;
    encBuf[3424] = 256'h0000000009090a08010105050405040203010108090b0b0b0a09010307030303;
    encBuf[3425] = 256'h0101000108090c0e0b0d0a0b0a0a0a0908010405030301000a0d0d0c0c0c0a0a;
    encBuf[3426] = 256'h0908010202030301080b0e0c0b0c0b0b0a0b0a0a0001040403020108090b0c0c;
    encBuf[3427] = 256'h0b0c0b0b0a090102030402020100080b0e0c0b0b0a080205040304020200080a;
    encBuf[3428] = 256'h0a0900040403010109090a09080003050603030100090b0a0b0b0a0a01040704;
    encBuf[3429] = 256'h030302000809090b0e0d0b0a0a00010200080b0d0c0b0b0a0900020302010a0f;
    encBuf[3430] = 256'h0d0c0c0b0b0a09000205020200090b0d0c0c0a0b0a0a09090808080103050402;
    encBuf[3431] = 256'h030108090c0d0c0c0b0a0a0001040304020200080a0b0c0b0a08080002020304;
    encBuf[3432] = 256'h0201010908020406040100090d0b0a0a0908090809080205050403030101090a;
    encBuf[3433] = 256'h0b0c0b0a0a08020406040201080d0b0c0a090204040403020100090b0e0b0b0b;
    encBuf[3434] = 256'h00020505030402010008090a0b0a0a0a0909000203050404030503030200090b;
    encBuf[3435] = 256'h0d0b0a0908020403030403020101000008090a0c0b0c0a090001020305030202;
    encBuf[3436] = 256'h02030406040301080c0d0d0a0a0901010302010009090908030504030301080b;
    encBuf[3437] = 256'h0f0c0b0a090004050403020202010101090a0d0d0b0a0a020406040402030101;
    encBuf[3438] = 256'h0108090a0b0d0a0a0803050504030303020100080b0b0c0a0908020504030303;
    encBuf[3439] = 256'h030202010101080a0b0c09090802030205040306020200090b0b0c0b0a0b0c0b;
    encBuf[3440] = 256'h0c0b080001030302000a0f0d0b0d0b0b0c0a090a080908090a0c0a0b0a000101;
    encBuf[3441] = 256'h000d0e0d0c0c0b0a0b0909010204030400080b0c0d0a0b0a0a0a000003040302;
    encBuf[3442] = 256'h02000808080a0c0c0d0c0b0a090001040305030201010009090a0c0b0c0b0900;
    encBuf[3443] = 256'h02030403020304030201090d0c0b0a0b0b0c0c0c0a0a08010404030401000a0b;
    encBuf[3444] = 256'h0d0c0b0b0b0b0a0801010201090a0b0c0d0b0e0b0c0a0a08080800080009090a;
    encBuf[3445] = 256'h0b0b0c090909090b0a090a0a0d0f0b0b0a0801000a0c0d0a080000000c0b0b09;
    encBuf[3446] = 256'h0207030303010203010202090a0c0f0c0c0b0b09090003020405030403010808;
    encBuf[3447] = 256'h0b090909090a0e0b0b0a00040405030302030200080b0f0b0d0a080803040302;
    encBuf[3448] = 256'h0109090809010403060403030301090b0e0a0a09080809090808050604050302;
    encBuf[3449] = 256'h030100090b0d0b0c0a090900030504050303010108090a0c0c0c0a0a08000304;
    encBuf[3450] = 256'h0402030203020200080a0d0b0c0b0a0a08000203040403030202000a0a0c0b0b;
    encBuf[3451] = 256'h09000104030504020201000809090b09080101080c0f0d090003070403020102;
    encBuf[3452] = 256'h010100080a0b0b0902040403050304040303020201010108080a0a0801050402;
    encBuf[3453] = 256'h050403070303040201010808080a090800020504030303020102080100090009;
    encBuf[3454] = 256'h0a0b0a0a05060405040204030201000a0d0c0c0b0a0908000002020303030101;
    encBuf[3455] = 256'h090b0d0e0c0c0b0a0a0908000204040302010a0d0c0d0a0b0a0a0a0a09080102;
    encBuf[3456] = 256'h0101090a0c0c0b0d0a0b0908080000090a0d0b0b0c0a0a08010302000d0e0c0c;
    encBuf[3457] = 256'h0b0b0a090900010303030200080809080b0e0d0c0a0a0900010303040300090c;
    encBuf[3458] = 256'h0d0b0c0a0a0b0a0b090908010304040403040301080b0d0b0c0a0b0a0b0b0c0b;
    encBuf[3459] = 256'h0b0908010405030302080b0e0c0c0b0a09000102040202010a0d0c0c0a090801;
    encBuf[3460] = 256'h030306030201080c0c0c0c0a0a0a0a000103060304010100000008090a0a0909;
    encBuf[3461] = 256'h000100090a0b0b000105050305040303030108080a0a0b0b0a01060704040201;
    encBuf[3462] = 256'h010809090a0a0909010406040302020108090a0b0b0b0a090207050404020208;
    encBuf[3463] = 256'h090b0c0b0b0a09000204050403030108090c0b0c0b0a09090101020203020402;
    encBuf[3464] = 256'h01000b0e0c0b090900010102020303080c0f0d0b0a0002040403010008080a0b;
    encBuf[3465] = 256'h0b0e0b0b0a090802030505020302010100090a0d0d0b0b0a0104040402020101;
    encBuf[3466] = 256'h0100080b0d0c0b0b0a080802050404030402020108090b0c0b0a080204040303;
    encBuf[3467] = 256'h02020100080b0b0c0901020503020304030703040402030202010008090a0b0d;
    encBuf[3468] = 256'h0a08000505040402030203020201090b0c0c0900020503040203020304020201;
    encBuf[3469] = 256'h00000809080808090a0d0b0900070403040100090b0b0c0b0b0b0b0901050305;
    encBuf[3470] = 256'h0200000a0a0b0d0c0c0d0c0b0b0b090908010001000009090c0c0c0c0c0b0b0b;
    encBuf[3471] = 256'h0b0a0909080000090a0d0d0d0b0c0a0b090a090a0a0a090908090a0b0d0b0b0b;
    encBuf[3472] = 256'h0b0b0c0c0b0b09090009090c0b0c0b0a0b0e0c0d0b0c0909000101000008090b;
    encBuf[3473] = 256'h09010206030402020108080d0d0c0c0a0a09000002020504020300080a0b0d0a;
    encBuf[3474] = 256'h0a08080003040304030101000800000808010001010d0e0c0d0a0a0801030504;
    encBuf[3475] = 256'h030402010809090a08000001000800020100000d0b0a09030707030502020301;
    encBuf[3476] = 256'h00080b0d0d0c0b0b0901040603040303020101090b0e0b0d0a09080102040304;
    encBuf[3477] = 256'h03020100000a0b0c0c0a09080002030303040304030100090b0d0c0b0c090908;
    encBuf[3478] = 256'h0203040403030201080a0b0d0b0c0b0a0c0a0a08020504040302020108080c0c;
    encBuf[3479] = 256'h0d0b0b0b090801030304040202020008080b0d0c0b0b0a090001010101030405;
    encBuf[3480] = 256'h0303030100090a0d0c0d0b0a0a0801030503040302020100080809090a0c0c0a;
    encBuf[3481] = 256'h0a080003030703060304030200090a0d0b0b0b0a080004050503040201010808;
    encBuf[3482] = 256'h09090b0b0b0c090902030704030403020108080a080908090b0b0b0a00040404;
    encBuf[3483] = 256'h0503050403030100090a0a0b0c0b0a0a0802050404030402010108080a0a0a0a;
    encBuf[3484] = 256'h090808090002060603020100090a0b0c0b0d0a0b09080102030603030300090b;
    encBuf[3485] = 256'h0d0b0c0b0d0b0c0a09080001010103020302080c0c0d0c0a0c0b0d0b0a0a0900;
    encBuf[3486] = 256'h0103030304030201090b0e0c0b0d0c0b0c0a0a0908010202040304030200090c;
    encBuf[3487] = 256'h0c0c0c0b0b0c0909080102030304030201080a0e0d0b0b0a0a00000102020101;
    encBuf[3488] = 256'h090809090a0a0b0a0a0b0a0a0d0a0b0b09010307030302000a0f0c0d0b0b0a09;
    encBuf[3489] = 256'h0802040504030201000a0c0c0a0909000102020304030201080b0d0d0b090902;
    encBuf[3490] = 256'h04040403020101000101000009090b0b0a08040604030302030203040300080c;
    encBuf[3491] = 256'h0e0b0b09080102030505060403040200090a0d0b0a0b0a090102050404020202;
    encBuf[3492] = 256'h0009090b0c0b0c0b0a0a09010505040302020108090a0b0c0d0b0b0b09010304;
    encBuf[3493] = 256'h040304020200080a0d0b0b0c0a0b0a0908030404040202020100080a0b0d0c0b;
    encBuf[3494] = 256'h0c0b0c0a09080204030302020108090b0e0d0b0b0a0908000203040203010101;
    encBuf[3495] = 256'h01000a0f0d0c0c0b0a09080203060304020100090c0b0c0b0a09080003040503;
    encBuf[3496] = 256'h030402010000090b0c0c0b0b0a09000305040403030202010000090a0d0b0c0a;
    encBuf[3497] = 256'h0001040403040503030300090c0c0c0a09090801010204030403020000080809;
    encBuf[3498] = 256'h0a0a0b0c0a0a0802040503030208090a0908000201090c0f0d0c0b0b0b0a0803;
    encBuf[3499] = 256'h07040403030108090b0d0a0a0a090a0a09090102040302000001010303000d0e;
    encBuf[3500] = 256'h0c0b0a0908000002030502030101080a0a0c0a08000204000a0f0d0b0b090a08;
    encBuf[3501] = 256'h090908020505030300080a0a09090800080a0c0c0c0b0c0a0908010305030301;
    encBuf[3502] = 256'h090f0d0c0c0a0a08010104030402030100080b0c0b0b0a0800000008090b0d0b;
    encBuf[3503] = 256'h0a0a08010504040200080a0b0b090901000103050505030301000a0c0c0b0c0c;
    encBuf[3504] = 256'h0a0a08010303040201080a0a0c0a090207040202000b0e0b0c0b090801040405;
    encBuf[3505] = 256'h030200080b0c0c0a0b0a0a09090800030404020100080a0a0a09000406040302;
    encBuf[3506] = 256'h000b0e0c0c0a0a08080102020203020301090c0d0b0b0a080204030304030202;
    encBuf[3507] = 256'h00080a0c0c0a0b0a0003050301090c0c0901050303080a0c0a08030403030303;
    encBuf[3508] = 256'h040401000a0d0a0a01040403030203040300090f0d0c0b0a0900020504030302;
    encBuf[3509] = 256'h00090b0a09000404030302000a0d0f0c0a0b08000204040203030201080b0e0c;
    encBuf[3510] = 256'h0b0b0a0808010203030404020402020100090c0b0c0b0b0b0d0b0b0a00030605;
    encBuf[3511] = 256'h03020201010009090b0d0b0a0a0908000101030305040403040100090c0b0b0a;
    encBuf[3512] = 256'h0a090a0b090805050403020009080801020202000908090809090b0d0b0b0a08;
    encBuf[3513] = 256'h040605040302000a0c0d0c0a0a09080002050403030201080a0c0a0a09090001;
    encBuf[3514] = 256'h0002030302090e0e0c0b0b0b09000102050504030301010a0b0d0c0b0a0a0801;
    encBuf[3515] = 256'h0203050304030302000a0c0e0c0b0b0b0a0a09010307050403030200000a0c0c;
    encBuf[3516] = 256'h0c0b0c0a0800020305030202020001080a0c0b0c0b0a09090000010102020403;
    encBuf[3517] = 256'h04040402010008090a0a0b0c0e0b0b0a0002040403010008000100090d0e0b0b;
    encBuf[3518] = 256'h0900030404020201030101000b0c0c0c0b0c0a0b0a0808020304040304020109;
    encBuf[3519] = 256'h0c0c0c0a090800000008010204030100090a0b0a0c0b0e0b0b0a080202020100;
    encBuf[3520] = 256'h0908080000090d0d0b0b080106040302000a0c0c0b09010304050201080a0d0c;
    encBuf[3521] = 256'h0c0a0a080104030301090c0c0a0902050503030101000000080a0c0e0c0a0a08;
    encBuf[3522] = 256'h01030203020303030301090c0c0b090002020202010206040404020201000a0b;
    encBuf[3523] = 256'h0e0b0b0902030402080a0c0a0004060403030302080d0d0c0b0b080103030502;
    encBuf[3524] = 256'h0303030201090c0c0c0a0b0a0b09090802020203020404030502000a0b0e0b0b;
    encBuf[3525] = 256'h0b0a09090900020405040302000b0f0d0c0b0a0a0801030604020200080a0c0c;
    encBuf[3526] = 256'h0c0b0c0a08000304040301010008090a0b0c0c0a0a0a09090a0b080104050402;
    encBuf[3527] = 256'h03020200080b0e0c0a0a080008090a0a0908020403040504040401080b0d0c0b;
    encBuf[3528] = 256'h0a08000001000000000102050503040200090b0b0b0b0a0a0b0c0a0b08020305;
    encBuf[3529] = 256'h04030403020201080a09090900080a0f0d0b0b0a080304050304030200080a0c;
    encBuf[3530] = 256'h0b09080101010a0d0c0a00030604030100090a0c0c0a09080002030402010101;
    encBuf[3531] = 256'h010203050303000b0f0e0b0c0a00020305020108090a09090809090801050503;
    encBuf[3532] = 256'h0201080a0b090801020300000b0f0d0d0c0b0a0a000205030402020201000008;
    encBuf[3533] = 256'h0909090a0b0d0c0b0c0b0b0a09000306040202080a0b0a0004050302080a0c0b;
    encBuf[3534] = 256'h0a0a0809080808000200080d0d0c0a09020405040302010808080808080a0e0c;
    encBuf[3535] = 256'h0b0a08010201010809000103020204040505040201090b0d0b09000306030200;
    encBuf[3536] = 256'h090a0c0b0b0a0b0b0b0a0005060404020108080801030405020108080a0b0b0d;
    encBuf[3537] = 256'h0d0b0c0b0a0808020404040303030201000800000800090b0c0d0c0c0b0a0902;
    encBuf[3538] = 256'h03050301000909080001020102020201090c0d0b0a0802030403020201020109;
    encBuf[3539] = 256'h0a0f0d0c0c0b0a0900010404030302010a0e0c0b090104050302080a0c0c0a0a;
    encBuf[3540] = 256'h0a0808010103040303020200080c0d0c0c0b0908080101030404040201090c0c;
    encBuf[3541] = 256'h0a080001000808080101010a0c0c0802060302000800020402090f0e0b0a0900;
    encBuf[3542] = 256'h01010100020403040201020102020108090a0d0e0c0d0b0a080204050200080b;
    encBuf[3543] = 256'h0a0b09010304040200090a090901030304010202030302090f0f0c0b0b0b0a09;
    encBuf[3544] = 256'h000103030503040305020201080a0909000000090d0c0c0a0a0909090a080802;
    encBuf[3545] = 256'h030404030504020301080a0a0c0d0b0b0a0105050402010808080000000a0d0d;
    encBuf[3546] = 256'h0c0a090908000000020305040304020201000809090909090b0d0d0b0c0b0909;
    encBuf[3547] = 256'h0900010204050403030200080a0c0b0c0b09090801030404030201090b0b0b08;
    encBuf[3548] = 256'h0001090d0e0b0b0b0a090b0a0901070504030101090a0a090104060301080b0e;
    encBuf[3549] = 256'h0c0a0a080808080a0a0908010205040404030302010000090a0d0e0c0c0b0a08;
    encBuf[3550] = 256'h00020304020101020202040201080c0d0c0b0b09080000010000010101020201;
    encBuf[3551] = 256'h0103050303080d0e0c0a0901040304030000090a0b0d0c0b0d0a0b0908000001;
    encBuf[3552] = 256'h020105050504040201080a0b0c0a090809090b0c0b0c09080002030503030303;
    encBuf[3553] = 256'h03030200090b0e0b09080001000a0d0d0c0a09080003030201080a0900020502;
    encBuf[3554] = 256'h000b0c0a020706040100090c0c0b0b0900010101080800010305030302010000;
    encBuf[3555] = 256'h08090c0c0e0c0b0d0a090801030304030102020304040202080b0e0c0b0c0a0a;
    encBuf[3556] = 256'h090801010101090a0b0902070604030201000a0c0d0a0a0901020202000a0a0a;
    encBuf[3557] = 256'h08010302010b0e0c0b0a0908020404050304020200090a0c0c0b0a0a09090809;
    encBuf[3558] = 256'h0909080106040502030000090b0b0c0a0a08000002020201090e0e0b0b090206;
    encBuf[3559] = 256'h040402010808080a0908090909090b0e0c0b0c0a080003060503030301080a0b;
    encBuf[3560] = 256'h0c0908000200080b0c0c0b09000000090d0b08020706030300000a0808020302;
    encBuf[3561] = 256'h090f0c0c0a09000102010108000001030302020101010405040302080c0e0c0b;
    encBuf[3562] = 256'h0b090a0909080003050403030203040305020108090a0c0b0c0c0c0b0b0a0901;
    encBuf[3563] = 256'h010303030304050303030301010008090b0d0a0a0000000a0f0f0c0a0a090103;
    encBuf[3564] = 256'h04030203020202030302080b0f0b0c0b09090900020204030302090a0c0b0800;
    encBuf[3565] = 256'h0303030200010101090d0f0c0b0b0a08080204050503040302020000090a0e0c;
    encBuf[3566] = 256'h0b0b0c0a0908080103050304010108000900080103030201080b0b0c0a0a0c0e;
    encBuf[3567] = 256'h0b0c09000205020108090909000001000101050604040201090a0b0b0a0a0b0d;
    encBuf[3568] = 256'h0d0b0a00010403030304040302000b0f0c0a09080202030100090a0901040603;
    encBuf[3569] = 256'h0301090c0d0c0a0b080001040303020203020303010a0f0c0c0b0b0a0a080801;
    encBuf[3570] = 256'h0303040403030504030401000a0d0c0b0b0c0a090800030603020200080a0a09;
    encBuf[3571] = 256'h090801020305030302080d0d0d0c0b0a0a080103040404020102010101090b0e;
    encBuf[3572] = 256'h0c0b0b0908020303040201080b0d0c0a0908020405030301080c0b0a09010303;
    encBuf[3573] = 256'h080d0d0b0b08010304020100090b0c0b090106030401080a0a09080101090b0d;
    encBuf[3574] = 256'h0900040402000b0d0c0a080002010100080909000104040301080a0e0b0b0b0b;
    encBuf[3575] = 256'h0c0a000506040301080a0d0b0a0a0800010304030200090d0b0a080204030209;
    encBuf[3576] = 256'h0d0d0a0a00030503020100080909090b0e0b0c0a08000100090b0a0803070403;
    encBuf[3577] = 256'h0000000102040208090d0b0c0a0b0c0b0a090205060304010108090a0b0b0c0c;
    encBuf[3578] = 256'h0b0c0a0a0001030303010000010205040403030200090c0c0a090800090d0f0b;
    encBuf[3579] = 256'h0c0a09010305030101080a0a0a090001020303030504030202090d0e0c0b0a09;
    encBuf[3580] = 256'h08020108090c0b09000304030108000307050303020100090a0a0c0b0d0b0c0c;
    encBuf[3581] = 256'h0b0a0900010202000809090105060404020100090d0b0b0a0002040302080a0b;
    encBuf[3582] = 256'h0a08010302080b0f0d0b0a0b0909000205040402020101000100000a0b0c0b0a;
    encBuf[3583] = 256'h0909090a0b0b080101090f0e0d0b0a0801040403020102020405040301080a0d;
    encBuf[3584] = 256'h0c0c0a09090808000908080002050503020208080908000000090b0d0d0c0a0a;
    encBuf[3585] = 256'h080204030200090a0a08020404010108080103070202080b0d0b0a0908080a0d;
    encBuf[3586] = 256'h0c0a090305050302010009090900000108080b0c0a09000a0c0f0d0b09000204;
    encBuf[3587] = 256'h0403030305020200080b09090001000c0f0c0c0a09000204040202010809090a;
    encBuf[3588] = 256'h090a0a0a0a0a0a0001040304030304030403030302080a0d0c0b0b0b0d0b0c0a;
    encBuf[3589] = 256'h00020704030200080a0b0a090908000000010205040301000b0e0c0b0a0a0800;
    encBuf[3590] = 256'h03060403030208080808010101090c0b0c0a0909090908000205030201090c0b;
    encBuf[3591] = 256'h080307050201090b0b0a02050402000a0a0c0a0b0c0c0c0b0802060504030201;
    encBuf[3592] = 256'h00090a0a0b0a090a090b0b0c090901030201090a000507060201080a0c0a0801;
    encBuf[3593] = 256'h0304020108090a09000001080c0d0c0b0a090000000800030606040304010008;
    encBuf[3594] = 256'h0b0c0c0b0908010203020000010101000b0f0e0a090002020202030305030301;
    encBuf[3595] = 256'h090b0e0b0c0a0a0900000108090900040603040201080908080809090a0c0b0a;
    encBuf[3596] = 256'h090004040302090e0c0c0909010102020303040202080b0c0d0b0c0a0a080206;
    encBuf[3597] = 256'h05040301010a0a0d0c0a0b0b090801030404020202030301010a0e0b0c090900;
    encBuf[3598] = 256'h090a0d0c0b08010604040200080b0c0b0a080102030202010001010101000a0d;
    encBuf[3599] = 256'h0c0c0a0a080008090b0c0a0a0800080909030707070302000008090a0b0d0d0b;
    encBuf[3600] = 256'h0a09000204020100000102030302080c0e0c0b0a090102050202000909090800;
    encBuf[3601] = 256'h00090b0e0b0901030403010809090809080909090206050201080c0c0b0a0802;
    encBuf[3602] = 256'h0201090c0d0a0a090908090804070404030200090a0b0c0a0c0a0c0b0a090102;
    encBuf[3603] = 256'h0603040201010001010202080b0f0d0c0a0b0908000102020303020201020303;
    encBuf[3604] = 256'h0401080b0e0b0a00020402000c0e0c0c0a0a00010403020202000000080b0c0b;
    encBuf[3605] = 256'h0b00030603020809090a08090b0c0d0b0c0a0a00010305020108090a01030605;
    encBuf[3606] = 256'h030201080b0d0d0b0a0a0a0909090003070403040101080809090a0b0c0b0d0a;
    encBuf[3607] = 256'h0b0a09090002040303030100020407040303080b0f0b0b0a0801020200090a09;
    encBuf[3608] = 256'h08010202090d0d0b0a020605030201080909080808090b0e0b0b0a0800010100;
    encBuf[3609] = 256'h000001010008080002040403020001010305030301010307050302090e0e0c0a;
    encBuf[3610] = 256'h0b0a0908000204040402020808090908090a0c0c0b0908010000080104070403;
    encBuf[3611] = 256'h010101020304010a0f0d0b0b0808010100090800010204020008080104060303;
    encBuf[3612] = 256'h00080b0c0b0b0b0d0c0b0a090103060203010001020503050201090b0f0c0a0b;
    encBuf[3613] = 256'h0900010404020201090a0b09000202010a0d0c0b090801010201010305030201;
    encBuf[3614] = 256'h0108080a0a0c0c0a0901050403030201010008090b0d0b0b0a090c0f0c0c0b09;
    encBuf[3615] = 256'h0801030303040306030303000808080001000a0e0c0b0c0a0a0b0a0908040504;
    encBuf[3616] = 256'h0302010102020303000a0f0d0b0a090008000a0b0a0805070403030200080a0b;
    encBuf[3617] = 256'h0e0b0c0a0a0801030303020008090802030503030202010203040303000a0f0e;
    encBuf[3618] = 256'h0c0c0b0b0a080001020203030303020008010204040202040506040302090c0d;
    encBuf[3619] = 256'h0b0c0a0809000008080808000104040303010100020304040201080a0b0d0b0d;
    encBuf[3620] = 256'h0b0d0b0c0a090803040502030102010101010a0c0d0b0b0801020302080a0b09;
    encBuf[3621] = 256'h000403040108000204030300090b0c0a090e0d0e0c0a09000304040101090909;
    encBuf[3622] = 256'h0801030503030008090a08080000000b0e0e0c0b0a0800020302020002040504;
    encBuf[3623] = 256'h0200080909000101080d0d0c0b0a080100000800000205030302030204050202;
    encBuf[3624] = 256'h090d0e0c0a0900010302020000000001080a0d0b0a0105040302080b0d0c0a0a;
    encBuf[3625] = 256'h0a0a080900010205040405030200080b0c0b0a09080008090909010505030208;
    encBuf[3626] = 256'h0a0d0a09000303020a0e0d0c0b0a090104050403030200080a0a0b0d0b0b0b0a;
    encBuf[3627] = 256'h08010203020008000306040302090a0c0a000303010b0f0f0a0a080101020303;
    encBuf[3628] = 256'h05030401080b0d0b0a000203010a0d0c0b0a0001020201000000010100000204;
    encBuf[3629] = 256'h06030401080b0b0d0a0b0a0b0909000101020205040302000c0c0c0908000101;
    encBuf[3630] = 256'h000809090b0a0a09020503080d0f0c0b0a0900020405040304020100090a0a0c;
    encBuf[3631] = 256'h0c0c0b0b0a08030504020108090a090801030301080b0e0d0c0b0a0a09010103;
    encBuf[3632] = 256'h0101010207060304020100090a0a0c0b0d0b0b0a08010303030302020200080a;
    encBuf[3633] = 256'h0d0d0b0a08000301080d0c0b0a0106040203010001000100090c0e0c0c0a0a08;
    encBuf[3634] = 256'h00030503030302020101080b0f0c0b0d0a0a0908000102030404020201010008;
    encBuf[3635] = 256'h0b0b0d0a0a0900010102010008080901040704030201090c0c0c0a0b0c0c0b0b;
    encBuf[3636] = 256'h0a0802040403030202000008090801040604030302090d0c0c0b090901010100;
    encBuf[3637] = 256'h090a0c0c0b0b0a0a000106050403030200080909090800080a0c0c0b0c0a0a08;
    encBuf[3638] = 256'h080108000801050604030301080a0b0b0a0909090b0b0a000403000c0f0f0a0a;
    encBuf[3639] = 256'h080102030302020303060304020109090b0b0c0b0d0d0b0b0a08010404040202;
    encBuf[3640] = 256'h01000009090a0c0b0b0a08080101000001000009090900040706030403020101;
    encBuf[3641] = 256'h090a0e0c0b0b0b0801030302000009000000080a0c0c0b090800010307050303;
    encBuf[3642] = 256'h0200080a0801040201090e0c0a0a00020101090c0a080407040302000a0c0b0c;
    encBuf[3643] = 256'h0b0a0a090808010000020407050403030008090b0a0a0a0c0c0c0b0a08010305;
    encBuf[3644] = 256'h02020200010100000809080102050303000a0f0d0c0b0b090001030404030303;
    encBuf[3645] = 256'h0202020100080b0f0e0b0b0900020503020200090b0c0a0900020202080a0c09;
    encBuf[3646] = 256'h00050504010108090a0a0a0a080003050303000a0c0c0a090003040404030304;
    encBuf[3647] = 256'h01090c0f0b0c0a090000010202030404020300080b0b0c09020405030101090b;
    encBuf[3648] = 256'h0b0b0b0c0c0b0a090105050201090a0a09000302000a0e0c0908010403030202;
    encBuf[3649] = 256'h020403050201090d0d0b0a0900020302000a0c0b0b0a0a090800040505030202;
    encBuf[3650] = 256'h0000080000080a0d0b0a090008090b0a01070602000b0f0b0a08030405020201;
    encBuf[3651] = 256'h0008090a0a0c0a090908090908000307040202080a0b0e0a0b0a0a0908010504;
    encBuf[3652] = 256'h0403020200080809080800000008090c0c0d0c0b0c0b0a0a0902050404030202;
    encBuf[3653] = 256'h08080908000101010a0e0d0c0b0a0808010202030503030301080a0a08010201;
    encBuf[3654] = 256'h090e0e0c0b0c0a090808020305020200080808020405030101090a0909080101;
    encBuf[3655] = 256'h080c0f0e0c0c0c090900030404030302010008080a0a090a0a0b0d0b0c090908;
    encBuf[3656] = 256'h0800010001010101010506040402000008080008080c0e0c0c09090800010000;
    encBuf[3657] = 256'h010204030201000a0a0a08010403000b0f0e0a0a0102050302010a0a0c0a0809;
    encBuf[3658] = 256'h080a0909000305040301000808090a0c0d0c0c0b0a0801030503040202000008;
    encBuf[3659] = 256'h0909080800000a0d0d0d0a09000102000a0c0b09010603030008090803060303;
    encBuf[3660] = 256'h00090c0c0b0b0c0b0b0c0a08000304050303030201000808090a0b0c0c0c0c0a;
    encBuf[3661] = 256'h0a08010304040200080b0c0c0a0900020201080a0b0902070502010809000104;
    encBuf[3662] = 256'h02010b0e0c0b0a0a08080000080009090908050605030301080b0c0b0c0a0909;
    encBuf[3663] = 256'h080a09090a080003050604030301080b0c0b0a0a0a0a09090105040303030000;
    encBuf[3664] = 256'h090a0c0b0a0a0a0e0f0c0c0b0a0003040403030303040201080b0d0c0b0a0908;
    encBuf[3665] = 256'h010008090b0a090204040301000000000008090b0c0901040604030200090b0c;
    encBuf[3666] = 256'h0a0b0b0e0d0b0c09080204030202010204040301000b0c0c0a0900010100090b;
    encBuf[3667] = 256'h0d0b09000206030301080a0c0b0d0b0c0a0a08010405040304010108090a0a09;
    encBuf[3668] = 256'h0808090b0e0b0a090802020304030504030200090a0a0a0a090b0e0c0b0a0909;
    encBuf[3669] = 256'h0808000307060403030101080a0a0b0d0b0b0a0908090a0c0a09010506040303;
    encBuf[3670] = 256'h03010200090a0b0d0b0a090801030201090d0d0c0a080003050201080b0a0902;
    encBuf[3671] = 256'h05040402020008080a0a0c0c0a0a000103020101010405030402020201080d0f;
    encBuf[3672] = 256'h0d0c0b0b09010305030202000001010304030201090b0c0c0b0d0b0c0b0a0002;
    encBuf[3673] = 256'h05030300090a0a0003050303010909090801020200090a0c0b08010200090f0c;
    encBuf[3674] = 256'h0a0902040302080b0d0a090800020405040503020100090a0b0c0c0a0b0a0a0a;
    encBuf[3675] = 256'h0b0900050604030200000808000100080b0d0b09090008080908010604040202;
    encBuf[3676] = 256'h000809090b0c0b09010503020a0f0c0b0a0908000900020704030301090a0a01;
    encBuf[3677] = 256'h050504020208090a0b0b0a0b0b0d0c0c0c0a0a09080103040303030401010808;
    encBuf[3678] = 256'h01020604030201080a090909080b0e0e0b0d0a09090001000101010204050303;
    encBuf[3679] = 256'h0202000809090b0d0e0b0d0a0a0001030504020101080808090808090b0b0c0c;
    encBuf[3680] = 256'h0b0a0909010203040403040404020200080a0a0c0a0b0c0c0b0b0b0a0b0a0a09;
    encBuf[3681] = 256'h0104040503050403040301000a0d0c0b0b090801010201010808080808080a0c;
    encBuf[3682] = 256'h0c0b0a0a08000000010104040302000a0b09010706030301080b0d0c0a0b0b0b;
    encBuf[3683] = 256'h0908030503010a0c0c0b09010203030201000909090a0a0b0d0b0c0901040404;
    encBuf[3684] = 256'h0203030303000d0e0c0b080102000c0e0c0b090803030503020200080a0b0b09;
    encBuf[3685] = 256'h0802030202000a0c0d0d0b0a00030403090e0d0c09000404040100090a0a0a09;
    encBuf[3686] = 256'h080a0b0b0a08030603030100000102040201090c0d0c0b0a09000008090a0b0a;
    encBuf[3687] = 256'h0b0a0908030707050202010009090a090a0b0b0b0a0000000b0f0d0b08030505;
    encBuf[3688] = 256'h030100090a0b0a080002040201080d0d0c0a0a010206030302090a0d0b0a0003;
    encBuf[3689] = 256'h030400090b0a090205050201090b0e0b0b0a0a000001020404040303000a0b0d;
    encBuf[3690] = 256'h0a00010402000a0c0d0a09000103010100090801010108090b0a000505040100;
    encBuf[3691] = 256'h0a0c0a09000100090d0d0b0b090002030100080001060504030302010008080a;
    encBuf[3692] = 256'h0b0f0d0c0b0a0802040402000909090800020201090c0a0a0003050302090d0c;
    encBuf[3693] = 256'h0d0a09080102020203050404030201090b0c0b0b0b0b0a0801040401000a0b0c;
    encBuf[3694] = 256'h0b0e0c0c0b0901050603030100090a090900000101080a0c0c0a090101010009;
    encBuf[3695] = 256'h0901030503000b0c0b00040402080c0d0a09010203010009080800080a0b0e0a;
    encBuf[3696] = 256'h0a0801030605030502030203040303080c0f0e0b0c0909000000010204030303;
    encBuf[3697] = 256'h01080a0b0908010202090b0e0b0a00000202020001020302010a0c0c090a0a0d;
    encBuf[3698] = 256'h0d0b0a00050504030203020201080c0f0c0c0b0c0a0900010404040303020108;
    encBuf[3699] = 256'h090c0b0b09000302000a0e0c0a08020403030009090a08000000090b0d0c0a09;
    encBuf[3700] = 256'h0908000003070605030201090c0c0a09010201000a0d0b0a0002050303010809;
    encBuf[3701] = 256'h090908090a0b0d0a08030604020208080a09000008090c0b0a00050503000a0c;
    encBuf[3702] = 256'h0d0b090802020402030402030108090a0a0a0a0b0c0e0b0c0908030604030200;
    encBuf[3703] = 256'h090b0c0c0a09000003030303030200000009080a0908020402090f0f0b0a0902;
    encBuf[3704] = 256'h040302000008000001000a0c0c0a08020405040303030200080a0b0c0c0d0c0c;
    encBuf[3705] = 256'h0a0a0a0001020304030302020101020304030200090a0c0c0b0a000307020109;
    encBuf[3706] = 256'h0e0c0b0b0a0a0909090002050405030403030200090b0d0b0a08090a0c0d0c0b;
    encBuf[3707] = 256'h0a0901030502030303030403040301080b0d0d0b0b0b0a0a0a08020506030100;
    encBuf[3708] = 256'h0a0a0b080101010a0d0b0b00010201000a0004070503030208090b0b0b0c0a0a;
    encBuf[3709] = 256'h0c0b0d0a080205050202000808090808090b0d0c0b0908010204020303030403;
    encBuf[3710] = 256'h02000a0c0e0a0b08080101000a0b0b0a0900090b0a0804070602020100010002;
    encBuf[3711] = 256'h0201080a0c0c0b0c0c0b0c0b0b09080101000100020506040201080b0d090002;
    encBuf[3712] = 256'h050201090b0c0a08000201010100000000090b0f0d0b0b0a0106040303080b0e;
    encBuf[3713] = 256'h0c0b090801010202020306040202000b0c0d0a0a080101020100090b0c0b0908;
    encBuf[3714] = 256'h01020203040305030201080a0a0b0b0a0c0d0c0b0c0a090102060302080c0d0c;
    encBuf[3715] = 256'h0b0800040305020201080a0c0b0b090104040200090b0c0a0a09090909080205;
    encBuf[3716] = 256'h0404020000090a0909090b0f0c0d0b0b08000205030302020202020303010009;
    encBuf[3717] = 256'h0b0e0c0d0b0b0b09080102040202010109090e0c0b0b0a080103040403030303;
    encBuf[3718] = 256'h02010001010304000b0f0f0d0a09080101010008090908010203030302010102;
    encBuf[3719] = 256'h0200080c0c0b0a0901020401010b0f0e0b0c0b08080001000809080103040304;
    encBuf[3720] = 256'h04030504040202010009090a0d0b0d0b0c0b0b0b0c0909080002040504040302;
    encBuf[3721] = 256'h010009090a09090800010101080b0e0c0b0b08000202080c0d0c090105050502;
    encBuf[3722] = 256'h0200080b0c0b0a0a09080008000801020403040301010100010000000808090c;
    encBuf[3723] = 256'h0e0d0c0b0b0b080001020403030504030402010808090a090a0b0c0d0b0d0a0a;
    encBuf[3724] = 256'h0909010102040404040402030100090b0c0b0c0b0a0a0a0a0a08030706030301;
    encBuf[3725] = 256'h080a0c0b0b0908000102030404030101090b0b0b0a000202000b0f0e0b0a0808;
    encBuf[3726] = 256'h0101020305050403020108090a080000010a0f0d0b0c0a000003020200080001;
    encBuf[3727] = 256'h030603040201020301000b0f0c0c0b0b0a080801020303030100010306040303;
    encBuf[3728] = 256'h0200090c0c0b0a0003060301090d0c0a080102000a0e0c090002050301090909;
    encBuf[3729] = 256'h000404030208090b0c0a0a0900000304020200090a0a0b0a0b0a090a0b0e0d0a;
    encBuf[3730] = 256'h0903070503030301000009090a0b0b08020402090f0e0b0b090004040202090a;
    encBuf[3731] = 256'h0b0b080307040302010008080808090d0c0b0b0902020301090c0b0a00040504;
    encBuf[3732] = 256'h02010808090b0b0b0b08020704030301000a0a0909000008090b0c0b0b0b0a08;
    encBuf[3733] = 256'h03070703020300080c0c0c0c0a0808020202010000010205040303020200080a;
    encBuf[3734] = 256'h0b0b0c0b0d0d0d0b0b0900030403030000080900080103060504030201080b0d;
    encBuf[3735] = 256'h0c0a0a0a080a0a0d0b0a08040604030208090a090801010108090c0a0b0b0a09;
    encBuf[3736] = 256'h08010405030302010100020201010a0d0d0c0b0c0a0a0909090c0c0d0a090104;
    encBuf[3737] = 256'h0504030203040303000a0e0c0b0a08000008090a0a0900020201010808010305;
    encBuf[3738] = 256'h040200000a0908000001080b0d0b0b080206040402000a0e0c0c0b0b09080203;
    encBuf[3739] = 256'h0404040201000000010100080b0f0c0c0a0a0908000101020303030101020406;
    encBuf[3740] = 256'h030401080c0d0b0b0a090a080909000002020302050504040201090c0c0b0909;
    encBuf[3741] = 256'h0000080a0c0a0a010505040201090b0d0b0900020201080a0a0a080304040101;
    encBuf[3742] = 256'h00080a0b0d0d0b0a090803040503020108090b090a090a0d0e0c0c0a09000306;
    encBuf[3743] = 256'h0404030201080a0b0b0b0b0a0b0b0e0b0c0a09010404040302020008090a0b09;
    encBuf[3744] = 256'h09090008090a0c0b0b080307040201090c0c0a0900010201080a0c0b09010403;
    encBuf[3745] = 256'h0401000a0b0b0908080b0f0d0b0c09010306030301010001020402080c0f0c0b;
    encBuf[3746] = 256'h0b090000010102010303040100090b0c0a090802010100090b0b090003060303;
    encBuf[3747] = 256'h03030402000b0f0e0b0c0a090900000001040604040201080b0c0c0a09080000;
    encBuf[3748] = 256'h00090a09080104040302000101020302090e0d0d0b090800010208090a0a0803;
    encBuf[3749] = 256'h0706030202080a0b0d0b0a0a0908090000020404020200080800010302080c0f;
    encBuf[3750] = 256'h0c0b0a090002040403020200080a09090001040402000b0f0e0b0a0800020402;
    encBuf[3751] = 256'h020200000800080808080b0d0a0902060303000a0b0a0808090d0e0b0a000404;
    encBuf[3752] = 256'h04020203020201090f0c0b0b0a09000101020305020302010101080b0f0c0c09;
    encBuf[3753] = 256'h0900010000010204040302000a0b0b0b090100080c0e0c0b0a00050604030201;
    encBuf[3754] = 256'h01080008090c0d0d0b0c0908000102020303030402020208090c0b0a09030703;
    encBuf[3755] = 256'h01080b0d0b09010201090c0d0a0a000203040201000000000002040405030302;
    encBuf[3756] = 256'h01080c0e0d0c0b0b09090001030404040203010108090a0a0a09090808080809;
    encBuf[3757] = 256'h0a0a0c0a0b090003060503020200000000090a0f0c0c0b080205050302020808;
    encBuf[3758] = 256'h0a0a09080101000b0f0c0b0a0003040401000809080103030401010201040202;
    encBuf[3759] = 256'h000c0e0d0b0b0b090001010202020205040303030100080908090b0d0c0b0801;
    encBuf[3760] = 256'h040502010a0c0c0c0a08000305040201080b0e0c0a0802040404030200090a0b;
    encBuf[3761] = 256'h0c0b0b0a0b0a09080002050404030303040201090c0d0b09080204030200090c;
    encBuf[3762] = 256'h0c0c0b0a08010305020201010001020100090c0d0b0b0901030703040100090a;
    encBuf[3763] = 256'h0b0b0c0b0c0b09000307050302020009090b0b0d0b0a09080204030200090c0b;
    encBuf[3764] = 256'h0b0a00040403040202020202090b0e0c0a09080000090b0b0a00060503030109;
    encBuf[3765] = 256'h0b0d0b0a08000202020201000202000108000405050200090d0d0c0a0b090908;
    encBuf[3766] = 256'h0002040403040202010101000000090d0e0c0d0a090002040202000808010103;
    encBuf[3767] = 256'h02090d0e0b0b0a09000202030304030503030201090c0c0c0c0a0a0a090a0900;
    encBuf[3768] = 256'h000203040304030303020108080a0b0d0d0d0b0d0a0908010304040202000808;
    encBuf[3769] = 256'h0908000008090b0c0b090808090d0d0b0b08030703030200090b0b0c09090002;
    encBuf[3770] = 256'h04040202080c0d0c0a0802040401080b0c0b0a0901020100080a090001020208;
    encBuf[3771] = 256'h0b0c090206050201080a0b0b0a0b0b0e0d0c0b0a0802050402010a0e0c0b0900;
    encBuf[3772] = 256'h01040303030301000009090c0d0d0b0c0b09080204020300080a090900010202;
    encBuf[3773] = 256'h01000009080a0a0d0c0c0c0b080206050301090c0e0b0a090801020202020101;
    encBuf[3774] = 256'h0102040303000a0f0d0b0b0a08000001010000080a0d0c0b0901070404020008;
    encBuf[3775] = 256'h0a0c0a0a0900010101080b0e0c0a0a0808010102040504020200090a0c0b0a09;
    encBuf[3776] = 256'h080908090b0c0b0b09010603040200000808090a0d0b0a0a0803040403010201;
    encBuf[3777] = 256'h0108080d0c0c0c0b0a0a0a0a08010404060304030303000b0f0c0c0a08080101;
    encBuf[3778] = 256'h010008000002010008000103050300080c0a09080102090c0d0e0b0b0a000505;
    encBuf[3779] = 256'h040201080a0b0b0a0808000a0a0a0901040505030303030108080b0b0c0c0c0b;
    encBuf[3780] = 256'h0c0c0a0b0a00030704020301080000000100090c0d0a090103040200090a0a08;
    encBuf[3781] = 256'h0000080a0c0c090802050403020301020002020201010a0b0c0a08080a0e0d0c;
    encBuf[3782] = 256'h0a090000000001060504040200080a0a0801020200080909080000000b0f0e0b;
    encBuf[3783] = 256'h0a00040704030108090b0c0a0900010203040201080a0d0b0b09010307030301;
    encBuf[3784] = 256'h000808080001080b0d0d0a09000204040303040302000a0e0c0b0b0900020201;
    encBuf[3785] = 256'h010001030604040302020000090a0b0e0b0d0b0b0a0801030603040201000008;
    encBuf[3786] = 256'h00020202010009090c0b0e0c0b0b0a08020305040203030203020108090d0d0c;
    encBuf[3787] = 256'h0b0a090104060304020108090b0b0b0b0909000000080b0e0c0a080106050403;
    encBuf[3788] = 256'h03030202080a0b0e0b0a0909090b0e0c0a0a0803050503030202000009090909;
    encBuf[3789] = 256'h0a0a0b0d0b0b0a08000201020204030502010000000201010a0d0d0b0b090103;
    encBuf[3790] = 256'h060403030100090d0c0b0c0a09080801020203030302030406040302010a0e0c;
    encBuf[3791] = 256'h0b0c0a0908010002010100020305030200090a0909000801080a0a0c0d0e0c0c;
    encBuf[3792] = 256'h0a0900020306030402020009090b0a0a0a0c0d0b0b0801040403000009080001;
    encBuf[3793] = 256'h00080b0b0c090808090c0b0c090104040503040201080b0f0c0b0a0900010101;
    encBuf[3794] = 256'h00090008020305030401000a0e0c0c0a090002020302000a0d0c0b0900020503;
    encBuf[3795] = 256'h020109090a0909080a0a0c0b09080001000b0c0e0a080205040308090e0b0a08;
    encBuf[3796] = 256'h0103030108090a09080a0c0f0b0c0a000102040202020100080a0e0c0b0a0900;
    encBuf[3797] = 256'h02030308090c0a0901000a0f0f0c0b0a0902040403030100080909090909090b;
    encBuf[3798] = 256'h0c0d0b0c0b0a0800010108080003060402080a0d0b090003030301090a0d0c0c;
    encBuf[3799] = 256'h0b0a09080108080a0a0a0a09090a0005050502010808090800080c0d0e0b0a00;
    encBuf[3800] = 256'h010301090d0d0a0801030401080a0b0b080203020008080a0a0f0f0c0c0b0901;
    encBuf[3801] = 256'h0405030201090a0a0a08010208090c0c0a0809090b0f0d0a0901020302010101;
    encBuf[3802] = 256'h0406040301090b0e0a0a08010001090c0c0b090802030301080b0a0001040402;
    encBuf[3803] = 256'h02030203010009090b0a0c0d0d0d0b0c09080103040301080b0b0c0801010200;
    encBuf[3804] = 256'h09090307070301000b0c0a09010303080b0f0b0b080002020201000101020101;
    encBuf[3805] = 256'h00090808090908010606030302090a0a0900000a0f0d0c0b0900010403050202;
    encBuf[3806] = 256'h01010008080b0c0e0c0a0900030503040101010201020208090c0b0b0a090a0c;
    encBuf[3807] = 256'h0e0b0c090003040302000001040704030301090a0b0d0a0a0a08000002030405;
    encBuf[3808] = 256'h040202000a0b0d0b0a090909090a090307050403030100080a0a0a0801030303;
    encBuf[3809] = 256'h000b0f0d0c0a0900010202020102030403030202010201000a0d0d0a08000303;
    encBuf[3810] = 256'h0402020202000c0f0d0b0a0901030405030202020009090a0908030603030108;
    encBuf[3811] = 256'h0a0d0d0a0a090003050202000a0a09080205040304010100080a080801040303;
    encBuf[3812] = 256'h080c0f0c0b0b0901030502030101020304040202000808090b0d0c0c0b0b0900;
    encBuf[3813] = 256'h010203050201000a0a0903070705020100090a0a0a0a0a0b0a0b090800010001;
    encBuf[3814] = 256'h02050404040203020100080808000202000c0f0b0c0b09080909090901050505;
    encBuf[3815] = 256'h030101000909080800080909080801030303080b0f0d0c0c0a0a000204030401;
    encBuf[3816] = 256'h020101030303040200090b0d0a0b0c0b0e0d0c0b0b0901030604020201000108;
    encBuf[3817] = 256'h00010008080b0c0b0b0b09090b0c0b0b08020304000909000506040202080809;
    encBuf[3818] = 256'h090909080900010402000d0e0c0c0a0b0a09080203060304020101010101080a;
    encBuf[3819] = 256'h0c0d0b0b0c0b0a09080203030300000304050401080a0b0c09090a0d0d0b0900;
    encBuf[3820] = 256'h03050300090c0b0a0003060302080a0d0b0a09020201000b0d0b090002020108;
    encBuf[3821] = 256'h090909080a0a0a0903050401000a000305020b0f0f0e0a090800010302020008;
    encBuf[3822] = 256'h0a0a0802040301090c0a080102080f0f0b0c09080103030303030108090b0a0b;
    encBuf[3823] = 256'h0a0a0d0c0c090801040202080a0b0b0a0b0c0b0c0900030603020109090b0c0c;
    encBuf[3824] = 256'h0a09010405040100090c0b0a0a09090b0d0c0c0a090801020306040304020100;
    encBuf[3825] = 256'h0a0d0b0c0b09090908090800010403030108090a000205030108090c0a0b0c0d;
    encBuf[3826] = 256'h0d0c0b0a0800040403030200080b0a0909000108090b0e0b0b0b0a0802050402;
    encBuf[3827] = 256'h01090c0a0902040301090b0d0a08080a0a0d0b0909080108020605040401080b;
    encBuf[3828] = 256'h0e0b0b0900010403050201000a0c0d0b0c0a0a08000203040303030202010008;
    encBuf[3829] = 256'h0a0c0b0a0b0a090c0c0c0b0b0a0a0909080207050404020100090b0c0c0a0900;
    encBuf[3830] = 256'h00020200000800020303020a0f0d0b0b0908000008080103070503030201080a;
    encBuf[3831] = 256'h0c0c0b0b0a0a0a0c0a0a0803060403010008090003040403010a0d0f0b0b0908;
    encBuf[3832] = 256'h010303020008000102040208080b0c09090a0909000406050301090a0d0b0a0b;
    encBuf[3833] = 256'h090a0b0c0909010404040403020402020401010a0d0d0b0b090908090a0a0803;
    encBuf[3834] = 256'h060502010008080103040302090c0d0c0b0b0a09000104050302020009090a08;
    encBuf[3835] = 256'h02040402000b0c0d0b09090800000002040403020100080001080a0e0d0a0a00;
    encBuf[3836] = 256'h02040302020201020008080808000a0f0c0d0a09080000080802030705020304;
    encBuf[3837] = 256'h02020201080a0d0c0b0d0a0a0a08000104030504020300080a0b0b0b0909090a;
    encBuf[3838] = 256'h0a090207050402020001080000000a0b0c0c0a0a09090b0b0b0a020706040303;
    encBuf[3839] = 256'h0202000909090a0a0a0a0b0b0d0b0b08010306030303030504040301080c0e0b;
    encBuf[3840] = 256'h0c09080103030302010202050302080a0d0d0a0a090908080808010504050303;
    encBuf[3841] = 256'h0202000909090c0b0e0b0c0909000202020305030502020200000808090a0d0c;
    encBuf[3842] = 256'h0b0b0a0909090900010505040303020201020100080b0e0c0c0b0a0802040403;
    encBuf[3843] = 256'h02010008080909090a0c0c0b0b090103070304040203010100090a0a0c0b0b0b;
    encBuf[3844] = 256'h0b090a0a0c0b0b0901060505030503020201090a0b0d0a0b0a0a090802040304;
    encBuf[3845] = 256'h00080808000203030402090b0f0c0b0a0003050303010203030302080d0a0a0a;
    encBuf[3846] = 256'h0b0f0e0c0a0a00030504030201000009090a0a090808090a0a0b0c0801010403;
    encBuf[3847] = 256'h0305030201090d0b0c0b09080104040303000a0c0b0901040301080b0c0a0800;
    encBuf[3848] = 256'h000a0b0d0a08010306030203020000000003010a0f0f0c0b0b0a080008000103;
    encBuf[3849] = 256'h0705020201090a0b0b0a080802040302080e0d0c0b0a0802030303030108090c;
    encBuf[3850] = 256'h0d0b09080202030101000101090d0e0b0a08010201090c0c0b08080001080008;
    encBuf[3851] = 256'h090c0d0c0c09080002030505030302090c0e0b0a09010001090b0e0b0b0a0908;
    encBuf[3852] = 256'h000304030301090c0b08030506030201080b0d0d0c0b0a090808080809080001;
    encBuf[3853] = 256'h01040405040302080c0d0b0b09090008080808000101020201010201010a0e0e;
    encBuf[3854] = 256'h0c0c0a0b0908020504030200090c0b0b0b0a0808000100000a0d0c0b09010406;
    encBuf[3855] = 256'h03030201090b0e0c0b0b0908010100090c0d0b0a0a08030705030301000b0c0c;
    encBuf[3856] = 256'h0a0a09080000010100080a0b0c0a0a00010200080a080802050403040201000a;
    encBuf[3857] = 256'h0c0c0d0c0b0d0b0b0900020202080c0b0a02070503030300080a0d0c0b0c0a09;
    encBuf[3858] = 256'h090808000801000202030404030201090c0c0b09090809080b0b0c0c0b0c0b0b;
    encBuf[3859] = 256'h0802060503020209090a0b0b090a09010003040108090e0c0b0d0a0a0a000102;
    encBuf[3860] = 256'h010208010505040400080a0c0b0a0a09090b0c0909020604040300000a0d0b0a;
    encBuf[3861] = 256'h0a080102030300080a0e0b0a0901050503030108080b0a090a09000900010d0e;
    encBuf[3862] = 256'h0d0c0a090105040303020000080a0909080001090a0b0f0a0a0a0b0a09010705;
    encBuf[3863] = 256'h0403020000090a090a0a0b0a09000101030003060405030201000a0b0a0c0b0b;
    encBuf[3864] = 256'h0d0b0a0a0004040503020101020305040201080a0c0b0c0a0a0b0a0c0b0a0902;
    encBuf[3865] = 256'h070405040202020009090a0b0b0c0b0a0a090001040403030302010001020503;
    encBuf[3866] = 256'h03020a0e0c0c0a090000020203030503030300090b0c0b090801000100000105;
    encBuf[3867] = 256'h050404020100080a090801020302000b0c0c0b0c0a0a00060704040100080a0a;
    encBuf[3868] = 256'h090802030303020200080c0d0b0c09010404050200080a0c0a08010303020000;
    encBuf[3869] = 256'h0801030504020202030202080c0f0d0b0a090104040301010009080002030402;
    encBuf[3870] = 256'h0108090b0c0b0a0908020504030202010203070302000b0d0a0a00020200080a;
    encBuf[3871] = 256'h09010405040201000000030502030109090a0902060304010a0c0d0b0a010104;
    encBuf[3872] = 256'h030102030306030101000002040101090d0c0a0b0b0a0902070504030100090a;
    encBuf[3873] = 256'h090909080908010305040202010208080b0e0b0a080203020303020603020200;
    encBuf[3874] = 256'h09000108000b0f0c0908020303050200080b0f0a0a0006030402000a0a090a00;
    encBuf[3875] = 256'h01080404040501090b0e0c09090801080801020206020100000001010000090e;
    encBuf[3876] = 256'h0b0d0c0a0a000205030202090a0a0b090809000103050401000a0b0b0b0a090a;
    encBuf[3877] = 256'h0a0a0a0c09090a030703060301000a0d0b0d0c0a090802020403030101010202;
    encBuf[3878] = 256'h000d0f0c0c0b0909000001020304030100080909020303020a0f0d0d0b0b0b0a;
    encBuf[3879] = 256'h00020403040102000000080b0b0d0b0b0a0c0b0c0a000206040201000809090a;
    encBuf[3880] = 256'h0c0c0b0a08000101080b0c0a0a080a0b0a0802070403010108090b0f0b0d0b09;
    encBuf[3881] = 256'h080000080a0b0c0a010204040302000a0f0c0b0b0800010100000808090a0d0d;
    encBuf[3882] = 256'h0b0a00030402000a0d0c0b0a0b09080204040201080a0909090c0f0d0c0b0a08;
    encBuf[3883] = 256'h0102020101010103030301090a0c0c0d0b0d0a0b0a0a0b0b0a0a000203020809;
    encBuf[3884] = 256'h09020604030100080b0c0c0d0c0b0c0a09090909080003040301090b0c0d0b0b;
    encBuf[3885] = 256'h0d0b0a0908010008080900070305020100080a0b0e0d0c0b0b0b08090a090801;
    encBuf[3886] = 256'h0605040303010109090c0d0c0b0b0a0808000001030304030201000100020200;
    encBuf[3887] = 256'h0a0c0e0c0b0d0c0a0a09080101020203060303030000000808000b0f0c0c0a0b;
    encBuf[3888] = 256'h090a080801050404030108090a0a0909090009090a0c0c0a0901040503040202;
    encBuf[3889] = 256'h030201090d0f0b0a0a000001020001010000000800020102030809090b080301;
    encBuf[3890] = 256'h05050404050200090d0b0c0a0900080001080001080002030704040202000908;
    encBuf[3891] = 256'h0802020200080d0b0b0c0b0b0d09080205050304030101080b0b0a0901030000;
    encBuf[3892] = 256'h090b0006040302000801020505010108090a090a090a0b0a090a020606060404;
    encBuf[3893] = 256'h03020008080a0a0b0c0c0b0b0901020504040203020102000203030401090d0c;
    encBuf[3894] = 256'h0d0a0a08080000000000000304070305030302030100080b0c0c0b0b0a080000;
    encBuf[3895] = 256'h00090a0b0a0903070704030203010808080001020200080b0c0d0a0908000103;
    encBuf[3896] = 256'h04030201080c0c0c09000405050304020201000809090909080909090b0c0b0b;
    encBuf[3897] = 256'h0a0207040403010100090808010305040304020100080b0c0c0a090002030402;
    encBuf[3898] = 256'h0008080908020206030503030302000808080001020008080b08000901000207;
    encBuf[3899] = 256'h070503030201080b09090105050303020808090801040102080a080105050300;
    encBuf[3900] = 256'h0a0d0c090003060302020101050403050200090b0d0b0c0a0a0a0a0900020703;
    encBuf[3901] = 256'h0403030202020103010008090b0b0e0d0b0c0b0a090800010104030604030302;
    encBuf[3902] = 256'h0008080a0908010202080a0c0c0b09000002080a09090902000d0c0c0a010605;
    encBuf[3903] = 256'h050303020109090a0a0800010401090b0e0d0b0a0b0900000304020302010302;
    encBuf[3904] = 256'h030402010402040402090b0f0d0a0a0900000808090a08000803030306020304;
    encBuf[3905] = 256'h030303000b0d0d0c0a090000000a0b0e0c09090801010304040304020100090a;
    encBuf[3906] = 256'h0b0c0d0a0a0c0a0c0b0b0a0802040305020002000001000808090b0c0e0c0b0b;
    encBuf[3907] = 256'h0a090008080a0c09090900080b0a0b0b08080801080b0809020707030300090d;
    encBuf[3908] = 256'h0e0c0b0c0a0b0a0b0a0909090a0908000405040203020101000a0b0f0d0c0a0b;
    encBuf[3909] = 256'h0a0a090a090b090908010204030201080c0c0c0d0a0a090a090a0b0b0c0a0909;
    encBuf[3910] = 256'h08090900010205010b0f0f0c0b0b0908010101090c0c0b0b0908000103030202;
    encBuf[3911] = 256'h08090d0c0c0b0c0b0b0b0909090a0f0d0b0b0a0002030401080a0c0b0c0a0800;
    encBuf[3912] = 256'h0000000a0c0c0c0b0b0c0a0a0800020200080d0d0b0b0b09090001090c0b0f0b;
    encBuf[3913] = 256'h0a0b0a090a09000205050201090c0c0b0c09000808080c0c0b0d0b0909000101;
    encBuf[3914] = 256'h010301020301090c0f0c0b0b090000020300090a0d0a090900010a0a0a0f0b09;
    encBuf[3915] = 256'h0b0b090b0a090d09000104050108080d0a080804040202000b0c0b0f0a0a0c09;
    encBuf[3916] = 256'h090800030203020a0b0b0c08060403040108080b0c0a0c0b090a010403030400;
    encBuf[3917] = 256'h090a0c0a09080306030202090c0b0d0a00000305010202000000090801000307;
    encBuf[3918] = 256'h020302090b0c0d0b0909010303040301010301050502040402020308090a0c0b;
    encBuf[3919] = 256'h090902040204030101000b0a0103070703020108000000020302040302030300;
    encBuf[3920] = 256'h09090b0802050605020302080808090207040403020000090800080101010405;
    encBuf[3921] = 256'h0305030201000909080803060304020100080003050404020201010001000001;
    encBuf[3922] = 256'h0202040203040403040202020305050404020100090909000102030401020008;
    encBuf[3923] = 256'h0001060504040303020202010008080808080100000809080204070703050203;
    encBuf[3924] = 256'h0202000808080801000101000200080001000407040603020301000808090001;
    encBuf[3925] = 256'h0105020101000b08090904060305040203020101010909080b01020305020900;
    encBuf[3926] = 256'h0a0a02060307030202020002010801010904030206010808090b010108040209;
    encBuf[3927] = 256'h030201070402040301040201020209010a0d080a0b02000a0301090603010703;
    encBuf[3928] = 256'h0104010003000900090d08090a03030204000c09090b05030206030103010a00;
    encBuf[3929] = 256'h0c0f080909010200030109080b0e08000904020105020001090e090b0c080000;
    encBuf[3930] = 256'h03030003000a080c0d08090a01090d090b0e08080a02010006020102010b080c;
    encBuf[3931] = 256'h0d090c0b0a0a0a020008000c0e090a0a020100040109000b0e090b0d090b0a08;
    encBuf[3932] = 256'h00000401090a0d0e0a0b0a00080801080a000c0d0a0b0c090909000809080a0d;
    encBuf[3933] = 256'h0a0e0b0a0a09010008080b0e0a0d0b0b0c0b08090900090c0b0d0b0a0c0a090a;
    encBuf[3934] = 256'h09000808080b0d0b0e0b0b0b0c090a09090c0d0c0c0b0b0a0909000001000809;
    encBuf[3935] = 256'h0e0c0b0c0b090809090a0a0b0d0c0b0b0b0b0b090b0b0b0c0c0c0b0d0b0c0a0a;
    encBuf[3936] = 256'h090a090b0b0a0d0b0b0c0c0a0a0b09090a090c0b0b0d0b0c0d0b0a0c0b0a0b0b;
    encBuf[3937] = 256'h0a0b0c0a0b0b090b0a000a0d0b0e0c0a0c0a090b0a090b0a090c0c0a0e0a090a;
    encBuf[3938] = 256'h090a0c0b0a0c0b090b0b080a0a000b09090e0a090c0d0a0d0b0a0c0b090a0a00;
    encBuf[3939] = 256'h0a0a080d0c090b0b000908010a0b090f0c0a0c0a0a0b09080a0a000c0b090d09;
    encBuf[3940] = 256'h080a08000c0b0a0f0b080a09000b0b0a0f0b080b09010900030900030c0b0a0f;
    encBuf[3941] = 256'h0a080b0a010b0a080f0c090d0a000901030001020a09080c09010900040a0902;
    encBuf[3942] = 256'h0e09000c09080c0a010802050808090f09000801040102030002040908000c08;
    encBuf[3943] = 256'h010a00030901060a0a010c00040206040002030102030808020b010600020309;
    encBuf[3944] = 256'h0004000306000203010307010305010203080002090103010405010304000203;
    encBuf[3945] = 256'h0003050306040203030000020802040103050203040002020801030205050304;
    encBuf[3946] = 256'h040202010002030206040203030102010808080a010404050502030302030201;
    encBuf[3947] = 256'h0203040405020102000000000203040504030303030101020403030503010302;
    encBuf[3948] = 256'h0203030304050305030403020203020203040306020203000100010303050403;
    encBuf[3949] = 256'h0403030303040303030403030203060203030203030304030304030203050304;
    encBuf[3950] = 256'h0303040304030401030301040302040301020300020401030402060302040401;
    encBuf[3951] = 256'h0302010302010203080304000203040602020403010403000402000303000402;
    encBuf[3952] = 256'h0803010806040104020002020803020804030107020001080902020005020805;
    encBuf[3953] = 256'h020104010901010803020804030007030801080d00010804030003010b01090f;
    encBuf[3954] = 256'h00010004030104010903080b000b0e01030005010a000a0e08090b0001000703;
    encBuf[3955] = 256'h0802080b09090a01090d01080a01000c080a0c03010904000e08080a080b0e00;
    encBuf[3956] = 256'h080a01000b01090d01080c09090d010809010d0d090a0a00010900080a02090d;
    encBuf[3957] = 256'h000b0f09080908090b090a0b080f0d0a0a0a01010001000a090a0d080c0c0008;
    encBuf[3958] = 256'h0900090f0b0c0c090a0a09080901010002090d090a0a080a0c090b0f0a0d0d0a;
    encBuf[3959] = 256'h0a0a000008000008000009090f0b0b090a00090b0c0e0c0a0a0b090a09000008;
    encBuf[3960] = 256'h080a0c09090a000a0d0b0c0c090b0d0b0d0b0b0a0a090b0c090a080800090008;
    encBuf[3961] = 256'h090a0d0c0b0c0d0a0a0a0c0c0b0a0a0b090a0b090a08080a0a0c0c0b0b0d0a0b;
    encBuf[3962] = 256'h0d0a09090a0c0d0c0b0a0b09090a08080009090a0e0c0b0c0a08090a0a0b0c0c;
    encBuf[3963] = 256'h0c0c0b0c0b09090002010808090c0c0c0b0b0b090009090a0d0e0a0c0a080908;
    encBuf[3964] = 256'h08080a090c0c0b0c0a09080800090a00080a090e0c0a0a0b08090c0b0e0c0a0a;
    encBuf[3965] = 256'h0908090002000001090b0b0e0a08090a0a0b0c0a0c0c0a0d0c080a0001000009;
    encBuf[3966] = 256'h0c0a080b0a080a09030000080d0c0b0c0b0a0c09000909020909080b0a010003;
    encBuf[3967] = 256'h060000020a0c0b0f0c0a0b0808000801090801010304080003000404000c0a0d;
    encBuf[3968] = 256'h0b0b0c0b0a0a09020204030008010003050808080a010500080a0f0b0a090900;
    encBuf[3969] = 256'h0a00030206030009080a00030101000801040000090f0b0a0a00030102050202;
    encBuf[3970] = 256'h03090b0d0c09010205030100030000080f0c0a09020503030308090a0d0c0a0a;
    encBuf[3971] = 256'h01030504040000090909080909000205040201000b0d0a080001010304010303;
    encBuf[3972] = 256'h090b0a0c090104070301030308090b0f0b090902040203020100010908080904;
    encBuf[3973] = 256'h07030402000b0a0d0a090a08010205050202000909000001020102020008080d;
    encBuf[3974] = 256'h0b0a0901040204030102050100000909010106040008000908000908010a0802;
    encBuf[3975] = 256'h010304000104030404010103010202090b0d0c0a000203050100010101030203;
    encBuf[3976] = 256'h030306030200080a090800020501000202030401000008020302020302010200;
    encBuf[3977] = 256'h030402030603020100090a090005030303010202010201000004040403020000;
    encBuf[3978] = 256'h0908030303030407030200080b0d08000204040303020201080a0a0a01070405;
    encBuf[3979] = 256'h02010100090a0b0b0a08040605030200000909090801020505030302000a0b0b;
    encBuf[3980] = 256'h0a0a0103060403040201090b0c080204060302020200090b0b0c090802050403;
    encBuf[3981] = 256'h0201010009090a0804070403020108090b0b0c09090203070303020108090908;
    encBuf[3982] = 256'h0002020405030402080a0b0d0a000002040304040201010a0b0a080103060303;
    encBuf[3983] = 256'h030202080b0d0c0900030405020102020008090c0a0802060304020009000a0b;
    encBuf[3984] = 256'h08000004060304020000090a09090b08080207030303080a0a0a0a0204030604;
    encBuf[3985] = 256'h0203080b0b0d0b000001040201050200080a0c0a080105030102080908090d08;
    encBuf[3986] = 256'h080802030104000a08080a08090b01010107030201000a0b0b0b00010801000a;
    encBuf[3987] = 256'h090b0e0a090004030306020000000b0b0c0c090800040200080b0d090a090003;
    encBuf[3988] = 256'h04060400000a0c0a0a0a01010002010800090d0a0c0b0000000403020301090a;
    encBuf[3989] = 256'h0b0d0b0b0c00000802010b0a0b0d0a0a0b01030405020101080d0b0d0c090a09;
    encBuf[3990] = 256'h01030201080b0a0b0d09090b02020103080d0a0b0f0a090a080001020401010a;
    encBuf[3991] = 256'h0f0b0a0b0a080902010103000e0b0c0e0a0908000203020109080d0e0a090a00;
    encBuf[3992] = 256'h010101010a0b0e0d0a0b0b09000205030100090d0b0b0c0909000102080a0c0e;
    encBuf[3993] = 256'h0a0b0b0a0a0801030305010a0c0d0c0a0a0908000001080a0a0e0d0b0b0a0a08;
    encBuf[3994] = 256'h00030201080b0e0c0b0b090908000009090e0c0c0b0b0b0a0a0800010201080a;
    encBuf[3995] = 256'h0e0c0b0b0a0a0a090a0c0c0b0d0a0b0a090a090900090008090b0d0d0b0b0c0a;
    encBuf[3996] = 256'h0b08090809090c0c0c0b0b0a090101090a0b0c0c0a0c0b0b0b0a0a0a0b0a0d0c;
    encBuf[3997] = 256'h0a0a0b0c0b0a09090001090a0b0e0a0a0b0a0b0b0d080b0b0b0c0b0b0f0a0808;
    encBuf[3998] = 256'h00010000090e0b0c0c0b090a09000809010a090a0c08000b0a080b0a080e0b0b;
    encBuf[3999] = 256'h0c0b0a0b0801010204080a0a0e0900080002090a080d0c090c0b090900030000;
    encBuf[4000] = 256'h030800000d0a080c09020102040809090f0a090b09020803050001010b0a000c;
    encBuf[4001] = 256'h09020002030808090d0b090d00020801030103040800000d0900090002000304;
    encBuf[4002] = 256'h0001080d0a080b01060202010000020900020900020801050102030808020b0a;
    encBuf[4003] = 256'h000802040103060101040001010800030003050102040809080b000304060402;
    encBuf[4004] = 256'h0302000000080102000303020306010202000102010305020503030402080900;
    encBuf[4005] = 256'h0802050303040303030202020a08000004060305030201000900000205050201;
    encBuf[4006] = 256'h0100010800000202040503040303030201010809010403040403020302030403;
    encBuf[4007] = 256'h0502030303040403040100080000030405040304030102000001020203030401;
    encBuf[4008] = 256'h0305020204020302030602020304010202000103050403020201000101030403;
    encBuf[4009] = 256'h0403000104020305020203030303020203020103020003010306020102080104;
    encBuf[4010] = 256'h0304040100010008020101040100020101040203070201010800020203050100;
    encBuf[4011] = 256'h02080801080803020103000803010205020104010104010203000a0100080200;
    encBuf[4012] = 256'h0802080902000004000804020306020001000002000900090b01080902010004;
    encBuf[4013] = 256'h020104010801080801080a010100050000000b0a000800020100020100050108;
    encBuf[4014] = 256'h000b0c090b0a03030307010808090b08080802000902000902000a0808090301;
    encBuf[4015] = 256'h0002000a08080a010a0b080808010109000808010009010a0b090b0d09090802;
    encBuf[4016] = 256'h020201080b09090a00080a09090a09090a090b0e09090801020101090b0a0a0c;
    encBuf[4017] = 256'h090b0c0a0a0a0a090b09090b00090c0a0a0a010108090c0d0b0b0a0908090800;
    encBuf[4018] = 256'h0b090c0d0b0b0c09080900010908080c0a0c0c0b0a0b0a0a0c0a0b0d0b0a0c09;
    encBuf[4019] = 256'h090a09090a0a090c0a0a0e0b0b0c0b0a0b0a0a0b0b0b0b0b0a0b0b0b0b0b080b;
    encBuf[4020] = 256'h0c0c0d0b0a0b0a090b0b0b0d0a090a0a0a0c0d0b0b0a0808080a0b0e0b0c0b0a;
    encBuf[4021] = 256'h0b0c0a0b0a0a0b0d0a0a0b0a090c09090908090b0f0b0d0a0b0a0a0a0b0a0908;
    encBuf[4022] = 256'h000108090b0d0b0b0d0b0a0b0c0a0b0b0b0c0a0a0b09090a09090b0c0b0e0a0b;
    encBuf[4023] = 256'h0a0a0a0a0a080b0a0a0b0b090c0b090d0a090b0b0b0e0a08080802080a080b0b;
    encBuf[4024] = 256'h090c0a0a0e0b0b0b0a08090801080002080000090a080b0e0a0d0b0909000201;
    encBuf[4025] = 256'h01010808020000010b0b0a0d0b090b0a080a09020002060100010a0a090b0a01;
    encBuf[4026] = 256'h0a09020a08000909010003050101020809010b0c0a0c0a000801070102040100;
    encBuf[4027] = 256'h02090001090002080902080802080205020305010002010103000a080b090403;
    encBuf[4028] = 256'h0505010202000102000102080804020405010101080103020205000204020404;
    encBuf[4029] = 256'h0202020101010a09010104060303030302020100010808020004060305030203;
    encBuf[4030] = 256'h010808090a0901000404020304030505020301000000080008090a0000040703;
    encBuf[4031] = 256'h0304030201010800080000000008000205030503020303040403020200010009;
    encBuf[4032] = 256'h0a0b0b0a0908010405060305020201000008080a0b0b0b0b0003070403030302;
    encBuf[4033] = 256'h010008090a0b0a09010104020404040304020100080b0b0d0c0a090004050303;
    encBuf[4034] = 256'h030101080b0b0d0a09010306030101090b0c0b0b010203060303040201080a0e;
    encBuf[4035] = 256'h0b0b0a090808020204050402030100000b0e0b0c0c0908080204040403010109;
    encBuf[4036] = 256'h0c0b0c0a0a080800020204030202020100000b0c0d0d0b0b0c09080005030403;
    encBuf[4037] = 256'h020001080808080b0b0b0f090a0b0b0d0c0909010404040403030201090b0e0c;
    encBuf[4038] = 256'h0b0b0c0a0909010304050303020201080a0e0c0b0b0a09080103030502020200;
    encBuf[4039] = 256'h090a0a0c090809000009000101030309090c0b0a0a0c0b0b0b04070403020008;
    encBuf[4040] = 256'h0a0c0b0d0b0a000406040201090a0d0b0c0a090802040503030200080a0c0b0d;
    encBuf[4041] = 256'h0a090900020203030201010008080909090a0a090b0908030705030401080a0c;
    encBuf[4042] = 256'h0d0b0c0a0a0001050403030201010809090a0b0a0b0d0c0b0b0b090002050305;
    encBuf[4043] = 256'h040303040102010808090c0d0d0c0b0b0a08000306040304030101000a0b0c0c;
    encBuf[4044] = 256'h0b0c0a0908010303050303020301090b0f0b0b0a0800020305030302080a0d0b;
    encBuf[4045] = 256'h0b0a0900010204040302000a0a09080101080b0d0a0a00000808090802010a0a;
    encBuf[4046] = 256'h0f0a00050604030202080a0d0e0c0b0a0a0103040503020100090b0c0d0a0a08;
    encBuf[4047] = 256'h01020202010100010008080909080a0d0f0c0b0a0003050404020100080b0d0d;
    encBuf[4048] = 256'h0b090900020302030100080a0c0b0a010505030300090c0e0b0d0a0b09000204;
    encBuf[4049] = 256'h05020302010109090c0b0c0b0b0b0a090800030604020202000008090b0d0b0c;
    encBuf[4050] = 256'h090a08080800010202040201000909090b0c0c0b0b080008000a0a0a0a080102;
    encBuf[4051] = 256'h04050303020c0f0f0c0a0a0800020304040302000a0d0d0b0b09080101020201;
    encBuf[4052] = 256'h0108090b0a08000303000b0e0c0a0a0a0a0a0902060303000c0d0c0b0c0b0b0a;
    encBuf[4053] = 256'h0004060404030201080a0c0e0c0b0b0a09000203040503030302000a0d0b0c0b;
    encBuf[4054] = 256'h0a0908000101000a0b0d0a0804050504020202080a0d0c0c0b0a090001010304;
    encBuf[4055] = 256'h02030202010809090a0b0c0b0c0b0a0a090908010405050302010009090b0a0a;
    encBuf[4056] = 256'h0a09090908080a0b0c0b0a010307030503030301080c0e0b0c0a090001030603;
    encBuf[4057] = 256'h0401080b0e0b0b0a0902030703030300090b0d0b0b0a09000202040302020009;
    encBuf[4058] = 256'h0a0909080101020300080d0e0c0b0a00040604030200090c0c0c0b0a08010405;
    encBuf[4059] = 256'h0304020108090b0c0c0b0a09080003040403030200080b0d0b0b090103060402;
    encBuf[4060] = 256'h02000a0c0d0c0b0b080004050403030101090b0d0c0b0b090801030404020101;
    encBuf[4061] = 256'h0009080808000008090c0c0c0a0a0901030504040102000000080909090b0c0c;
    encBuf[4062] = 256'h0b0b0b0a0801040504040403030302080a0f0c0b0c0b09080204040304020008;
    encBuf[4063] = 256'h090b0b0b0a08010204020200080c0b0c0b0a0002060404030201080a0d0b0c0a;
    encBuf[4064] = 256'h09000204030201080b0d0b0b0902050504030202080b0c0d0b0a0a0801020304;
    encBuf[4065] = 256'h02010109080908010204040200080b0e0c0a0b09000203040303020100080808;
    encBuf[4066] = 256'h0a090a0a000105040302080c0f0c0c0b0a0002060503040201080a0d0b0b0b09;
    encBuf[4067] = 256'h010204030301080a0b0c0b0a0002060403030301090a0d0c0b0b090800020302;
    encBuf[4068] = 256'h0108090a0803070603050200080a0d0c0b0c0909010203040303010108090808;
    encBuf[4069] = 256'h080000090b0e0d0c0b0a080004050403030201080b0d0b0c0b09090002020403;
    encBuf[4070] = 256'h04020100090b0d0b0c0908020405030303000a0e0c0b0b0a0802050304020109;
    encBuf[4071] = 256'h0a0c0b0b090102050304020000090b0d0b0b0a090002050304030101080a0c0c;
    encBuf[4072] = 256'h0b0b0a08010304040302010008080a09090809080a090908000303000a0f0e0c;
    encBuf[4073] = 256'h0a09010405030402010809090a0909080a0a0b0d0a090802030504030302090b;
    encBuf[4074] = 256'h0e0c0a080204050302000a0e0c0c0a090002040503020100090c0c0b0b0a0002;
    encBuf[4075] = 256'h0304020208080a0a0a080001030201000a0c0c0b0b0908020203080d0d0b0b00;
    encBuf[4076] = 256'h04070403030100090d0c0c0b0b0a080001030403030200080a0c0b0a09000101;
    encBuf[4077] = 256'h010108000808090e0d0d0c0b0a0a00040505020300090b0d0d0b0a0a09000103;
    encBuf[4078] = 256'h050303030108090a0c0b0b0a080008080c0d0c0b0a090104040200080b0c0c0a;
    encBuf[4079] = 256'h08020505030301000a0e0c0c0b0a09000203030101080000020203080b0f0f0b;
    encBuf[4080] = 256'h0b0a090102050303020108090a0b0b0b0b090a0b0c0e0b0a0a01040404020208;
    encBuf[4081] = 256'h080c0b0c0a0a080204030401090a0d0c0c0a0908010304030302090c0d0c0b0a;
    encBuf[4082] = 256'h08020406030201090c0c0d0b0a0800030404020208090b0c0a0a000103040301;
    encBuf[4083] = 256'h080a0d0c0b0a090003030403020109090b0b0b0a0a0a0a090a09030705050302;
    encBuf[4084] = 256'h01080b0c0c0b0a0800010101080a0a0c0a0908000307040403040200090b0c0c;
    encBuf[4085] = 256'h0a090800010100010000080a0c0b0a00050604030201080b0c0c0a0800020303;
    encBuf[4086] = 256'h00080a0a0802050504030302080a0f0c0a0a0801020000000901030504040304;
    encBuf[4087] = 256'h020200090d0c0c0b0a09080103070304030100090b0c0b0a0a09080204040303;
    encBuf[4088] = 256'h00000909000102030202080b0f0e0b0908030604020200000808080a0c0c0b0a;
    encBuf[4089] = 256'h0901020503030403020108080809080a0b0e0b0b0a090103070505030201080c;
    encBuf[4090] = 256'h0b0c0b0900010303040302010a0c0e0b090801040503030301080a0c0c0a0b09;
    encBuf[4091] = 256'h0800010305040200090a0c0a090800010103050503030300090b0c0c0b0c0b09;
    encBuf[4092] = 256'h0002060304010109090b0b0b0a09010503040201000809090908090003040300;
    encBuf[4093] = 256'h0c0f0b0b08030604020200090c0b0c0b09000305030201000a09080808000801;
    encBuf[4094] = 256'h020203000a0e0c0c0a090900030504040202000809090a0a0c0c0a090001090b;
    encBuf[4095] = 256'h0d0b00070604030208090b0c0b0b09000104030301090c0e0a0a080205030402;
    encBuf[4096] = 256'h08090c0b0a09000303030101080000000a0b0d0900030502090e0c0c09080205;
    encBuf[4097] = 256'h03030200080a0c0c0a090801030503040200090c0d0b0b090001030203030304;
    encBuf[4098] = 256'h0402080a0d0c0b0a0908080000020306040203020100090c0b0e0b0b0b0a0001;
    encBuf[4099] = 256'h0504040302080b0d0c0a080003040301010809090a0a0b0c0b0c0a0802040603;
    encBuf[4100] = 256'h030301000a0c0d0c0b0c0908020404030100090b0b0b090103030401080b0d0c;
    encBuf[4101] = 256'h0a0a0001030402010a0c0f0b0a0900030504020201020108090e0c0c0c0a0a09;
    encBuf[4102] = 256'h080002030504020302000108090b0b0e0c0b0c0b0a0a08010405030303010009;
    encBuf[4103] = 256'h080a0c0b0c0a0908010100090a0a090800000a09000407040200080c0b0d0b0a;
    encBuf[4104] = 256'h090801020302010a0b0b0b090908080002060302080d0e0b0c0b0a0a09080101;
    encBuf[4105] = 256'h0200090a0004060401080b0d0b090000090c0c0c0b0908080000000203040404;
    encBuf[4106] = 256'h040202090c0f0b0b0b090a0b0b0c08040604030200080909090a0b0d0c0a0900;
    encBuf[4107] = 256'h020201080a0b0c090102050502030100080a0c0c0c0d0b0a0901030602010009;
    encBuf[4108] = 256'h0000020200090d0c0b0b09090900000305030402010109090a0b0c0a0a090809;
    encBuf[4109] = 256'h090a09000201010009010707050301090a0c0b0b0b0a0a0a0901040504030303;
    encBuf[4110] = 256'h010100090d0b0e0b0a0a09000102040203040204030401000a0d0c0b0c0b0b09;
    encBuf[4111] = 256'h08030505040202010008090a0d0c0b0a0900030503030102010808090a0b0b0d;
    encBuf[4112] = 256'h0b0b0b08020505030102010104040202080b0e0c0c0b0c090901040503040201;
    encBuf[4113] = 256'h0008080a0b0b0d0a0a0a08010304030302010808000204040200080c0b0c0c0a;
    encBuf[4114] = 256'h090900030505020208090a0a080801010800080000030405030301090a0b0802;
    encBuf[4115] = 256'h070501000a0c0c0c0a0b090802070503040201080a0b0c0b0c0a090800010404;
    encBuf[4116] = 256'h0403030200080a0c0a0909090b0c0c0a0900040305030304030201090c0d0b0b;
    encBuf[4117] = 256'h0a00010303020208090a0a080405030301090a0b0b0b0a0c0a09010605040302;
    encBuf[4118] = 256'h010100080b0e0c0c0a0900030503040200000009080909090c0b0c0a09010304;
    encBuf[4119] = 256'h030200010205050402020109090c0d0b0d0a0908020404020101000809000001;
    encBuf[4120] = 256'h02020200080d0c0c0c0b0a090003060404030302010008090c0c0c0c0a0a0a08;
    encBuf[4121] = 256'h0802020504040303020100080a0b0c0c0c0a0a0a090001030504030302000809;
    encBuf[4122] = 256'h09090a090a0a0909090103030603020300090b0d0b080101000a0e0c09010706;
    encBuf[4123] = 256'h0304020008090c0c0b0c0a0a0901020404030303030200080a0c0d0c0a0a0908;
    encBuf[4124] = 256'h000203020101010002030304020000090a0b0f0e0b0c0a090801030304040403;
    encBuf[4125] = 256'h050201080b0d0c0b0b0a0a080001030404030304010108090c0b0d0b0b0b0a08;
    encBuf[4126] = 256'h0205040203010008090908090b0c0b0c090802030302000a0c0b0b0b09000307;
    encBuf[4127] = 256'h040202080d0c0d0b0a0801050304020108090a0a0a0b0c0b0d0a090801020303;
    encBuf[4128] = 256'h03020101080a0c0c0b0a080004030200090d0b0d0c0a0a0a0908020603030208;
    encBuf[4129] = 256'h0d0d0c0b0a090800020405040202000a0b0e0a0a0a0801000100080a09090901;
    encBuf[4130] = 256'h03030301080b0f0c0b0b0b0801030301090b0c0b010407030201080b0c0c0c0c;
    encBuf[4131] = 256'h0b0d0b0b090803070304020108080a0a0b0b0b0c0b0a0a090900020205050503;
    encBuf[4132] = 256'h0302000a0d0c0c0a0a0a080909090001040503020109090b0a09090808080101;
    encBuf[4133] = 256'h0302000b0f0d0b0b0a0b090a0a080802040305040200000a0c0c0b0a09080102;
    encBuf[4134] = 256'h030304010a0f0d0b0b0a01030303000b0c0c0a090808090a0a0a010206040100;
    encBuf[4135] = 256'h00090908090000010206010a0f0f0f0a0a09010305030301090a0b0c0a080101;
    encBuf[4136] = 256'h0101080a0c0c0b0b0a080104060403030200080b0c0c0b0c0b0a0a0901020403;
    encBuf[4137] = 256'h03030109090a0a08030504030100090d0c0c0b0a0a0a0103040603020000090b;
    encBuf[4138] = 256'h0c0d0a0b0a0802030603020008090b090801030404030302080d0e0c0b0b0900;
    encBuf[4139] = 256'h0204030201000000020203000a0d0d0b0a0002050302010809090908080a0b0a;
    encBuf[4140] = 256'h09050704030200090a0b09090a0c0c0c0a080104050303020000020205030200;
    encBuf[4141] = 256'h0a0d0b0a0a080808000201040301090c0f0a0a08020503050203020100080909;
    encBuf[4142] = 256'h08010506030302090d0d0c0b0a0a080102050405030201090b0d0c0a08000204;
    encBuf[4143] = 256'h030304010100090b0c0c0b0b0900010304030201000103040301000c0d0b0a08;
    encBuf[4144] = 256'h0002010000010405040301080a0a0a0002050202080b0e0b0b0a000102010001;
    encBuf[4145] = 256'h050704040200080a0a0a08080a0b0c0a010605040202000a0a0c0b0a09080101;
    encBuf[4146] = 256'h0102020402030101080001030402000a0e0a09020306020009090a09090a0c0b;
    encBuf[4147] = 256'h0c0902060504020100080808010000090c0b0a0005050301080b0b0b00020302;
    encBuf[4148] = 256'h090c0c0a08030502030304050403010a0f0c0c0a080102040201010008000100;
    encBuf[4149] = 256'h0108090b0b0d0a0b0a09080307040302000a0b0a09020301090f0c0b0b000206;
    encBuf[4150] = 256'h03040301010009090b0d0a0b0a0a090800080900010205030200090b00030605;
    encBuf[4151] = 256'h030203010102080c0e0e0b0c0b0a080102050302010809090909000800000002;
    encBuf[4152] = 256'h04040301090e0c0d0b0c0a080004040403020008090b0b0d0c0b0c0908010404;
    encBuf[4153] = 256'h0201000809080001000008090909090c0c0d0b0a080003040303020000080809;
    encBuf[4154] = 256'h0a0f0c0d0b0b080004050203010000090b0c0a0900040402080d0c0c0a090000;
    encBuf[4155] = 256'h010108010204040401080a0c0c0a0a0808020204040302080a0e0c0b0b0a0002;
    encBuf[4156] = 256'h02030008080003070303000a0b0d0a08080a0d0c0c0a08030503030201000101;
    encBuf[4157] = 256'h01090d0f0c0a0b080002030302010100000000090c0c0a08010302000c0e0c0a;
    encBuf[4158] = 256'h0800020102000203050302080e0d0b0b0a080000000001020504040100090b0c;
    encBuf[4159] = 256'h0b0a090000080909090900080a0c0c0a0004070304020108090a0c0d0b0d0a0a;
    encBuf[4160] = 256'h09000203040303030100090c0d0c0a0a0900010403020300090b0b0c0b0b0b0c;
    encBuf[4161] = 256'h0a0a000001000b0e0b090107050304020200090a0c0d0b0b0c0b0b0a08020405;
    encBuf[4162] = 256'h0403020100090a0b0d0b0c0a0a0801040503030301000a0c0c0b0d0b0a090801;
    encBuf[4163] = 256'h02050302020100080a090a0808010001000a0b0d0e0b0b0b0902040503030301;
    encBuf[4164] = 256'h0808090b0d0b0b0a080205040200080c0b0b0b090001030703040201090a0c0a;
    encBuf[4165] = 256'h080800000a0a080105050302080c0b0c0a09000103030404040303010a0d0d0c;
    encBuf[4166] = 256'h0a080003040402010100000a0a0e0c0b0b0a00030603040302020108090b0c0b;
    encBuf[4167] = 256'h0b0b090a080002050504020108090b0a0a0801040403040208090c0c0b0b0801;
    encBuf[4168] = 256'h030703040201080b0e0b0b0800030503020101080009090a0a08000203050108;
    encBuf[4169] = 256'h0c0e0c0b0900030504030402010100090a0c0c0b0c0a0a000003050304030201;
    encBuf[4170] = 256'h0808090b0b0b0a0a0800010100080801060604030200090a0b0b0b0d0c0a0a09;
    encBuf[4171] = 256'h0205050403020200080a0a0c0a0a0b0b0c0b0800040403030201010102030402;
    encBuf[4172] = 256'h0201090c0d0d0c0a0b09090809080004070404030100090b0d0b0a0b09000104;
    encBuf[4173] = 256'h0403030200090a0b0c0a0a090a0a0b0b0b09030705030403010100000101000a;
    encBuf[4174] = 256'h0f0e0c0a0b0900010204040203020200080b0c0c0b0b09000203030302080809;
    encBuf[4175] = 256'h0a0b0c0b0d0a090104050303010000090008090b0e0b0901040403000a0c0c0c;
    encBuf[4176] = 256'h0a0a090800020604040304020208090c0e0c0a0b08080203040303020100090b;
    encBuf[4177] = 256'h0b0c0b0a080001030302020008090800030403010b0f0d0b0a0103040301080a;
    encBuf[4178] = 256'h0800030403010002060402080f0e0c0a09010305030101080908080000000909;
    encBuf[4179] = 256'h0909010201080c0d0d0a08010404040202010000090b0d0c0c0a080204040402;
    encBuf[4180] = 256'h020000080a0c0d0b0c0a09000204050304020208090b0d0b0a09080001030302;
    encBuf[4181] = 256'h030008080a090a090900010506030302080a0c0d0a0b09080101040304030201;
    encBuf[4182] = 256'h000a0f0b0c0a0802040403020100090a0d0c0b0a090205030402080a0c0b0b09;
    encBuf[4183] = 256'h0003030403020008090a0a0b0c0d0b0b080205040200090a09010303000c0e0b;
    encBuf[4184] = 256'h0b0800080a0b0c09030704030401000a0b0d0c0a0a0808000800010305030300;
    encBuf[4185] = 256'h0a0c0c0a0a09090800040503020a0d0d0b0b08010102010103040401000b0e0c;
    encBuf[4186] = 256'h0a0a080003030200080a0c0a0b090a0b0a080207060201080b0c0b0900010000;
    encBuf[4187] = 256'h0a0c0908000100090a00030502000c0e0a0a080000080b0b0a0a010306030300;
    encBuf[4188] = 256'h0a0e0d0a09080201010809000202080f0f0c0b0908010102020305040201080a;
    encBuf[4189] = 256'h0d0b0a0b0b0c0b0c0a0901030706030201000a0c0c0a0a090a0a0a0802060403;
    encBuf[4190] = 256'h02010a0a0c0a0908090808010104030302080b0c0c0b0b0b0b09090909080107;
    encBuf[4191] = 256'h05040301000a0d0a0a0801030201080b0d0c0c0b09080204030403020201090c;
    encBuf[4192] = 256'h0e0c0b09080103030203010100080a0c0d0a0a0800010203030101090c0e0c0a;
    encBuf[4193] = 256'h0a0002040403030200090b0f0c0a0b090802030603030301080a0c0b0c0b0b0b;
    encBuf[4194] = 256'h0b0902050504020208090b0a0a0a09090a09000307040302000a0c0b0c090000;
    encBuf[4195] = 256'h010009090902050403080b0e0b0801030401000b0a0a0909090a090102050301;
    encBuf[4196] = 256'h0000010403000a09080206080f0e0c0b090104040200000a0a09080004040403;
    encBuf[4197] = 256'h00090d0d0c0a09000103030404030201080d0c0c0b0a08000103040304030100;
    encBuf[4198] = 256'h0a0b0d0a0a08000103040301000c0c0c0a09000204040202010008080a08090a;
    encBuf[4199] = 256'h0b0c0c0a080205030201000104050302000a0d0c0a080001030108090a0a0205;
    encBuf[4200] = 256'h050302080b0c0a01030503020000010102080e0c0c0a00030603030108080a09;
    encBuf[4201] = 256'h0800020200080b0e0a08020604020109090801050403020009090a0a0c0b0c0b;
    encBuf[4202] = 256'h0002060302000000010504030301000a0d0c0c0b0901040504010008090a0800;
    encBuf[4203] = 256'h010203030301090d0e0c0b0b08010305040403030201080c0c0c0a0a08010202;
    encBuf[4204] = 256'h0303040101090b0c0c0a09000204040303020108080a090a0a0b0e0c0b0a0803;
    encBuf[4205] = 256'h06050402020101090b0b0d0a0b0900010203020102030304030200080a090a0a;
    encBuf[4206] = 256'h0a0c0c0a090207060304020100080b0d0c0c0a09080304040302010108080001;
    encBuf[4207] = 256'h0001080c0e0c0b0a08030704020208090a0a0b09090000010103030204020102;
    encBuf[4208] = 256'h020002000a080a0b0d0e0d0b0b09020504030303030403010a0f0d0a0a000203;
    encBuf[4209] = 256'h0300090a0b0b0808090100000306040504030402080b0e0d0b0b0a0801010303;
    encBuf[4210] = 256'h0503030301080b0d0c0b0a0a090808000204030503030201090c0d0d0b0a0908;
    encBuf[4211] = 256'h000002020204020201080b0c0b09010101090d0d0b0b0a000203040202020200;
    encBuf[4212] = 256'h08090d0c0d0c0b0b0a00010204030402030201080b0f0c0c0b0a0a0000020403;
    encBuf[4213] = 256'h040302000a0e0b0c0a0900000101000008080809080004030401090e0c0c0a08;
    encBuf[4214] = 256'h000101000809090a0a0b0b0a0901070404030200080b0e0d0c0b0b0a00010303;
    encBuf[4215] = 256'h0201000101020203030402000f0e0e0b0c0a090001030503030302000a0d0d0b;
    encBuf[4216] = 256'h0b0b09080002030405030201080b0d0b0c0b0a0900000103030202020008090d;
    encBuf[4217] = 256'h0c0b0a09010101080c0e0b090803040302000a090909090d0e0c0c0a08080202;
    encBuf[4218] = 256'h02030302030201080a0f0d0c0b0c0a08010306030200080a0b0b0c0a0a0a0901;
    encBuf[4219] = 256'h03050402000a0d0c0b08000405030301000a0c0c0c0b0a0a0900010306030402;
    encBuf[4220] = 256'h00080a0a0a090900090a0a0900050304000a0d0c0c090001040404020201000a;
    encBuf[4221] = 256'h0d0b0d0a0b090800010305040303040201080b0d0d0c0a0a0900020304030402;
    encBuf[4222] = 256'h020008090b0c0b0b0b0a09000304030201080a0a08030704040101080b0b0c0b;
    encBuf[4223] = 256'h0b09090102030402000a0a0a080405030401080808080101090a0f0d0b0c0900;
    encBuf[4224] = 256'h03050503030300090a0d0b0c0b0b09080104050403020201090b0d0c0b0b0801;
    encBuf[4225] = 256'h040503020108090b0b0b0a0a0008020304040303030201090d0d0c0c09090103;
    encBuf[4226] = 256'h050304030101090b0d0c0b0a090002040403030301000a0d0c0b0c0a08010306;
    encBuf[4227] = 256'h0302020108090a0a0a0a0a0a0c0a0a0104070304010109090a0b0b0a09090002;
    encBuf[4228] = 256'h04040303020200090a0d0b0c09080002020204030305030200090c0e0c0b0c0a;
    encBuf[4229] = 256'h0801030703040302000a0b0e0c0a0a0802030402020108080908080008080b0c;
    encBuf[4230] = 256'h0c0b08000403040201010008080a0c0d0b0a08030606030201080a0d0c0a0b09;
    encBuf[4231] = 256'h0802030503030301080b0d0c0b0a080103030401010800090809090808020203;
    encBuf[4232] = 256'h0201090a0d0c0c0b0a08040503000b0e0b080307050201080a0c0a0a08000001;
    encBuf[4233] = 256'h0808090900040604030201090b0d0c0c0c0a0a08020704030201090a0c0b0a08;
    encBuf[4234] = 256'h09000808010205040301000a0d0b0b090002030200090b0c090106040401000a;
    encBuf[4235] = 256'h0b0e0a0a090002030503030100090b0c0d0b0a0a000204030201000808020304;
    encBuf[4236] = 256'h02090e0c0c0b090802020302030202030302080d0f0b0c090001020200090a08;
    encBuf[4237] = 256'h0105050202080b0c0d0a0a0800030304020009090a090800080002060403010b;
    encBuf[4238] = 256'h0f0d0b0b0801040304020100080a0a0c0b0a0a000205040202080b0d0b0a0003;
    encBuf[4239] = 256'h0502000a0d0a0a000102010808080204040200090b0b090908090c0d0a0a0801;
    encBuf[4240] = 256'h04040301000908010204020a0f0e0b0b0a0001030604030303080b0f0d0a0a00;
    encBuf[4241] = 256'h02020302000809000000080b0e0b0a0804040402000a0c0b0a08000100080900;
    encBuf[4242] = 256'h0207030400090b0d0a09000201000a0c0b0a000505030401000a0b0c0c0b0909;
    encBuf[4243] = 256'h01020303040101080808000001090b0e0c0b0908020304020108090b0d0b0900;
    encBuf[4244] = 256'h0206030302000c0d0d0a0a0801040403010108090909090a0b0d0c0b0a090001;
    encBuf[4245] = 256'h0404020301010103050301090e0d0c0b0a080001020102030303040200090c0d;
    encBuf[4246] = 256'h0c0b0a09010203040200090a0c0a090103060401000a0c0b0b0a000000090d0c;
    encBuf[4247] = 256'h0a00050605030200090c0c0b0c0a08080001030503020200090b0a090002010a;
    encBuf[4248] = 256'h0f0d0b0a000204030401010008090a0a0b0a0a09080808080801020405030301;
    encBuf[4249] = 256'h080c0c0a0802070301080b0f0c0a090801020305030401080b0e0c0a08000403;
    encBuf[4250] = 256'h0301090c0c0a090104040200000a0a0b0a0a09090103040302090c0c0a000306;
    encBuf[4251] = 256'h0302000a0c0c0b0a08010203030203020302080b0f0d0b0a0a08010303050304;
    encBuf[4252] = 256'h0201090d0d0b0b080204030300090a0a09000200090c0d0c0901030704030100;
    encBuf[4253] = 256'h090c0d0b0a0a090001030504030301010a0b0d0c0a0a08000102020201010102;
    encBuf[4254] = 256'h0202000c0d0c0c0a0908020307030402000a0c0d0c0a0901020404030101090a;
    encBuf[4255] = 256'h0a0c0a0909080808010103040305020200080c0c0d0b0a090003040303010101;
    encBuf[4256] = 256'h010202000a0f0c0b0b0a0001040302030101080a0a0b0a090003040403010009;
    encBuf[4257] = 256'h00000201090e0e0b0901050402000a0d0a090204040201090a0a0a0808080b0d;
    encBuf[4258] = 256'h0a09030605030100090a090802010108090a080204020b0f0e0a090104050202;
    encBuf[4259] = 256'h08090b0a090103030300090e0c0c0b0b0802070503040100090c0b0c0a0a0808;
    encBuf[4260] = 256'h010102050404020208090c0b0b0a0808000808000104040304010009090a0b0c;
    encBuf[4261] = 256'h0c0b0a08030603040200080b0c0b0c0a09010305040302020100090b0e0b0c0a;
    encBuf[4262] = 256'h0a080002040403030301080a0b0d0b0a0a090909080102050303030404040302;
    encBuf[4263] = 256'h090d0d0d0a090801020302000108000009080a08000405040302090b0f0b0c0a;
    encBuf[4264] = 256'h0908010305030402010108090a0c0a0c0a0a090a0a0a00020705030302010809;
    encBuf[4265] = 256'h0a0a0c0c0c0a09000404030200080a0a0a0a090908080206050202000b0d0c0a;
    encBuf[4266] = 256'h090001030200080908030602010a0e0c0a090204030108090b0a00020401000a;
    encBuf[4267] = 256'h0908010202090f0d0b090206040401080b0c0b0a090102020301010101090a0e;
    encBuf[4268] = 256'h0c0a0a08010202010201010100080800040602010b0f0c0b090003060303010a;
    encBuf[4269] = 256'h0b0e0b090800000008000206040400080c0d0a09000201010809080002040300;
    encBuf[4270] = 256'h090b0c0c0a0908010204020201000000090c0f0b0c09010404030108090a0909;
    encBuf[4271] = 256'h09090a0b0b090900000800000405040301000a0d0d0c0c0b0908020603040100;
    encBuf[4272] = 256'h0809090908080a0d0c0c0a08020505020208090b0b0b08000001090c0b0c0a08;
    encBuf[4273] = 256'h02040502020008090a09090b0d0d0b0a0a000101030604050302010b0e0c0b0a;
    encBuf[4274] = 256'h0801030301000a09090104060303000b0f0c0b0b0a0802030504020208090a0c;
    encBuf[4275] = 256'h0a09080808090a0a09030705030300090b0d0b0b090000020303030302010a0d;
    encBuf[4276] = 256'h0d0b0b0a08010102010303040402000a0d0d0a0b0a0808000008080206060403;
    encBuf[4277] = 256'h02000a0d0c0b0b0908000202040305020200080a0c0b0b0b0908010101080a0b;
    encBuf[4278] = 256'h0b080606040302080a0e0b0b0b0900020403040200080b0b0b0a080003040403;
    encBuf[4279] = 256'h040101090a0c0c0b0b0b0b0b09020707030302000a0c0c0a0a08000000000909;
    encBuf[4280] = 256'h0901020604030200090c0c0b09080103030201080b0c0b0a0805050503020009;
    encBuf[4281] = 256'h0b0b0b0b0908090a0b0b0a00050705030402000a0c0d0b0b0b09000305040302;
    encBuf[4282] = 256'h0200090b0b0c0a09000103030302010008090000010108090c0d0c0b0a010506;
    encBuf[4283] = 256'h04030200090c0d0a0b0a080801020403040202010000080a0a0e0c0b0b0a0004;
    encBuf[4284] = 256'h060304020008080a080908080b0c0b0b08050604030208090c0b0c0909080101;
    encBuf[4285] = 256'h0102020304020201080a0e0c0c0b0a0002060403030108090c0b0a0908010201;
    encBuf[4286] = 256'h080909000505040201000a0a0c0b0a0b0a0808020204040302030301090c0d0c;
    encBuf[4287] = 256'h0a0b090901030704040200080b0b0b0a01020303010808090001010304030503;
    encBuf[4288] = 256'h03010a0d0d0c0b0909010103020208090800020405020301010000090a0f0d0d;
    encBuf[4289] = 256'h0c0a0901040703030201090a0b0b09080808080a0a080105040303000a0c0c0a;
    encBuf[4290] = 256'h0003060401090a0c0b090801000009090001050403030302040303020b0f0f0d;
    encBuf[4291] = 256'h0a0908020404030200080909090808090c0c0c0b09010307020301080a0b0c0a;
    encBuf[4292] = 256'h0808010202010200010100080a0f0b0c0a0900020504030402020200090c0c0d;
    encBuf[4293] = 256'h0c0a0a08000104030403020200080b0e0c0b0b0a090102040303020100010100;
    encBuf[4294] = 256'h080b0e0c0b0b0908010203040403030200080b0e0b0c0b0b0908020404030101;
    encBuf[4295] = 256'h00090809090c0d0d0b0a09010306030201000a0b0c0b0b0a0900010403040303;
    encBuf[4296] = 256'h01000a0d0c0b090900010008090901050402090c0d0c0a090101020301000809;
    encBuf[4297] = 256'h0a0c0c0b0b080000080a0a090107050201090d0c0b0b09010307040303010a0c;
    encBuf[4298] = 256'h0d0b0b0a09000102030404040201080b0d0c0b0b0a0800030404030100090c0c;
    encBuf[4299] = 256'h0b0a090002030403010008090a0a0a0b0a0c0b0c0a0801070404030302080a0d;
    encBuf[4300] = 256'h0d0c0b0a0a00020304020201000008080a0a0d0b0b0a00010200090901050704;
    encBuf[4301] = 256'h0301090d0c0c0a000104030401000a0c0b0a0908000200010801010304020208;
    encBuf[4302] = 256'h0a0b0e0b0c0b0b0b0b09000206050404020100080a0a0c0b0c0b0a0900040503;
    encBuf[4303] = 256'h040200080a0a0b0b09080100000909080207060301090b0f0b0a090002030403;
    encBuf[4304] = 256'h02030200080c0e0c0b0a090102040303020201010808090c0d0c0c0a09000303;
    encBuf[4305] = 256'h0502010008010001080a0d0d0b0a080304040201080a0b0b0a09000102040203;
    encBuf[4306] = 256'h020201000b0d0b0b0a010304020a0c0d0a010605030302090c0c0b0a09080202;
    encBuf[4307] = 256'h0108090b0b0b090204060404030201090c0d0c0b0b0908020405020301080a0a;
    encBuf[4308] = 256'h0a08000301080b0e0a080204040108090b0c09080204040201080b0c0c090800;
    encBuf[4309] = 256'h01020201010200090c0c0b0a02030603010102030402000c0f0c0c0a09080204;
    encBuf[4310] = 256'h0503020201080a0c0c0c0a0a09010103050203020101080a0d0e0b0a09010304;
    encBuf[4311] = 256'h030303020101080b0e0c0c0a0a080102040403040101080a0a0b0c0a0b090900;
    encBuf[4312] = 256'h03040302010202060403000a0e0d0a0a08010102020201020200080c0c0b0b08;
    encBuf[4313] = 256'h030405030100080a0a090a090a0c0b0b0804070404020208080a0a090909090b;
    encBuf[4314] = 256'h0c0b0c09010306050304020200090d0c0c0a0a080204030401010809090a0b0b;
    encBuf[4315] = 256'h0b0b08020706030301000a0c0c0c0b0908000303050303020100090c0c0c0b0a;
    encBuf[4316] = 256'h09000204030402000009090a0a0a0808010204040302080b0c0c090802020100;
    encBuf[4317] = 256'h0a0b0a00050604040101090c0c0b0b0a08000204030304030301090d0d0a0a08;
    encBuf[4318] = 256'h0203030302090b0e0c0c0908010306030201000a0a0a0a0a0908080103030100;
    encBuf[4319] = 256'h0c0d0b0b080307040304020100090c0d0c0b0b08000305030202000008080809;
    encBuf[4320] = 256'h0b0c0c0b0c09080003050403030300090b0e0b0c0a0808010101010103070503;
    encBuf[4321] = 256'h03000b0f0c0b0a0900020402020201010000090b0d0b0a09010101000a0a0802;
    encBuf[4322] = 256'h06040302000a0c0b0a08000103010100090009090c0f0c0c0a08030504030108;
    encBuf[4323] = 256'h090a090808090c0d0d0a0a080204030503030200080a0d0b0b0c0a0909080101;
    encBuf[4324] = 256'h0303040304030302000a0d0e0c0a0b09000204040201000a0b0b0a0900010303;
    encBuf[4325] = 256'h050202000a0d0d0c0c0a08000404030401000a0b0b0b0b0a0a0b090105060303;
    encBuf[4326] = 256'h01090c0c0b0a08010303030101080909090b0c0c0c0b0c0a0800050504030303;
    encBuf[4327] = 256'h080a0d0e0c0a0a08000303050202010008090a0b0d0b0b0b0a09010307040302;
    encBuf[4328] = 256'h01000a0c0b0c0a090900000100010304040302000a0f0c0b0b0b080103050404;
    encBuf[4329] = 256'h020101080b0d0c0c0a0a0001030503030200080b0b0d0b0c0a09000203050302;
    encBuf[4330] = 256'h0008090a0b090900080a0b0c0a08020604020100090a0a090a0b0a0b0a090104;
    encBuf[4331] = 256'h0603040201080a0c0d0b0c0a0a08010307030301000a0c0b0c0a0a0001030305;
    encBuf[4332] = 256'h0101080a09090800010108090b0c0b0b0a0103060301080b0b0805060303090d;
    encBuf[4333] = 256'h0e0b0c090002030403030008090a090008090d0e0c0b09000404040202000908;
    encBuf[4334] = 256'h0a090908090a0c0c0d0a08020405030100090a09090101020100090b0d0c0c0a;
    encBuf[4335] = 256'h0a0001040503040201000a0c0c0b0900020302080b0d0c090102050302030001;
    encBuf[4336] = 256'h00090a0b0f0c0a0b09010304030108090a000405040201090b0d0b0b0b0a0a09;
    encBuf[4337] = 256'h080204050504030201080a0d0b0b0b0a0808000203040403020202030403010a;
    encBuf[4338] = 256'h0f0f0b0b0a08010204040202020008090a0b0c0a0b0909010205030302080a0c;
    encBuf[4339] = 256'h090803050402000a0e0b0b0a08020204020202030203080c0e0c0b0900040303;
    encBuf[4340] = 256'h01080c0b0a0802030301090d0a000406040301080a0c0a0a090a0a0b0d090004;
    encBuf[4341] = 256'h0604030301000a0c0b0a0b0a0a0a0a000207040402010109090a0a0b0a0c0a09;
    encBuf[4342] = 256'h09000204050403020108090b0c0b0a0a0800030703030300090d0c0b0a090802;
    encBuf[4343] = 256'h040404030101080a0b0b0b0b0a09090104060403020200080a0d0c0a0b090802;
    encBuf[4344] = 256'h05030402020000090a0a0a0b090800020404030201000a0b0a0002060303010a;
    encBuf[4345] = 256'h0d0d0b0b00020604030201080a0909000000080800020703000b0f0d09080204;
    encBuf[4346] = 256'h050303010108090c0c0c0b0a080104030403030201090c0d0c0b0a0801030403;
    encBuf[4347] = 256'h030402010100090b0f0b0c0a0a0002050403010109090909000809090b0a0802;
    encBuf[4348] = 256'h0403000b0d0b0805050403010a0c0c0b0801040303000a0d0b0a090801010102;
    encBuf[4349] = 256'h040604040202080b0e0c0c0a09080103040402020108090a0c0b0a0a09080001;
    encBuf[4350] = 256'h02030404020208090b0d0a09000102030201080b0f0c0b09000206030300080b;
    encBuf[4351] = 256'h0c0a00020502000a0d0c0b090103040201080a0900010301090a0c0a08080a0d;
    encBuf[4352] = 256'h0d0c090104040302000a0a0a09000201090d0e0c0a0800030503010108090001;
    encBuf[4353] = 256'h0101090d0e0c0a0b0800030304030101080909080908090c0c0d0b0c09080203;
    encBuf[4354] = 256'h050301000808000102000a0e0d0b0a0800000808090803060304010100000009;
    encBuf[4355] = 256'h0d0d0d0b0b0b090801030605030201080a0c0b0c0a0a09080103040302010809;
    encBuf[4356] = 256'h0a090b0b0b0a00030502080a0b0b080204000a0f0e0b0b09000404040202080a;
    encBuf[4357] = 256'h0c0c0a0a0909000001020108090a0802070502010a0c0d0b0a08000303030201;
    encBuf[4358] = 256'h08090c0b0d0a0a090001040302030208090d0c0c0c0b0d0a0a08020604030301;
    encBuf[4359] = 256'h080a0c0c0b0c0a0908000204030402010008090a0b0a090b0b0d0b0a08000203;
    encBuf[4360] = 256'h0503040402010a0e0c0c0a0908000102030201000a0d0d0a0a08020304030201;
    encBuf[4361] = 256'h0100000a0c0f0d0b0c0a0001050403030200090a0c0b0b0b0c0b0a0a08020505;
    encBuf[4362] = 256'h03040100090a0b0a0b0b0a0a09080104040200090b0b0805050303010a0b0d0a;
    encBuf[4363] = 256'h090908000101000a0e0b0b000505040208090a0a0a0800080a0c0d0c0b0b0a01;
    encBuf[4364] = 256'h060504030100090a0b0b0a0a090a0b0b0a0104070504020108090a0b0b0b0908;
    encBuf[4365] = 256'h080808090801030704030200080b0c0b0b090008080b0b0d0900040504020202;
    encBuf[4366] = 256'h0201080a0d0c0c0b0900010305030302000000080001080a0f0e0a0a00020403;
    encBuf[4367] = 256'h0200090a09080001010100090a0c0b0a080104030304020203000a0a0a080706;
    encBuf[4368] = 256'h040304020100090c0d0d0a08000404030200090a0a00010201080c0d0c0b0900;
    encBuf[4369] = 256'h03050303020009090800010101080a0a0b0a00010205070505030302090a0c0b;
    encBuf[4370] = 256'h090800000a0a0a00060604030201090c0c0c0b09080102040303040101080a0a;
    encBuf[4371] = 256'h0c0b0b0a0802060502020108090800020302000a0c0c0a090802040302020103;
    encBuf[4372] = 256'h06040401080c0e0c0a090803040303020808090908090a0b0d0a080206040302;
    encBuf[4373] = 256'h020100000a0a0d0b0b090803070403040108090b0c0b09000102030200090a0c;
    encBuf[4374] = 256'h090103060301000a0d0b0b0a08020305030302010000000104040302080b0e0b;
    encBuf[4375] = 256'h0c0a000206050203010809090a080a0b0c0d0a0a08000202030604030401080a;
    encBuf[4376] = 256'h0e0c0c0a0800030403030100080908080800090a0b0b0a000507040202010a0b;
    encBuf[4377] = 256'h0e0b0b090802030503020008090c0c0b0c0a090102030302010000030201000a;
    encBuf[4378] = 256'h0e0c0c0b0b08020605020200090a09090101020100090b0d0d0b0c0a09000205;
    encBuf[4379] = 256'h030401000a0c0b0c090a0a0a0b0a08010605040303000a0c0c0c0a0908020304;
    encBuf[4380] = 256'h03020100090a0a0b0d0b0a0901020303010a0b0b0803010c0f0f0d0a08000304;
    encBuf[4381] = 256'h0302080a0d0b0b09080202020109090902040502000b0d0b0b08020203010008;
    encBuf[4382] = 256'h0909090a0c0b0c0b0b0b08020503000b0f0e0b0908000001080a0b0b0b080306;
    encBuf[4383] = 256'h03010a0e0c0a0802030301080a0a0900020303090d0c0c0a000203080d0e0b0b;
    encBuf[4384] = 256'h080101080b0d0b0a09080100080b0f0c0c090802030401080b0a0b0908090809;
    encBuf[4385] = 256'h080405030300090c0b0a090800080d0e0b0c0a0801030302080b0f0d0c0b0c09;
    encBuf[4386] = 256'h0802040302010a0c0b0c0a0909080808010505040200080c0b0c090900000000;
    encBuf[4387] = 256'h010003040401000b0e0c0b09080001010009090a09000102010a0e0d0c0a0909;
    encBuf[4388] = 256'h01020203040101080d0c0b0908010202020101020800010a08080d0b0b0b0902;
    encBuf[4389] = 256'h08000a0e0005080a0f0e0a09000202000b0c0c0a000101010008000003050402;
    encBuf[4390] = 256'h010c0e0b0b0803070303010809090800080a0a0f0b09080205040301080b0c0b;
    encBuf[4391] = 256'h09080000080a0b09090106030403010a0c0d0900010303010001000305010202;
    encBuf[4392] = 256'h000a090c0a0900060401010100040402000c0f0b0a080204030201090a080908;
    encBuf[4393] = 256'h00080000090102020604010301090002020502090a0a00070705020008090a0a;
    encBuf[4394] = 256'h09000103030203000801020101080f0b0a0a01050304020101000a0900010604;
    encBuf[4395] = 256'h0302000800010307030101090a0a010607030301090d0a0902040402000a0b09;
    encBuf[4396] = 256'h080204030300090b0b0b08040504020200000000080a0c0a0007050402010009;
    encBuf[4397] = 256'h0a0a090001040302030304030202080a0c0a0802050401010001020304020108;
    encBuf[4398] = 256'h01010104000b0c0908050603040201010101030401080c0e0a09030705030208;
    encBuf[4399] = 256'h09090a0801020100090a00020507020200090c0b0a0803030402000800010102;
    encBuf[4400] = 256'h000b0b0b090505040403010100090808090a0a0b00050704030202000908090d;
    encBuf[4401] = 256'h0b0b0b00050504030200090b0b0b0b08010203040203020202080a0808010501;
    encBuf[4402] = 256'h0c0b0f0c08000404040201010808090b090b0d0a09000404040301080a0a0901;
    encBuf[4403] = 256'h0302080f0d0b0a0804050303000a0c0b0b08010201080d0a090004050302080a;
    encBuf[4404] = 256'h0b0d0a09000102010001080801020202080e0b0d0c0909090002010401010009;
    encBuf[4405] = 256'h0b0b0d0d0a0b0b0a080106030303000c0c0d0b09090102030100090b0a0a0b08;
    encBuf[4406] = 256'h0a0c090a0c080a0a020301030a0f0f0b0b0b0c0a0900010402080009090a0d0e;
    encBuf[4407] = 256'h0c0c0b09000103030202080b0d0c0c0a0909090b090104040402080a0d0d0a0b;
    encBuf[4408] = 256'h09090001000100010100000a0f0b0d0b0a0a0a0a090003050401000b0c0c0c0a;
    encBuf[4409] = 256'h0a0a0908000103040302080c0f0b0c0a08000102000008090801000a0e0e0c0a;
    encBuf[4410] = 256'h0a0802030401000a0d0b0a0a08080008090b0b08010302000a0e0b0b0e0c0b0c;
    encBuf[4411] = 256'h090003050301080a0c0b0a0a0a0a0a090a0002050403000a0e0c0c0a0a0a0808;
    encBuf[4412] = 256'h00000100010800010a0f0c0d0b0a0900020303050201000b0e0b0b0a08080000;
    encBuf[4413] = 256'h080105030403080b0e0d0c0a0908020302020a0a09090801080a0b0e0a0a090a;
    encBuf[4414] = 256'h08000307040302090b0b0d0a090909000800020104050303000c0f0b0c090800;
    encBuf[4415] = 256'h020201010201040300090c0f0c0a090004030303000809090a090b0c0c0c0a00;
    encBuf[4416] = 256'h0003060303020108090c0b0d0b0908020504020201010000090a0a0d0b090901;
    encBuf[4417] = 256'h05040302080a0a0a080109090b0f0c09000307030202000b0a0c090800010102;
    encBuf[4418] = 256'h04060302030100090a0c0c0d0a080003060202020008090c0b0b0a0808080002;
    encBuf[4419] = 256'h040704020201090a0a0a090808000304050403040201080b0e0b0b0908020203;
    encBuf[4420] = 256'h0503030300080b0e0b0a09000302030202040604040200080b0c0c0909010204;
    encBuf[4421] = 256'h02020202020202080c0d0d0a0a0000020402040302020208080b0d0b0b080306;
    encBuf[4422] = 256'h04040202010000090a0c0b0c0a08010205030302020101090b0f0c0b09080305;
    encBuf[4423] = 256'h050302020100090b0b0a09010303040202040305030108090c0d0c0a0a080104;
    encBuf[4424] = 256'h040202000808080908080a0a0902070604030300090a0b0a0801020200010102;
    encBuf[4425] = 256'h07040202090c0d0c0a09000202030304020101080a0a0a0b0a0a080407050303;
    encBuf[4426] = 256'h02010008090b0c0b0c0a0901040403020300080a0a0c0c0b0c09010307030302;
    encBuf[4427] = 256'h0100000808090b0c0b0a0803060405020201080b0a0c0c0a0b0a080102040303;
    encBuf[4428] = 256'h04030301090f0c0a0a080102030504040200080b0b0a0908080a0a0104050401;
    encBuf[4429] = 256'h000a0b0e0a0a090808010101020305030400090b0e0b0a080003040404020202;
    encBuf[4430] = 256'h080a0b0d0c0b0b0a080102040302040101090c0d0c0c0a090801030404030202;
    encBuf[4431] = 256'h00080a0d0c0c0a0a080304030201010101090b0f0f0a09080001010203020301;
    encBuf[4432] = 256'h080a0d0d0a0b090901020603030300090a0b0b0d0c0b0b0a0802050304020808;
    encBuf[4433] = 256'h0b0b0c0b0b0a0a0900020405040303000a0b0c0a0a0a0b0c0b08030704020009;
    encBuf[4434] = 256'h0a0a0b0b0c0d0b0a0802020302010100080b0c0d0b0c0a090002040503030201;
    encBuf[4435] = 256'h080c0e0b0b0a080800080801040401090e0c0b0a090808000003030302000809;
    encBuf[4436] = 256'h0a0e0d0b0a0104030208090a0103030b0f0f0c0908000008080001020100090b;
    encBuf[4437] = 256'h0d0c0b0c090801040503020200080a0b0b0b0d0b0b0c0a0004040301080a0b0b;
    encBuf[4438] = 256'h0b0e0d0b0c090102030302020101090a0c0b090a090b08050705010009090900;
    encBuf[4439] = 256'h000a0f0b0b09010202090a0a000302090f0c0b08010001080003050502000808;
    encBuf[4440] = 256'h08090008090b0c0a09030703000a0d0c0a0101000b0e0b0a0802030108090002;
    encBuf[4441] = 256'h0301090900040501000800050501090b0b090402080c0c0a0000000d0d0b0801;
    encBuf[4442] = 256'h01080c0b0a01060302080800030303080c0d0901050403010908090002010b0f;
    encBuf[4443] = 256'h0e0a0a00010108090a000304010a0e0b09010101000902070503010009080001;
    encBuf[4444] = 256'h080b0d0a080204020008080000090d0e0c0a0a08080800020503030208090809;
    encBuf[4445] = 256'h0009090b090207060403030109090909080a0e0c0b08010303000b0d09010301;
    encBuf[4446] = 256'h0c0f0a0901030400000801050302080b0a08020501080909020503010b0d0c09;
    encBuf[4447] = 256'h080008090a0b080102010000080008000800040505040203030404030100090a;
    encBuf[4448] = 256'h0908000102000a0c0c0a090a0b0f0d0b0909000108080207050201080b090005;
    encBuf[4449] = 256'h030209090007060202090a090802010a0d0d0908030200090b080204020a0f0c;
    encBuf[4450] = 256'h090002030008080104050301000908000101080a0b0902060401000a0b080001;
    encBuf[4451] = 256'h0a0f0d0a08010302000b0b00050402080b0b01050501080900020503010a0c0a;
    encBuf[4452] = 256'h010401080c0c08020402090c0b0a010302090c0c0803040301090a0003050300;
    encBuf[4453] = 256'h0a0b00030702010a0c09010403000c0c0a000303000c0c0a000304000b0d0902;
    encBuf[4454] = 256'h0403000a0a08050402000b0b00040401080b0b000404000a0d0a000302000c0c;
    encBuf[4455] = 256'h09000402080b0c09010503080a0a09050403000b0b0a020503000c0b09030503;
    encBuf[4456] = 256'h080b0c090103010a0f0b08020303080c0b08040402080b0c08010403000a0a08;
    encBuf[4457] = 256'h020502080b0b090103010a0d0b08030500090d0b000203010a0d090205040009;
    encBuf[4458] = 256'h0b0a00040300090c0a00040301090c09080102090e0c0908020200090a0a0204;
    encBuf[4459] = 256'h02010b0f090802040301090909020403010c0e0b0a000102000a0d0902050208;
    encBuf[4460] = 256'h0c0e0b08000200090b090107040100090b080001000a0c0a0802060100080a08;
    encBuf[4461] = 256'h01000b0e0d0b09010201090c0a08040501080b0c09000402000a0b0902040200;
    encBuf[4462] = 256'h0b0a0103030c0f0c080103010c0f0a09020302090e0a09020401080c0a080304;
    encBuf[4463] = 256'h02090b0b010405010a0c0a080203000b0e0a000305000b0d0b080202010b0e0a;
    encBuf[4464] = 256'h00030501080b0a00030400090d0908030401090b09010403090d0c090001010a;
    encBuf[4465] = 256'h0c0b080204010a0c0b000403000a0e0a00030401080a0a01040301090c090002;
    encBuf[4466] = 256'h03080d0d09080202090d0c0a000303080b0f0900020301090d0900030501080a;
    encBuf[4467] = 256'h0900030400090c0a080202010a0b0a0800090c0c0b0a09090b0c0b0902030404;
    encBuf[4468] = 256'h030201090a0803060402090a090207050108090a0900080a0c0e0a0909090909;
    encBuf[4469] = 256'h00030201090c0a000201090c0a000704020201020403030201080b0b0d0b0c09;
    encBuf[4470] = 256'h0a0b0b0c080102010b0f0d080202080d0d0a08040402080808030603000a0c09;
    encBuf[4471] = 256'h020303090d0b08040502090c0b0a0103010b0e0c09020303000a0b0803060208;
    encBuf[4472] = 256'h0c0b08040502080a0b00050402090c0b090204010a0c0b08040400090c0b0002;
    encBuf[4473] = 256'h03010a0d0a020503000a0b09020602000a0c08010502000b0b09010402090d0b;
    encBuf[4474] = 256'h0a010403080b0b09030601090c0c08020402080a0a01050402090b0b00030300;
    encBuf[4475] = 256'h0d0c09020403000c0b090203010b0f0a08020401090b08010503000b0b090205;
    encBuf[4476] = 256'h02000b0b00050401080b0b080203000b0e0a080303000b0e0a000303010b0d0a;
    encBuf[4477] = 256'h01050301090a08040502000b0b08030503090c0c090203020a0d0c080203010a;
    encBuf[4478] = 256'h0e0a08030302090d0a000503020a0c0900050401090b0b00040401090d0a0002;
    encBuf[4479] = 256'h03000b0d0b000303010b0d0b010403000a0d09020502000a0b08030503080b0c;
    encBuf[4480] = 256'h08020302090d0a080203000b0e0a000201090c0b09030402080b0a0107030108;
    encBuf[4481] = 256'h0b0901040400090a08020403000c0d090802010a0c0c09010200080c0a080303;
    encBuf[4482] = 256'h010b0e0900050302080900040503000a0b090203030a0f0b080202010c0d0a08;
    encBuf[4483] = 256'h0201090f0b09010402080a0b00060402080c0a08040401080b0b000503020a0d;
    encBuf[4484] = 256'h0a080203000c0e0a000302000b0d0a010402000a0d09020403000a0c09020502;
    encBuf[4485] = 256'h000a0c08010303080c0c090103020a0d0b090203020a0e0b00020401090c0a00;
    encBuf[4486] = 256'h040401080b0a01050301090c0a010304000b0c0b000204080b0e0a000103000a;
    encBuf[4487] = 256'h0d0a010303010a0c0b0005040108090a01030501080a0b09020401090c0c0a00;
    encBuf[4488] = 256'h0302090c0d0b080102000b0c0a0104050208090908030303000a0a0804050201;
    encBuf[4489] = 256'h090a080001090e0d0b0b090000080b0a09010201090c0d090003030301020605;
    encBuf[4490] = 256'h0403010008000100080b0e0b0a000202090e0b0b0900080d0e0b09000302080c;
    encBuf[4491] = 256'h0a00060502000a0a08030602080a0b01040501090c0b080202000c0e0a080202;
    encBuf[4492] = 256'h000b0d0a010402080a0c09030502080a09000503020a0c0a010502000b0c0901;
    encBuf[4493] = 256'h03020a0e0c080102010b0e0a000303010a0d09010403010b0c09020702010a0b;
    encBuf[4494] = 256'h09010502080b0d09000401080c0b08010303090d0b09010302090b0b00060302;
    encBuf[4495] = 256'h08090a01040301080a08010201080a0a0801080d0e0b0a09080a0c0a09020100;
    encBuf[4496] = 256'h0b0d090206040100090803060401080a0900030402080a0c0a000102090e0c0a;
    encBuf[4497] = 256'h090800080b0d0908030201090a0a010603030000030704020009090003060109;
    encBuf[4498] = 256'h0d0b090103000b0f0a080202000d0d0a000204000a0b09020703000a0b090405;
    encBuf[4499] = 256'h02000b0c09030502080c0b080203020a0f0b08020301090d0a08020400090b0a;
    encBuf[4500] = 256'h01040400090a09030502010a0b08010402080c0a09000202090c0b0b09080808;
    encBuf[4501] = 256'h0a0a0a0a080105050200090802060501080a0a01060402080b0a080203000c0e;
    encBuf[4502] = 256'h0a000102090c0c0a010202090b0d090103030009080106030301090800020203;
    encBuf[4503] = 256'h00000001000a0b0c0b0c0c0d0c0c0a090808080909080800020503010a0d0a02;
    encBuf[4504] = 256'h07060201080808020402000b0c0a000403090d0d09080202090c0c0b00010308;
    encBuf[4505] = 256'h0a0b0a04060201090b090206030208090901030401090b0c090000080b0d0b0a;
    encBuf[4506] = 256'h09000102080b0f0d0908020302090c0a01070402000a0b00040502080c0a0803;
    encBuf[4507] = 256'h0402090c0c080103000b0f0a09020201090b0b08040401080b0a00050303080b;
    encBuf[4508] = 256'h0a00040503000a0a0a090101000b0c0b090003010a0f0c0a000203080c0d0a00;
    encBuf[4509] = 256'h040302090a0903070400090a09020603000a0c09000202080d0c0a010202080b;
    encBuf[4510] = 256'h0d0a000203000a0d0a01030402090a08030603020a0c0a010304020a0b0b0104;
    encBuf[4511] = 256'h03000d0d0a080102000a0d0b09010301090b0b09040602000909000505030009;
    encBuf[4512] = 256'h0c09000203010b0c0a020502090e0c09010202090d0c08010402080a0b090305;
    encBuf[4513] = 256'h01090c0a00040402080a09000303000c0c0a000303080a0b090103000c0f0b09;
    encBuf[4514] = 256'h0800000908010305030201000100090c0c0902060402080a09080304010b0f0b;
    encBuf[4515] = 256'h0a000301090c0b09040502080c0d0a00020400080a0901050301090c0a000305;
    encBuf[4516] = 256'h01090b0a00050401090d0b090002010a0d0b08030602080a0b09000402000a0c;
    encBuf[4517] = 256'h0902050302090b0b000203000a0d0a0004020208090a08080a0f0b0c08000100;
    encBuf[4518] = 256'h0100020402010a0c0c090102010101030705010100080800090e0d0b09010203;
    encBuf[4519] = 256'h01090a090202000c0f0b0901030301080901030602080a0c0a00010102010305;
    encBuf[4520] = 256'h0503010a0d0c0a080808090c0b08040503000b0c0b080202000c0b0a02070502;
    encBuf[4521] = 256'h00090808010108090c0b090103040100080a0b0b0c0a0900090b0b0a03070402;
    encBuf[4522] = 256'h090a0a0003020b0f0d0804050301080a090304020a0f0c09010302080b0e0801;
    encBuf[4523] = 256'h0403080c0c0a000303080b0c0903060200090b09020502090b0c08020302090c;
    encBuf[4524] = 256'h0a08040400090d0a080202010b0d0a08030402090b0b09030602000a0b080205;
    encBuf[4525] = 256'h03000a0b09020502080d0c09000303000c0c09010302090e0b09010403080a0c;
    encBuf[4526] = 256'h08030503010a0d0908030201090b0a01050401090c0a090101010a0b0c080203;
    encBuf[4527] = 256'h010a0c0c09000200090a080307060200080908010100090c0c0901040303080a;
    encBuf[4528] = 256'h0c0800010a0f0c0b08020202080a08030702000b0c0a00030300090902070401;
    encBuf[4529] = 256'h090b0b090202010a0b0a010404000a0d0b0a0a0b0a0b0a00040504040302000a;
    encBuf[4530] = 256'h0c0a090100080a09030706020109090900090a0d0c0b08020303000909090102;
    encBuf[4531] = 256'h080a0f0b0a08030603020001000102000b0f0b0901050401080a09010403090f;
    encBuf[4532] = 256'h0d0a08000201080a09020603010a0c0b09010302080c0a00060403000a0a0900;
    encBuf[4533] = 256'h02000a0e0b09020402080b0c09010302090d0b09030403080a0b08030502000b;
    encBuf[4534] = 256'h0d0901050302080909080102080c0e0b0a000101080909010305010a0c0b0802;
    encBuf[4535] = 256'h01080a0b0007050300080a00020403080b0d0a09010201090d0c0c0901030301;
    encBuf[4536] = 256'h0a0c0a000404010b0f0a00020402080a0b0805050208090b0a000302000c0b0b;
    encBuf[4537] = 256'h010302090e0d0900030400090c0b00040402080c0c09010403010a0b0a030703;
    encBuf[4538] = 256'h010a0d0a090202010b0d0b08030502080a0b09010302080c0c0901030301090a;
    encBuf[4539] = 256'h0003060201090a0800020108090b0c0c0a0b0a090809090a030705010b0d0b09;
    encBuf[4540] = 256'h0304010a0d0b02070402000a0a000203010b0f0b080303020a0c0b000203080e;
    encBuf[4541] = 256'h0c09000302000a0b08040501090c0b0802050200080902040401080b0b0a0909;
    encBuf[4542] = 256'h090b0c090002040100090a0b0c0c0b0a090002040304020404040401090b0b09;
    encBuf[4543] = 256'h030602000b0c090204020a0f0c09000202080b0c09020403080c0d0908020301;
    encBuf[4544] = 256'h09090004060301000a0a090102000c0c0b08020502090a0c090102080c0d0b0a;
    encBuf[4545] = 256'h010302000a0801060302000808010201090900060402090c0b000503000c0f0a;
    encBuf[4546] = 256'h080102010a0c0b080304010a0d0b09020402010808000305030300090c0c0900;
    encBuf[4547] = 256'h0303080d0c08030602080c0d0a010201090d0b09030503080b0b08030602090b;
    encBuf[4548] = 256'h0c08030502000b0a09020402080c0c0901020100090b0a080101090c0c0a0802;
    encBuf[4549] = 256'h0302000002050403080a0b09020302090d0803070501090b0b0a0100080b0d0b;
    encBuf[4550] = 256'h08020202080a0b090008090b0803070304020205030108090b0a090a00020405;
    encBuf[4551] = 256'h0201090a0b08080d0f0e0a0a00020101080800030401000a0a09080001030705;
    encBuf[4552] = 256'h0201080a080304000c0d0b08020401090c0b090200090d0c0901020200090106;
    encBuf[4553] = 256'h0402080b0c0a010303090c0902070401080a0a0801000a0d0c0a000201010809;
    encBuf[4554] = 256'h010402000c0d0a08010301090a0005060301080a0b080001000a0b0b08040502;
    encBuf[4555] = 256'h000a0c0b0a080a0b0d0b00030603010008020402090e0c0a01040300090b0105;
    encBuf[4556] = 256'h0502000c0b0b0002000a0d0b00030601080a0b080203000c0d0a010404010909;
    encBuf[4557] = 256'h08020402000b0d0a08030301090b0b000204000a0f0b0a08010301000a080107;
    encBuf[4558] = 256'h0301090b0b0a0001000908030707010009080101000b0f0b09010302090c0b08;
    encBuf[4559] = 256'h0504010a0d0a080203000a0d08020503010a0c09020402080c0b09010502000a;
    encBuf[4560] = 256'h0c0a000302000c0c0b0802050100090b09010303000b0e0a0803060200090908;
    encBuf[4561] = 256'h020402000c0b0a000202090d0b090205020a0c0c09010401080c0a0802040300;
    encBuf[4562] = 256'h0a0b0901050400090a0901040400090b0b0a0002010b0c0b09020403080a0a0a;
    encBuf[4563] = 256'h0a0a0c0c0a0802050200000206040300080909000200090b0c010304000b0c0c;
    encBuf[4564] = 256'h0800090c0e0c08020201090d0a08040303080d0c0a02050401000b0b08030602;
    encBuf[4565] = 256'h080b0e09000204010a0a0b080305010a0c0b0a010301090c0a0803060200090a;
    encBuf[4566] = 256'h09010102000809090104030303000c0e0b080202080d0e09000405010a0c0a08;
    encBuf[4567] = 256'h0203010c0e0a08030602080a0a08010302080c0d090002030300080909020201;
    encBuf[4568] = 256'h080d0e0c0908020302000a0a08050400090d0c09010301080a0a01060302080d;
    encBuf[4569] = 256'h0b090203020a0d0a00040502090b0c09010301090d0b08020502000a0a090002;
    encBuf[4570] = 256'h010a0c0b080204030000000305020a0d0c0a010201080b0b01070402090b0d09;
    encBuf[4571] = 256'h0101010a0d0a00040302090b0a000401090e0a09030602080a0a000403020a0f;
    encBuf[4572] = 256'h0b08010402080b0b09030602080b0e0908020201090c0a01040401090c0a0803;
    encBuf[4573] = 256'h03010a0d0a010404010a0c09000303010c0c0a00030301090d0a08010202080a;
    encBuf[4574] = 256'h0b0a0803030501080c0c08020503000b0d09010503000b0c0a010304080b0c09;
    encBuf[4575] = 256'h010402090b0c080203010a0d0a000502010b0b09010403000b0b080205020009;
    encBuf[4576] = 256'h09010101080d0b090101000b0d0a01030403090f0b0a010403020a0c0b080505;
    encBuf[4577] = 256'h02000a0d0a01030401090b0b00040401090b0c09010201080b0a08020401090d;
    encBuf[4578] = 256'h0a080000010008000205040201090b09040401090d0b0801050400090b0b0b00;
    encBuf[4579] = 256'h0302010a0a0b0a01050502000a0e0b0902030401090b09030703010a0c0b0900;
    encBuf[4580] = 256'h0103020801010009010503010d0f0c09000403010a0b09020702000b0c0a0104;
    encBuf[4581] = 256'h01080a0a000504000a0c0b010402080c0d08020502000b0c09020402080c0b09;
    encBuf[4582] = 256'h020402080a0a080403010c0b0a010303090d0b08040502090c0b000203030a0e;
    encBuf[4583] = 256'h0b0002040200090a09010301000a0b0808000002010203080e0c0a0a0203010d;
    encBuf[4584] = 256'h0c0a080307030109090b08000303000b0d0a02070301000a090102000b0f0b08;
    encBuf[4585] = 256'h0304010b0e0a010504000a0e0a080304010a0b0b00060401080b0b0802050209;
    encBuf[4586] = 256'h0b0b09020602080b0a090103010b0d0a080304010b0c0a020602000b0c0a0104;
    encBuf[4587] = 256'h03010b0c09020602000a0a0a010202000b0c080102020a0d09080202090f0b08;
    encBuf[4588] = 256'h010403000a0d09010502020a0c0a08030602080a0b0a020404080a0d09080203;
    encBuf[4589] = 256'h000a0c0a010201090c0b000304000b0c09040602000b0c09030502090b0b0003;
    encBuf[4590] = 256'h0601090c0a000202080b0d09010401090d0a000303020c0e0900030402090c0a;
    encBuf[4591] = 256'h00030501090b0c08020402080b0c09010302090c0b0a000302090c0b08020501;
    encBuf[4592] = 256'h090d09080305010a0c0a01040501090b0b08030502080c0b09010303000c0d09;
    encBuf[4593] = 256'h000202080b0d09010203000b0b09030601080c0a08040302090c0b0804040109;
    encBuf[4594] = 256'h0b0c09000303080b0b0b00030503000b0d0a0002050401090b0a00050303000b;
    encBuf[4595] = 256'h0c0901030501090b0b0a0a000401090c0b0d09030402080c0b09010602000a0a;
    encBuf[4596] = 256'h08050402000a0b020503000b0e09010304000c0c0a000303000d0d0a08010201;
    encBuf[4597] = 256'h090c0a09010302010a0c0a0802050201080809090305030100090b0b00030305;
    encBuf[4598] = 256'h010a0b0b0c080502000b0d0c08000000090c0a09080a0c0c090800090e0d0c09;
    encBuf[4599] = 256'h0203000b0f0a090203020a0c0b08030702000909000304030000010204030101;
    encBuf[4600] = 256'h02030304000a09090304090c0c0c0a00000a0b0e0c0a0a080009090a0b0b0a0a;
    encBuf[4601] = 256'h080403010c0f0b00010502000b0e09000101080b0f0b0a0001000b0d0c0a0900;
    encBuf[4602] = 256'h080a0a0d0a080008080808020203020a0a050604030109000004060202080a09;
    encBuf[4603] = 256'h0003040208090b0b000300080b0f0d09090809080a0b0b090a0908090a000a0e;
    encBuf[4604] = 256'h0a0a000507010809090106040201090801050502010001010404030001000204;
    encBuf[4605] = 256'h0202080801030302090d0b0901010a0f0c0b0a09080a0c0d0b0a09090a0a0b0c;
    encBuf[4606] = 256'h0b09080808000009090a080107030100090a03050401090b0c0c0900080b0b0f;
    encBuf[4607] = 256'h0d09090a090b0e0a0c09090b0b0b0d0a090a0b0b0e0a09090a0b0d0b0b090000;
    encBuf[4608] = 256'h0b0e0c0a080102080a0d0a080204020008080206050203010104030504020103;
    encBuf[4609] = 256'h02050304010202020403030201010204040201080801020302000b0c09010202;
    encBuf[4610] = 256'h0a0e0a090802000a0a0b0a020501010102070402040202050402030303040502;
    encBuf[4611] = 256'h04030203030305030203020102030304020008080101010b0b0f0b09000b0b0c;
    encBuf[4612] = 256'h0c09000002000a02060505030202040405040203020304040303030302030403;
    encBuf[4613] = 256'h03020100000001090b0e0c0c0b0b0c0c0c0a0c0a0b0b0c0a0c0a0a0b0b0a0c0a;
    encBuf[4614] = 256'h0a0a09080a0a0a0b0a08090a0e0c0b0b0c0b0c0e0b0b0d0a0c0b0c0c0b0b0c0b;
    encBuf[4615] = 256'h0c0b0c0a0b0b0c0b0b0b0b0c0a0b0b0a0b0a09090a0909080102020301020603;
    encBuf[4616] = 256'h03050101030002030008080f0a080b0c0b0f0b0a0b0b0b0e0b0a0c0a0a0a0b0a;
    encBuf[4617] = 256'h0c0a090808000900020305050302040304050303030304040303040202030303;
    encBuf[4618] = 256'h050102020102030202030000050101030009030102060809000a09030b0d0a0f;
    encBuf[4619] = 256'h0b0a0d0b0c0d0c0a0c0b0b0d0b0c0b0c0b0b0c0b0c0a0b0b0b0b0b0b0a090808;
    encBuf[4620] = 256'h0104030605040305030503040403030404030305020304020304020303040203;
    encBuf[4621] = 256'h0203030303020302020201010808080a0b0c0d0a0c0c0a0c0b0a0c0b0a0c0a0a;
    encBuf[4622] = 256'h0b0b0a0a0b090a0a08080801010004020205030204020202020001090b0c0e0c;
    encBuf[4623] = 256'h0c0d0b0c0c0c0b0c0b0d0b0b0c0b0c0b0c0b0c0b0b0b0c0b0b0b0c0b0a0b0b0a;
    encBuf[4624] = 256'h0b0a0a0909090000020403060304040305030304030304030303040203030302;
    encBuf[4625] = 256'h020202010008090a0c0c0c0c0b0c0c0b0c0b0c0a0b0c0a0b0b0b0b0b0b0c0a0a;
    encBuf[4626] = 256'h0a0a0a09090808080100020202020201000209090a0e0c0b0c0b0c0c0b0c0b0b;
    encBuf[4627] = 256'h0b0d0b0b0b0b0b0c0a0909000203050504030404020402030304020402020402;
    encBuf[4628] = 256'h03030303050102020100020900000a0a000d0a080e0a0a0e0b0a0e0c0a0c0c0b;
    encBuf[4629] = 256'h0c0b0c0c0b0b0c0c0b0b0c0b0b0c0b0c0a0b0b0b0b0a0b0a0808000305040405;
    encBuf[4630] = 256'h0305030404030403040304030304040203030402030203020302020201000008;
    encBuf[4631] = 256'h080a0b0d0c0b0d0b0c0b0d0a0b0c0a0b0b0b0b0b0b0b0a0a0909000000030404;
    encBuf[4632] = 256'h040305030403040303040203030202010108090a0c0d0c0c0b0d0b0c0c0b0b0d;
    encBuf[4633] = 256'h0b0b0b0c0b0b0b0b0c0b0b0a0b0b0a0a09090900010204040404030503050303;
    encBuf[4634] = 256'h04040303040303040303030304020302030203020202010000080a0a0d0b0d0b;
    encBuf[4635] = 256'h0c0c0b0b0c0a0c0a0a0b0b0a0b0a0b0a0a0a0908080102030604030503030502;
    encBuf[4636] = 256'h0302030202010100080a0b0c0d0c0c0c0b0c0c0b0c0c0b0b0c0b0c0b0b0b0b0a;
    encBuf[4637] = 256'h0b0b0a0909000001030404040404030503040304030403040203030303020302;
    encBuf[4638] = 256'h020201000009090a0c0c0c0c0b0d0b0c0c0a0c0b0b0b0b0b0c0a0b0a0a090909;
    encBuf[4639] = 256'h0808000102030306030404040304030304030303020302010008090a0b0e0b0d;
    encBuf[4640] = 256'h0b0c0c0b0c0c0b0b0c0c0b0b0b0c0b0b0b0a0b0b0a0909080801020305030504;
    encBuf[4641] = 256'h0304040304030403040303040302030203020102000008080a0a0b0d0c0b0d0b;
    encBuf[4642] = 256'h0c0b0d0b0b0c0b0c0a0b0b0a0b0a0a0a09090808080001000201020303040403;
    encBuf[4643] = 256'h04040202030100000a0b0f0c0b0c0c0b0c0b0a0b0a090a080001020503050403;
    encBuf[4644] = 256'h0504040304040403040303040302030303030203030303040202020201010000;
    encBuf[4645] = 256'h090a0b0e0c0b0d0b0c0b0b0c0b0b0b0b0b0b0b0b0b0a0b0b0a0a0a0901010306;
    encBuf[4646] = 256'h0404040303050202030201010008090a0c0c0c0c0b0c0c0b0c0c0b0d0b0b0c0c;
    encBuf[4647] = 256'h0b0b0c0b0b0b0b0b0b0c0a0a090a090908080000020305040405030403050303;
    encBuf[4648] = 256'h0403040203030304020303030402030203020301020000080a0b0c0d0b0c0b0c;
    encBuf[4649] = 256'h0b0b0b0c0b0b0b0c0b0c0b0b0b0c0a0b0a0a0908080101030304040302030303;
    encBuf[4650] = 256'h020201020202020200020008090f0e0c0d0b0d0b0d0b0b0c0b0a0b0b0b0b0a0a;
    encBuf[4651] = 256'h0a0b0a0c090a0809080002060405030404030503030303040303030303040204;
    encBuf[4652] = 256'h020303020302030101090a0c0c0c0b0d0c0a0b0b0c0b0b0b0c0b0b0c0b0c0b0c;
    encBuf[4653] = 256'h0a0b0b0b0c0a0909090808080101000100000008000008000102050302030201;
    encBuf[4654] = 256'h020a0f0d0c0d0a0c0c0b0b0c0a0b0b0b0b0b0b0b0b0b0c0b0b0b0a0808020405;
    encBuf[4655] = 256'h060403050304030403030402030304020303020402010202000108090a0c0d0b;
    encBuf[4656] = 256'h0d0c0a0c0b0b0c0b0b0b0c0b0b0c0a0b0b0a0c0b0a0a0b0a0b0a0a0a0a0a0c0b;
    encBuf[4657] = 256'h0a0c0b0c0c0c0b0c0b0c0b0b0d0a0b0a0b0a0b0a080901030307040504040305;
    encBuf[4658] = 256'h0304040304030403030503030304030402030303020303030202020101000809;
    encBuf[4659] = 256'h0b0c0d0b0c0c0b0d0b0b0b0c0b0b0c0a0b0b0a0b0a0a09090808000101030603;
    encBuf[4660] = 256'h040305030304030402020202010100080a0b0d0c0c0c0c0b0c0c0c0a0c0b0b0c;
    encBuf[4661] = 256'h0c0a0b0c0b0a0c0a0a0b0a0a0a0a0a0909080000020204050403050304040304;
    encBuf[4662] = 256'h030403030304030304030203030303030303030202000008090b0d0c0c0b0c0c;
    encBuf[4663] = 256'h0b0b0c0b0c0b0b0b0b0c0b0b0b0c0a0b0a0a0a09080900000103030305030304;
    encBuf[4664] = 256'h0203030202020201010808090b0c0d0d0c0c0b0d0b0c0c0b0b0b0b0b0c0a0a0a;
    encBuf[4665] = 256'h0909080908000101030306040404030503030503030304030303030303030302;
    encBuf[4666] = 256'h030203010201010008090d0c0c0c0b0d0b0c0b0b0b0b0b0c0b0a0b0b0c0b0b0b;
    encBuf[4667] = 256'h0c0a0b0c0a0b0c0a0a0b0a0b0a0a0a0c0a0d0b0d0b0d0b0c0c0b0a0c0a0b0c0a;
    encBuf[4668] = 256'h0a0b0b0c0b0c0a0b0b0c0a0b0a0a0a0900000203070304040305030304030404;
    encBuf[4669] = 256'h03030403030502030303030402020202010000080a090c0c0b0c0b0c0c0c0a0c;
    encBuf[4670] = 256'h0b0b0d0b0a0c0b0a0b0b0b0b0a0b0a0b0a0a0a09090909090a090a0a0c0b0c0a;
    encBuf[4671] = 256'h0b0c0b0c0c0c0b0d0c0b0c0c0a0a0b0a0a0a0801010306030604040305040303;
    encBuf[4672] = 256'h050304030305020403020403030303030303030203020102010000080a0b0d0c;
    encBuf[4673] = 256'h0c0c0b0c0c0b0b0c0b0b0c0b0b0b0b0a0b0a090a080800010101040305030404;
    encBuf[4674] = 256'h040304030303030203010100090b0b0e0c0c0c0c0b0c0c0b0c0b0c0b0b0d0a0c;
    encBuf[4675] = 256'h0a0b0b0c0a0b0a0b0a0a0a090a08080001020304040405030403050303050303;
    encBuf[4676] = 256'h0304030402030302030303030303030202020000080a0b0d0d0b0d0b0c0b0c0a;
    encBuf[4677] = 256'h0c0a0b0b0b0b0b0b0c0b0b0b0b0b0b0b0a090900010204030503030403020303;
    encBuf[4678] = 256'h0302020102000000090a090c0a0b0f0c0c0c0c0c0b0c0b0b0b0b0a0909080000;
    encBuf[4679] = 256'h0202020202040504040403040404030403030403040203020302030201010100;
    encBuf[4680] = 256'h010102000000090a0c0e0d0b0d0b0c0a0c0a0a0b0a0a0a0b0a0b0b0b0b0c0c0a;
    encBuf[4681] = 256'h0b0a0b0a0a0b090800010202030401000a0e0c0d0c0b0c0b0b0c0a0b0a0c0a0b;
    encBuf[4682] = 256'h0d0b0b0d0b0c0b0c0a0b0a0a0a09080800010204020403030503040404030403;
    encBuf[4683] = 256'h040403040303030403020203010201010100080008090a0b0f0c0b0d0c0b0d0b;
    encBuf[4684] = 256'h0b0c0b0b0b0c0b0b0b0b0b0c0a0b0a0a0b0a0a0a0a0809080202040503050302;
    encBuf[4685] = 256'h03020000080a0a0a0a0b0c0b0b0d0c0c0c0c0b0c0a0b0a0a0809000202040604;
    encBuf[4686] = 256'h0504040305030404020304030304030403040303030304020202020201010101;
    encBuf[4687] = 256'h0000090a0b0e0b0d0b0c0b0b0d0a0b0b0c0b0b0c0a0b0a0b0a09090900000801;
    encBuf[4688] = 256'h01010304030603040403030402030201020008080a0b0b0e0c0c0c0c0b0c0c0b;
    encBuf[4689] = 256'h0b0d0b0b0c0b0c0b0b0b0c0b0a0b0b0a0a0b0909090008010204040503050403;
    encBuf[4690] = 256'h040305020304030303040303030402030302030302020201010808090c0b0d0c;
    encBuf[4691] = 256'h0c0b0c0b0b0c0b0b0c0b0b0b0c0a0b0c0a0b0a0a0a0a09000801020202050203;
    encBuf[4692] = 256'h0403030404020303030402020201020102010201080a0d0d0c0c0b0c0b0a0a0a;
    encBuf[4693] = 256'h0909080809080b0c0c0b0a080802040404040403030304030403040303030403;
    encBuf[4694] = 256'h02020201020402040202020301000a0c0d0c0b0b0c0b0b0b0b0a0a0c0c0b0c0c;
    encBuf[4695] = 256'h0b0c0b0b0c0b0b0b0b0c0b0a0a0a0a0a0b0b0b0d0c0b0e0b0b0c0b0a0b0b0a0a;
    encBuf[4696] = 256'h0a0a0c0b0c0b0c0b0b0c0a0b0a0a090809010204050503040403040202030302;
    encBuf[4697] = 256'h0404030404030403030203020202010001080008090a0b0d0c0b0c0c0a0b0c0b;
    encBuf[4698] = 256'h0c0c0c0c0b0c0b0c0a0a0b090a090a090a0b0b0c0b0b0b0a0a09000001020103;
    encBuf[4699] = 256'h0603040502030403020108090a0d0b0b0b0a090909090d0c0e0c0c0c0b0b0b0b;
    encBuf[4700] = 256'h0a0a0a0008000302050504040404040403030403040304030404030304020303;
    encBuf[4701] = 256'h0203020201020201020201010108090c0b0e0c0b0d0b0b0c0b0b0c0b0c0b0a0b;
    encBuf[4702] = 256'h0b0b0a0b090a0909080a00080802020505030504030303040202010101080909;
    encBuf[4703] = 256'h0a0b0c0d0b0d0c0a0c0c0b0c0b0c0c0b0b0c0b0c0a0b0a0b0b0b0a0a0a0a090a;
    encBuf[4704] = 256'h0800000103030703050404030404030304030402030303040203030303040203;
    encBuf[4705] = 256'h020201020008080a0b0c0d0b0d0b0b0c0b0c0a0b0b0c0a0b0c0a0b0c0a0b0b0a;
    encBuf[4706] = 256'h0a09090800010103040403030403040203040303030404030403040202020201;
    encBuf[4707] = 256'h0008090a0a0b0c0b0b0b0b0a0c0c0d0b0c0c0a0c0b0c0b0b0c0a0a0a0a0a0809;
    encBuf[4708] = 256'h0801000002020001080803050604040403040403030302030202020201010200;
    encBuf[4709] = 256'h0008090b0a0e0c0b0d0c0b0c0d0b0c0c0c0b0b0b0b0b0b0b0c0a0b0b0c0b0b0c;
    encBuf[4710] = 256'h0b0c0a0909080800000001030305030404030304030303030403030504030403;
    encBuf[4711] = 256'h030302020000000008000001010101000a0c0b0f0a0b0c0a0b0a0b0b0c0c0b0d;
    encBuf[4712] = 256'h0b0a0a0a000802020008090c0c0a0b0c090a08010306040101010a0a0b0d0a0a;
    encBuf[4713] = 256'h0a08080b0a090a08020908010b08050002000e0c0a0c0a090a08010800090f0d;
    encBuf[4714] = 256'h0c0d0a0c0b0b0b0d0a0c0b0b0c0b0b0a09080001040305040302050305050305;
    encBuf[4715] = 256'h0403040304030303040303040402030402030202020202010100010000090a0b;
    encBuf[4716] = 256'h0e0c0b0d0b0c0b0b0c0b0b0b0c0b0b0b0c0b0b0b0b0a0a080800080101020403;
    encBuf[4717] = 256'h040403030502040202030301020009080b0c0c0d0c0c0c0b0c0b0c0b0c0c0a0c;
    encBuf[4718] = 256'h0a0b0b0b0c0a0b0b0b0b0b0b0a0a0a0800010403050502040403030403040403;
    encBuf[4719] = 256'h0305020303040302030304020202020202010001000909090b0c0c0b0d0b0c0c;
    encBuf[4720] = 256'h0b0b0d0b0a0c0a0b0b0b0a0b0c090a0a09090900080001020204040205030405;
    encBuf[4721] = 256'h03040303020302020202020203030402030201000b0e0d0b0c0b0a0b0c0c0b0b;
    encBuf[4722] = 256'h0b0c0c0a0c0a0a0a0a0a0a0a0a0b0b0b0c0b0800020504030403040202010202;
    encBuf[4723] = 256'h04030503030403030303010100000808090b0a0d0e0b0e0c0b0b0c0a0c0a0b0b;
    encBuf[4724] = 256'h0c0a0c0b0c0b0b0c0b0b0a0a0909080908090800000100020204050403040403;
    encBuf[4725] = 256'h0305030304030304020202020102020202040204030202020008000800000a09;
    encBuf[4726] = 256'h080b09080c0c0c0c0b090801030303010c0f0c0c0b0a0b0b090908000100080b;
    encBuf[4727] = 256'h0f0d0c0b0b0b0a0809090a0c0d0a0b0b090a0a080003050201010b0d0b0d0a08;
    encBuf[4728] = 256'h01030703040301020108080a0c0c0b0b090a0a0a0b0d0b0d0b0c0b0d0a0b0b0b;
    encBuf[4729] = 256'h0c0a0a0b09080900020207060306040303050303040303040303050304040204;
    encBuf[4730] = 256'h020302020301020101000101000000080a0b0d0c0c0c0c0b0b0d0a0c0a0a0b0c;
    encBuf[4731] = 256'h0a0b0b0a0b0b0a0a0a0909090809080800010204050404040303040102010008;
    encBuf[4732] = 256'h08090a0b0c0b0b0c0d0b0c0d0b0d0b0b0c0b0c0b0c0a0b0c0a0a0b0a0a0a0a08;
    encBuf[4733] = 256'h0800010102030305040404040403040403040303040302030303030402030303;
    encBuf[4734] = 256'h03030203010208080a0c0c0c0c0c0b0c0b0c0a0b0b0c0a0b0b0b0c0b0c0b0b0b;
    encBuf[4735] = 256'h0c09090900000102020403040303040304030303040303040203020303020201;
    encBuf[4736] = 256'h00090b0e0c0d0c0b0c0c0a0b0b0b0b0b0b0b0b0b0c0b0c0b0b0b0b0a09080102;
    encBuf[4737] = 256'h040503050305020402030304030303020302020202020201010108090b0d0e0c;
    encBuf[4738] = 256'h0c0c0c0b0b0c0a0b0c0a0b0b0c0b0b0c0a0b0a0a090908080100010103030503;
    encBuf[4739] = 256'h04040304040402030303030303030303030102010808090b0b0d0b0b0b0b0a0b;
    encBuf[4740] = 256'h0b0e0b0e0a0b0a09080002050404030402020202040204030204030302030001;
    encBuf[4741] = 256'h000000020808080d0c0e0d0b0d0b0b0b0c0b0a0b0b0b0b0c0b0c0b0b0b0a0a0a;
    encBuf[4742] = 256'h0a09090900010204040404040204030303040202020103020203090a0b0f0a09;
    encBuf[4743] = 256'h0b0b0b0f0b090b0a0a0e0b0d0c0b0c0b0c0a0b0a0a0a090a09090a0a0c0d0a0a;
    encBuf[4744] = 256'h0a08000104040404050204030405030503040304030303040203040304040303;
    encBuf[4745] = 256'h040302030102010101010001000008090b0c0c0c0c0b0d0a0c0b0b0c0c0b0b0c;
    encBuf[4746] = 256'h0b0a0b0a090a09090908090a090a0b0909000404040504030402030302010100;
    encBuf[4747] = 256'h000a0a0c0b0d0b0c0b0b0c0c0b0c0c0b0d0b0b0c0b0c0a0b0b0a0b0a0a0a0909;
    encBuf[4748] = 256'h0800020403040403050304030503040304030403030402020302020303020402;
    encBuf[4749] = 256'h020203010101080a0b0d0d0b0c0c0b0b0c0b0b0b0c0a0b0a0a0a0b0b0c0b0b0b;
    encBuf[4750] = 256'h0c0a0a090001020504030503040203010202020102020201000109090b0c0e0c;
    encBuf[4751] = 256'h0b0d0b0c0a0b0b0c0c0b0c0b0c0b0a0b0b0a0b090a0909080808010104040603;
    encBuf[4752] = 256'h050303040202020203020403030403040202020000090a0a0c0c0b0d0b0c0c0b;
    encBuf[4753] = 256'h0c0b0c0a0a0b0a0a0a0a0b0c0b0b0b0b0b090800020504040303030302030305;
    encBuf[4754] = 256'h030503030403030303030302010108080a0b0c0a0c0b0b0d0b0a0a09090a0b0d;
    encBuf[4755] = 256'h0c0c0b0b0b0b0a0a000003070404040303030201020203040303040100010809;
    encBuf[4756] = 256'h0109090a0f0c0c0c0c0c0c0b0c0b0b0b0a0b090b0a0c0b0b0c0a0a0908080101;
    encBuf[4757] = 256'h02040305030305030304030303030303050303040201020108000a0c0b0d0b0c;
    encBuf[4758] = 256'h0b0c0a0c0b0b0c0a090908090a0c0d0d0b0b0c0a0a0a08080001020303010200;
    encBuf[4759] = 256'h0800020107050404040204030305040305030503030304030302030403040403;
    encBuf[4760] = 256'h050203030302020101000100080008090a0b0d0c0c0c0c0b0b0d0b0b0c0b0c0b;
    encBuf[4761] = 256'h0b0c0b0a0b0a09090a0808090808080800010304050404030402030302020202;
    encBuf[4762] = 256'h010108090a0d0c0c0c0b0c0b0c0b0c0b0d0b0c0b0c0b0b0b0b0b0a0a0a090909;
    encBuf[4763] = 256'h0809000001020504050403050304040203040303040303040203020302010201;
    encBuf[4764] = 256'h0201030203020201090c0c0e0b0c0b0c0a0b0a0a0b0a0b0c0b0b0d0a0a0a0909;
    encBuf[4765] = 256'h080800080000010104030703030402020201000008080000010200000a0f0c0d;
    encBuf[4766] = 256'h0c0c0c0b0c0a0b0b0a0b0c0b0b0c0b0b0a0b0a09000800000000080a09000307;
    encBuf[4767] = 256'h0705030303030302010101000001010201010100080a0d0c0c0c0b0c0b0b0d0c;
    encBuf[4768] = 256'h0b0b0c0b0b0b09090000010102010100090a0d0a090206060404040203020101;
    encBuf[4769] = 256'h00000800000000020304030101000b0b0c0b0c0b0d0c0b0d0b0b0a0a09090a09;
    encBuf[4770] = 256'h0909080000000008000802060504040304040203040203030101000808080a0b;
    encBuf[4771] = 256'h0d0d0d0a0c0a0a0b0b0c0c0b0d0b0b0c0b0b0b0c0a0a09080800010001010202;
    encBuf[4772] = 256'h0404040503040305030303020303020303030304020202080a0a0f0b0b0c0a0b;
    encBuf[4773] = 256'h0b0b0b0e0b0b0d0b0b0b0a0a0b09080802030302000909080205030603040305;
    encBuf[4774] = 256'h0203030201010801010206050304030304050404050304030304030303040304;
    encBuf[4775] = 256'h0403030503030402030201010108000808090a0a0a0b0d0b0d0c0c0b0d0b0c0b;
    encBuf[4776] = 256'h0c0a0b0b0a0c0a0a0a0a090a0908090808000001010303030603050503040302;
    encBuf[4777] = 256'h030201010008080a0b0b0e0b0d0b0c0a0c0b0b0c0b0c0b0c0b0c0b0c0b0a0b0b;
    encBuf[4778] = 256'h090a080800020204040403040402030403040403040304030304030302030202;
    encBuf[4779] = 256'h01020101020001000009090c0d0b0d0c0b0c0b0b0c0b0b0b0b0a0a0a0a0a0909;
    encBuf[4780] = 256'h0a080a090800010404060503040402020202010200000909090a0a0b0b0d0c0d;
    encBuf[4781] = 256'h0b0c0c0c0b0c0c0b0b0c0b0b0b0b0a090a090909080909080808000204050404;
    encBuf[4782] = 256'h0403040403020402020202010000000909090a0a0b0b0b0c0c0c0c0b0c0b0c0b;
    encBuf[4783] = 256'h0c0c0b0a0b0b0a09080808010204040403030303030304040303050305030303;
    encBuf[4784] = 256'h0403030101080a0a0a0b0a0e0b0d0b0a0a0a0908090a0a0c0d0b0d0b0c0a0b0a;
    encBuf[4785] = 256'h0a0800020504030303020303030403020202020101010002010203000a0c0f0b;
    encBuf[4786] = 256'h0c0d0c0c0c0c0a0b0b0b0c0a0b0b0c0a0a0a0908000102030503050403030301;
    encBuf[4787] = 256'h0202030505040304030403030203010008080a0b0b0b0b0b0b0c0d0c0c0a0b0a;
    encBuf[4788] = 256'h0a0a0b0d0b0c0c0b0b0c0a090800020403040202020101000800010104030402;
    encBuf[4789] = 256'h0202020001010800010a090a0e0a090a08010005070705050305030303040203;
    encBuf[4790] = 256'h03040303040304040304020303020201010008080a0a0b0d0b0b0d0b0c0c0c0b;
    encBuf[4791] = 256'h0c0b0c0b0b0c0a0c0a0b0a0b0a0a0a0908090000000100010202030504050304;
    encBuf[4792] = 256'h04030302030201080808090a0b0d0c0c0c0c0a0c0b0b0b0c0b0c0b0b0c0b0c0b;
    encBuf[4793] = 256'h0a0b090909000202030503040304040402040402040303040303030402030302;
    encBuf[4794] = 256'h0302010201010000090809090b0b0e0b0d0c0c0b0c0a0b0b0b0b0b0a0b0a0909;
    encBuf[4795] = 256'h0908080003040404040203030204030305030403040102000009090c0b0d0b0c;
    encBuf[4796] = 256'h0b0c0b0c0c0b0b0b0c0b0b0c0b0b0b0c0a0b0b0b0a0908000102030404030404;
    encBuf[4797] = 256'h0303040203020303030404020202000008080b0d0c0d0b0b0c0c0b0b0c0c0a0b;
    encBuf[4798] = 256'h0a0a0b0a0b0b0b0c0b0a09080103040403050304040303040203020303030303;
    encBuf[4799] = 256'h03040302020108090b0e0b0d0c0c0b0c0b0b0a0a0a09090a0b0a0c0a0a090900;
    encBuf[4800] = 256'h080103050504030503030503030302010101000001020403030302080a0a0d0b;
    encBuf[4801] = 256'h0b0e0c0c0c0c0b0b0b0a0a0808080808090a0c0b0c0a0a080203050304030403;
    encBuf[4802] = 256'h04040305040203030202010000000908000800010909080e0c0c0c0d0b0d0b0b;
    encBuf[4803] = 256'h0b0c0a090a08090808090a0a0b09080103050404040303030402030404030502;
    encBuf[4804] = 256'h020100090a0c0c0b0b0b0a09090a090c0c0c0d0b0b0b09000004030305040305;
    encBuf[4805] = 256'h040503050403030403040203020303040304030403030202010009090a0b0d0b;
    encBuf[4806] = 256'h0c0b0b0b0d0c0b0c0c0b0c0a0b0c0a0b0a0b0b0b0a0a0a080801020305030502;
    encBuf[4807] = 256'h030203030404030404030402030202010108090a0b0d0c0b0d0b0b0d0a0b0b0c;
    encBuf[4808] = 256'h0a0b0c0b0c0b0b0c0b0a0a090900000203030503040305030403040304030304;
    encBuf[4809] = 256'h03030304030303030202010109090b0c0b0b0b0b0b0d0c0b0c0c0b0c0c0a0b0b;
    encBuf[4810] = 256'h0a0a080908000001010205030503040303030304020303030402020202000009;
    encBuf[4811] = 256'h0d0c0c0d0b0b0c0c0b0b0c0b0c0b0c0b0a0b0b0a0b0a0a0a090a090908090001;
    encBuf[4812] = 256'h0306050403050302030303030203020202020202030200000b0e0d0c0b0c0c0b;
    encBuf[4813] = 256'h0c0a0c0a0a0b0a0a0a0a09090808000102020305030504040305020303040203;
    encBuf[4814] = 256'h030303030301000b0c0d0b0b0b0a09090a0b0d0d0c0c0c0b0b0a0b0908000002;
    encBuf[4815] = 256'h0301020000030505040403020304020402030302030203030303010a0c0e0c0c;
    encBuf[4816] = 256'h0a0a0a0a0b0b0b0e0b0c0b0c0b0c0a0a0909080809080a0a0a09080202040402;
    encBuf[4817] = 256'h03040202020304030503030201080b0e0a0b0a090800010808080b0d0c0e0b0c;
    encBuf[4818] = 256'h0a0a00020404020100090a0a0900050404040303030000090b0a090802040303;
    encBuf[4819] = 256'h03090c0d0e0a0a0a090008080a0b0e0c0c0b0b0b0b0c09090908010102040304;
    encBuf[4820] = 256'h0502040403040404030404040403040304030403020303030303030404030304;
    encBuf[4821] = 256'h02020100090a0c0b0c0c0b0c0b0b0c0b0c0c0b0c0b0b0b0c0a0b0b0a0b0a0a09;
    encBuf[4822] = 256'h0908000104030504040203030303040203030304020302020200090b0e0d0c0b;
    encBuf[4823] = 256'h0d0b0b0c0b0c0c0a0b0a0b0b0c0a0b0a0a0a0909090008010204050405030403;
    encBuf[4824] = 256'h03040303040303040203030303030202020201010008090c0c0d0c0b0c0b0b0b;
    encBuf[4825] = 256'h0a0a0a0a0a0a0a0b0b0a0a080104060304040204020403030403030304020101;
    encBuf[4826] = 256'h00090a0b0c0c0c0b0c0b0d0b0c0b0b0c0b0c0b0b0c0b0b0a0b0a0a0a09080801;
    encBuf[4827] = 256'h02020404030503030503030404020402030203020101000809090a0b0c0b0b0d;
    encBuf[4828] = 256'h0c0b0d0b0c0b0c0a0b0b0a0b0a0a090a08090800010305040503040304020303;
    encBuf[4829] = 256'h0303040203020302010100090a0d0d0b0c0c0b0b0b0c0c0b0a0c0a0a0b0a0909;
    encBuf[4830] = 256'h090000020205030305020305030306030403030402020101010008000008080a;
    encBuf[4831] = 256'h0a0c0d0b0d0b0b0b0c0a0c0a0b0b0c0b0d0a0b0a0b0909090808000102020303;
    encBuf[4832] = 256'h02010809080004050503040201000808090a0a0b0c0b0a0c0909080003020503;
    encBuf[4833] = 256'h0305040205030503060304030403040203030303020201010009080b0a0a0b0c;
    encBuf[4834] = 256'h0a0d0c0d0c0c0b0c0c0b0b0c0a0b0a0a0a090008010000000100010102010205;
    encBuf[4835] = 256'h0404040403030502030303040303020301020402030503040503050404040403;
    encBuf[4836] = 256'h0303040203020302030403030502040202020100080a0b0d0c0c0c0b0c0a0b0c;
    encBuf[4837] = 256'h0a0b0b0b0c0b0c0a0c0a0a0a0b09090a08000003040404040304030304020302;
    encBuf[4838] = 256'h02010201010101010100090b0f0d0b0e0b0b0c0c0a0b0b0b0b0c0b0a0b0a0a0a;
    encBuf[4839] = 256'h0908000102040404030404040304030403040302030402020202010201000008;
    encBuf[4840] = 256'h080a0a0c0c0c0b0b0c0b0c0b0c0b0b0b0b0b0a0a090900020306040304040303;
    encBuf[4841] = 256'h030403030304020303040303020101090a0d0c0d0b0d0b0c0b0b0b0c0b0b0b0c;
    encBuf[4842] = 256'h0a0b0a0b0a0b0a0b0b0a09080103050504040304030303030302030203030303;
    encBuf[4843] = 256'h01010008090a0d0b0d0c0b0b0c0b0c0b0b0c0c0b0b0a0a090801030404040304;
    encBuf[4844] = 256'h020302020102020303040303020101090a0d0c0d0c0c0b0d0b0c0a0b0c0a0a0b;
    encBuf[4845] = 256'h0a0a0a0a0a0a0908000002030503050305030403050203030203020100000809;
    encBuf[4846] = 256'h0a0a0c0a0b0d0c0c0c0c0b0d0a0c0a0a0b0b0a0a0a0a0a0a09090a0808010203;
    encBuf[4847] = 256'h040401020201030503020201000008090a0b0c0d0c0c0b0c0b0b0c0a090a0900;
    encBuf[4848] = 256'h0003050304040305040404030305030303040203030303030403030202010808;
    encBuf[4849] = 256'h0a0d0b0c0d0b0b0d0b0a0c0b0b0c0b0b0c0b0a0b0a0b0b0c090a080001010403;
    encBuf[4850] = 256'h050503040303020202010201010100000909090b0a0b0d0b0c0d0a0a0b0b0b0c;
    encBuf[4851] = 256'h0b08080307070306040305040303030403030303040203030304030203020100;
    encBuf[4852] = 256'h0a0b0e0c0b0d0b0c0c0b0b0b0c0b0b0c0b0b0b0b0b0a0a0a0909080002030504;
    encBuf[4853] = 256'h0503040403040303040202020201010100000008090b0c0c0c0d0b0d0b0b0c0b;
    encBuf[4854] = 256'h0c0b0b0b0a0b0b0a0a0a09080000030405030504030305030303040304020303;
    encBuf[4855] = 256'h03030201010808090b0b0d0c0b0c0b0b0c0b0c0b0c0b0b0b0b0b0a0908000104;
    encBuf[4856] = 256'h040404040304030304040203030302030202020108090a0b0e0b0d0b0d0b0c0c;
    encBuf[4857] = 256'h0b0b0c0b0c0a0b0a0b0a0b0a0a0a090808010205030503040402030402030304;
    encBuf[4858] = 256'h020302030302020100080a0a0c0b0c0c0b0c0b0c0c0a0a0b0a0a0b0909080801;
    encBuf[4859] = 256'h01020305040403050304030303030302020100080a0c0c0c0b0d0b0b0c0b0c0b;
    encBuf[4860] = 256'h0b0b0c0b0b0b0b0c0a0a09090002030603040403030403040203030402030201;
    encBuf[4861] = 256'h0108080a0c0c0c0c0b0b0b0c0c0b0b0b0b0c0b0b0b0a0b0a0a09080002020504;
    encBuf[4862] = 256'h0304040304020303040202030303030201080a0d0c0c0c0b0c0b0b0b0b0b0b0a;
    encBuf[4863] = 256'h0a0a080800020306040404030305030304040303050204020203020100000809;
    encBuf[4864] = 256'h090b0b0a0c0a0c0b0c0c0b0c0b0b0b0b0b0a0a0a0a0909080000020304050404;
    encBuf[4865] = 256'h040302010109090a0b0a0a08080001000b0f0d0e0b0d0b0c0a0b0a0a0a0a0a0b;
    encBuf[4866] = 256'h0a0a0a0800000405040504030404020304020303030404050305030503030303;
    encBuf[4867] = 256'h0402020201010201010101020000090b0e0c0c0b0d0b0b0c0c0a0b0b0b0c0b0c;
    encBuf[4868] = 256'h0b0a0b0a0a0a0908010102030504030404030403040303030202020200000809;
    encBuf[4869] = 256'h090b0c0c0c0b0e0b0c0c0b0c0b0b0c0b0a0b0a0b0a0909080800020203050404;
    encBuf[4870] = 256'h0304040304030402030303020203010200010809090c0c0c0c0b0c0c0a0c0a0a;
    encBuf[4871] = 256'h0b0a0b0a0a0a0a0a090001030505040403040403030403030303040201020108;
    encBuf[4872] = 256'h08090a0a0b0d0b0c0b0d0b0d0b0b0d0b0b0c0b0b0c0a0a0a0909090800010203;
    encBuf[4873] = 256'h0304040304030402030303040303040203020201010009090b0d0c0c0b0b0b0b;
    encBuf[4874] = 256'h0b0b0b0a0a0a0a0800000202020403020401010000090008080108090b0f0f0e;
    encBuf[4875] = 256'h0c0c0c0b0c0c0b0b0b0b0c0b0a0a090a09090800010102040303040403040304;
    encBuf[4876] = 256'h040202030202010200010009090c0c0b0f0b0c0c0b0b0c0b0a0a0b0a0a0a080a;
    encBuf[4877] = 256'h080808000302050403040502030402030202010200000009090a0d0c0b0d0c0b;
    encBuf[4878] = 256'h0b0d0b0b0c0a0b0b0a0c0a090a09000003060403060204030204020303030304;
    encBuf[4879] = 256'h030203030303020000090a0b0c0d0b0b0c0b0c0b0b0b0c0a0a0b0a0a0c0a0909;
    encBuf[4880] = 256'h08010101040305050304030203020100000a0a0d0d0c0c0b0d0a0c0a0a0b0a0a;
    encBuf[4881] = 256'h0a090909090a090a090a08010306050403050303040303030402010203020304;
    encBuf[4882] = 256'h0402040203050204030304040403050304040304030403030402030202020201;
    encBuf[4883] = 256'h010100080a0a0c0c0c0c0b0c0c0c0b0b0c0c0b0b0b0b0c0a0b0a090909000002;
    encBuf[4884] = 256'h030503050304030304030402030203020301020000090a0d0b0d0c0b0d0b0b0d;
    encBuf[4885] = 256'h0a0b0b0c0a0b0b0a0a0b0a090a08000102050404040304030403030303040203;
    encBuf[4886] = 256'h03020301010008090b0b0e0b0c0b0c0c0a0b0c0a0b0b0c0a0a0a090800010203;
    encBuf[4887] = 256'h060403050303050303030502030303030303020101080a0b0c0d0b0c0b0b0c0b;
    encBuf[4888] = 256'h0c0b0c0b0b0c0c0a0b0b0a0b0909080001030404030404020304020303030302;
    encBuf[4889] = 256'h0301010009090b0c0b0b0c0b0b0d0b0d0b0c0b0a0a0a09080000010101000001;
    encBuf[4890] = 256'h010306050403030202000a0c0d0d0b0d0b0b0b0c0c0a0c0b0b0c0b0b0c0a0a0a;
    encBuf[4891] = 256'h09080001010304030404030303040303030404030303030201010009090b0c0b;
    encBuf[4892] = 256'h0c0c0b0b0c0c0b0c0b0c0b0b0a09080802010304030402020202020203020101;
    encBuf[4893] = 256'h090b0e0c0d0b0d0b0c0a0c0b0b0d0b0c0c0a0c0a0a0a0a080001030404030403;
    encBuf[4894] = 256'h0303020403040503040402030303020201010008080a0a0c0b0d0c0b0d0a0b0c;
    encBuf[4895] = 256'h0a0a0a0a0a0a0a090a0908080801020405040404030402020302010202000108;
    encBuf[4896] = 256'h0a0b0c0d0c0b0c0d0b0b0d0a0a0b0a0a090a0909000808010002040405040305;
    encBuf[4897] = 256'h0203020201010808080a090a0a0a0a0b0a0b0e0b0b0d0a080802070404050304;
    encBuf[4898] = 256'h040403050304030305020303020302010101080809090c0b0e0b0d0b0c0b0c0b;
    encBuf[4899] = 256'h0b0b0c0b0a0b0b0b0b0a0b0a0909010205040503050304030303030304020201;
    encBuf[4900] = 256'h01010809090b0c0c0c0b0c0c0b0b0b0c0b0b0b0c0c0a0a0a0a09090801020503;
    encBuf[4901] = 256'h05030404020303040202020201010100080808090b0c0c0d0b0c0b0c0b0c0a0b;
    encBuf[4902] = 256'h0b0b0a0b090a0808000304050404030403030403030304030303040202020100;
    encBuf[4903] = 256'h0009090c0b0c0b0c0b0c0b0c0a0c0a0a0a0a0a0b0c0b0a0a0908080100080809;
    encBuf[4904] = 256'h0a0b0b0c0b0b0b0b090809090f0d0c0d0b0c0b0b0b0a0a0a0900020405030403;
    encBuf[4905] = 256'h0403050303040304020203030203020108080a0a0c0b0e0b0d0c0c0b0c0c0a0c;
    encBuf[4906] = 256'h0a0a0a0908080000090809080801020603050303030402020202020303040302;
    encBuf[4907] = 256'h02080b0d0d0d0b0c0b0b0b0b0a0a0a0800000000090a090b0903070505030304;
    encBuf[4908] = 256'h0202010101000808080a090a0c0d0c0c0d0c0b0c0b0a0b0a0a090a0908080000;
    encBuf[4909] = 256'h0101010404050305030304030304030402030102000100000008090a0c0d0b0d;
    encBuf[4910] = 256'h0c0b0b0b0a0908080808090a0a08000206040305030402020201020305050304;
    encBuf[4911] = 256'h02010108080a0b0a0b0c0a0a0a090909090b0d0c0c0b0b0a0a08080000020103;
    encBuf[4912] = 256'h05020402020202030604030403030302020108080b0c0b0c0b0c0c0c0d0b0d0a;
    encBuf[4913] = 256'h0b0a090801020404030402020202050404040404030304030403040304030402;
    encBuf[4914] = 256'h0201000009090a0a0a0b0b0c0b0d0c0b0d0c0b0b0b0c0a090a0a0a0a0a0a0a09;
    encBuf[4915] = 256'h08000304050403040402030402030303020301010808090a0b0c0c0c0c0b0d0a;
    encBuf[4916] = 256'h0b0b0a0b0a0b0b0b0d0a0b0a0908000203040503040303030303040403040202;
    encBuf[4917] = 256'h000009090b0c0c0c0c0b0b0c09090909080a0909000306050303010101000204;
    encBuf[4918] = 256'h0403040403040304030100000800000101090b0f0c0a0a0000020200090a0b0a;
    encBuf[4919] = 256'h08080100000202040402090b0f0d0b0b0b0b0c0c0b0b0b0b0b0c0b0e0c0b0b0a;
    encBuf[4920] = 256'h0a080801000008090a0a0901070604050402020101080000020203030108090a;
    encBuf[4921] = 256'h0b0a0b0c0d0c0c0b0c0b0a0c0a0b0b0a0909080b0c0e0b0b0a08000101010802;
    encBuf[4922] = 256'h040604030201000a0a0b0a0b0b0c0b0908010203010a0c0d0b09000304030201;
    encBuf[4923] = 256'h020307050302020008080103070404020200090b0c0b0b0a09090a0b0e0d0c0b;
    encBuf[4924] = 256'h0d0a0b0a09080101010108080a0b090802040503030402030304030302020202;
    encBuf[4925] = 256'h0504040200090c0d0b0b0b09000102030402030108080a080107050503040200;
    encBuf[4926] = 256'h000008080808080908090809080a0d0c0d0c0b0c0c0a0b090900020304020201;
    encBuf[4927] = 256'h00080800080000010307040403020008090d0b0d0c0b0b0b0b0c0a0a09090808;
    encBuf[4928] = 256'h00010102020108080a0b090005060403030202000202020402090c0f0d0c0b0b;
    encBuf[4929] = 256'h0b0900010504040303040404030504030304020303040203030302030108090a;
    encBuf[4930] = 256'h0d0b0c0c0c0b0c0b0c0b0c0a0b0a0b0b0b0b0a0b090908010205040404030304;
    encBuf[4931] = 256'h030403040203020202010009090b0d0c0b0c0c0b0b0c0b0b0b0c0a0a0a0a0a0a;
    encBuf[4932] = 256'h08000002020202020305050504030402020101080000000000080a0d0d0c0c0b;
    encBuf[4933] = 256'h0c0a0a0a09090a09090908000103040404030304040303040303030303030101;
    encBuf[4934] = 256'h010102030302000c0e0b0b0a08000108090a0902060504030203010203020108;
    encBuf[4935] = 256'h0a0b0c0a0a0c0e0d0d0c0b0b0b0a0c0c0b0d0b0a0a0909000008000001030405;
    encBuf[4936] = 256'h040304030403030303040202030202020101000808080b0d0e0c0c0c0b0b0b0b;
    encBuf[4937] = 256'h0b0b0c0b0c0a0b09090000010303040202000808080204040302080a0b0a0800;
    encBuf[4938] = 256'h02000c0f0e0b0d0a0b0909080102020102010002040505030302020102040305;
    encBuf[4939] = 256'h030202000909090b0c0c0d0c0b0c0a0a090909090809090a0a0a0a0909000304;
    encBuf[4940] = 256'h05030301010001050604040201080b0b0c0a0900080008090908080204030304;
    encBuf[4941] = 256'h010102080801020707060403020201000008000808090c0c0d0b0d0a0b0a0a09;
    encBuf[4942] = 256'h080008000909080102040301010008010405060404030403040302030100090b;
    encBuf[4943] = 256'h0d0b0c0a0a090a0c0b0d0b0c0b0a0a0a09090900000303030304030504040303;
    encBuf[4944] = 256'h0202010103030303010001020402080b0f0c0c090a09090b0c0c0a0802050503;
    encBuf[4945] = 256'h040203030505040305020303030403020401020001080009080b0b0e0b0c0b0b;
    encBuf[4946] = 256'h0c0a0b0c0b0c0b0b0b0b0b0b0a09080102040503030404030403020202020102;
    encBuf[4947] = 256'h0202010200090a0c0e0c0c0b0b0b0c0b0c0b0d0a0b0a08080001000201030404;
    encBuf[4948] = 256'h0402020000000102030201000800000203080e0f0d0d0a0b0a090809090a0909;
    encBuf[4949] = 256'h0801020304040304030503050302030202020303030201080a0d0c0c0c0c0b0a;
    encBuf[4950] = 256'h0b090a0808080808090002040603040303030403040201010101010101090b0f;
    encBuf[4951] = 256'h0d0b0c0c0c0b0c0b0b0c0a0b0b0a090a08000001020305030503040304030404;
    encBuf[4952] = 256'h03020201010001000000080a0b0d0b0b0a0b0b0d0b0d0b0b0c0b0c0a0b0a0909;
    encBuf[4953] = 256'h0908080001050504030201000809090a0b0d0c0c0c0a0b090909090a0a0c0b0c;
    encBuf[4954] = 256'h0a0a0b0a09080207050404020201010002030503030100080809080000080a0d;
    encBuf[4955] = 256'h0d0c0b0d0a0b0b0b090900000809090a090800020303050304030101080a0a0b;
    encBuf[4956] = 256'h0b0b0d0b0e0b0c0c0a0a0a0a0b0a0a090002030301090b080407070502020200;
    encBuf[4957] = 256'h0102020503040201010002010200090d0d0b0a0a090008090a0d0b0c0a080801;
    encBuf[4958] = 256'h0204020304030302010000080203050302080b0d0c0a0a09090b0e0b0c0b0a0a;
    encBuf[4959] = 256'h0b0b0b0b0804070404020108090a090b0900000203030404020201080c0d0d0c;
    encBuf[4960] = 256'h0a090908090b0d0d0b0b0b0a0b0a0b0c0c0a0b0a0a0c0b0b0a00050505050303;
    encBuf[4961] = 256'h0404030403030403040403030304020302020302010200090a0d0c0d0b0b0c0b;
    encBuf[4962] = 256'h0b0b0c0b0c0b0b0c0a0a0a080001020303030304030504040203030201020201;
    encBuf[4963] = 256'h0203020101080a0b0d0c0a0a0b0b0d0c0b0d0b0c0a0909080008000809090800;
    encBuf[4964] = 256'h03070503020208090b0c0a0b0b0d0d0b0c0b0a0a0908090b0c0b0c0908010303;
    encBuf[4965] = 256'h04020201030305030202020405040403020009090900030303090e0d0c0b0900;
    encBuf[4966] = 256'h010102020103060503050202010101010304030200080a0c0c0a0c0b0c0b0c0b;
    encBuf[4967] = 256'h0a0b0c0b0e0b0b0b0b0908080000000101030403050305030503040203020203;
    encBuf[4968] = 256'h0303020108090c0c0c0b0b0a0a09080000080a0b0d0b0c090808000100010201;
    encBuf[4969] = 256'h01010a0e0d0c0c0b0b0a0a0b0c0d0b0d0a0a0b0b0c0c0b0b0908020304020008;
    encBuf[4970] = 256'h08000307060303030303030402030100000800080009090b0d0c0c0b0c0b0b0b;
    encBuf[4971] = 256'h0c0a0b0c0b0b0c0b0b0a090002030304010809090901030403010a0c0d0b0b0a;
    encBuf[4972] = 256'h0d0c0d0b0c0a0800020402020202010203040404040403030402010101000101;
    encBuf[4973] = 256'h020101000809080000000c0f0f0c0c0a0a0a0908090808000305040202010001;
    encBuf[4974] = 256'h020204020108090a0909090a0b0d0b0b0a09090a0c0d0a0a0b0b0f0c0d0b0a08;
    encBuf[4975] = 256'h0204050402010008090909080809090808020303010a0f0c0b08010305020108;
    encBuf[4976] = 256'h080801030502080c0d0b0b090800000809090008010303070705030503030402;
    encBuf[4977] = 256'h03040204020303020303030403040304030304020100090a0b0c0b0c0b0e0b0b;
    encBuf[4978] = 256'h0c0a0a0909080b0b0d0b0a080203050203020203020301080b0a0a0006040302;
    encBuf[4979] = 256'h0809090a0901080a0b0f0c0b0b0b0c0c0c0c0b0c0a0a09080800010201020101;
    encBuf[4980] = 256'h010102040302000d0f0c0b0d0a0a08080008090b0d0b0c0a0908000102010202;
    encBuf[4981] = 256'h0102020404040304030205040305020201000808090808080908000104040301;
    encBuf[4982] = 256'h00090801050504020208080a0801030502010a0e0d0c0b0b0b0c0a0b0b0c0b0c;
    encBuf[4983] = 256'h0b0c0b0c0a0a0809000000080a0c0b0900040703040303010201010102010200;
    encBuf[4984] = 256'h0101030302010a0f0e0b0c0a09080008080b0a0b090800090a0d0c0a0a090a0d;
    encBuf[4985] = 256'h0d0c0b0b0a08000102030201080a0e0d0b0c0a0900020303020208080008090c;
    encBuf[4986] = 256'h0e0c0a09020604040200090b0c0b0808020404030304020108090a0b09010302;
    encBuf[4987] = 256'h000e0f0b0d0a0808000100080008010200080a0d0c0a090800080b0e0d0b0c0a;
    encBuf[4988] = 256'h0908080001020503040201080a0c0b0a000003020008000104060303000a0d0b;
    encBuf[4989] = 256'h0b09000201000b0b0a0805060302010000030605040202000808080800000008;
    encBuf[4990] = 256'h090b0b090800090c0e0c0c090a08090a0a090106070403040101080000020305;
    encBuf[4991] = 256'h02020000080908090b0d0a0b0a0909090c0d0d0b0b0909080801000205040404;
    encBuf[4992] = 256'h020201000800080800090a0c0c0b0a080104030301000a0c0c0d0b0c0b0b0a08;
    encBuf[4993] = 256'h01050504040303020302030304040202010101010103020200090a0a08030604;
    encBuf[4994] = 256'h0301090d0d0c0b0c0b0b0c090901040404020201080008010102020109090a00;
    encBuf[4995] = 256'h030604030100090a0c0b0b0e0b0b0b0802040603030203020201020201000009;
    encBuf[4996] = 256'h0b0a0d0a0a0909080b0c0b0d0c0a0a0a0a0a0d0d0d0d0c0b0a0a090000000101;
    encBuf[4997] = 256'h03030704040402020200080908000103030201010100080a0e0e0b0c0b0a0b0c;
    encBuf[4998] = 256'h0b0b0b0800010101000103060303010a0b0e0b0c0b0c0b090103040401080b0d;
    encBuf[4999] = 256'h0d0a0a0a080808090a0b0a00020602080b0f0d0a080103040202010102020200;
    encBuf[5000] = 256'h090c0b0a0104040301090d0d0b0b0a0a09080800020404050202010809090808;
    encBuf[5001] = 256'h08090b0b0007050303000a0c0b0c0a090a0b0a09010405030301080809000008;
    encBuf[5002] = 256'h0d0d0d0b090804040502020008090908010000090a0b0902050402080a0c0c0b;
    encBuf[5003] = 256'h0c0c0b0c0b0b080002020300080b0d0b0b090802040505040302020109090a0a;
    encBuf[5004] = 256'h0a0a0a0b0b0c0a09080808090d0c0b0a0801020304040505050202080a0c0c0b;
    encBuf[5005] = 256'h0a080102040203030303030300090c0b0b0a0800010000010303010c0f0f0b0b;
    encBuf[5006] = 256'h0a0a09080000000001020305030401000a0c0b0b08030706020208090a090003;
    encBuf[5007] = 256'h0402000b0c0a020705040201090a0b0c0b0b0d0b0c0b0a080204040302010800;
    encBuf[5008] = 256'h010504040200090b0c0a090008080a0c0b0a0801020201080004050603030303;
    encBuf[5009] = 256'h0303030302020009090a0c0b0c0c0a0a0a090802050704040303030201010008;
    encBuf[5010] = 256'h090b0d0d0b0d0a0a0a010203040100090a0b0808010101010505050403010009;
    encBuf[5011] = 256'h0b0d0a0a09080001020101010003050302000d0d0c0c0b0a0b0b0b0b0b0a0800;
    encBuf[5012] = 256'h030505030200090a0c0b0a0909090a0c0c0b0b090004060403030208090b0d0b;
    encBuf[5013] = 256'h090908000809090a0909000105060505040303020100090a090a0a090a0c0c0d;
    encBuf[5014] = 256'h0c0b0b0b09000104040402030202020008090c0b0c0b0b0b0e0b0c0b0a080002;
    encBuf[5015] = 256'h020304030303040204020201090d0d0b0b0a0a0a0a0d0b0b0a09010204050305;
    encBuf[5016] = 256'h03030202000101080a0f0c0b0a090808090b0b0804060303080a0a0a00020208;
    encBuf[5017] = 256'h0d0d0b0900010100090c0d0c0c0c0b0b0a08010203040303020108080a080207;
    encBuf[5018] = 256'h0402000a0b0d09080001010101030201080b0c0a09000009090803070502080b;
    encBuf[5019] = 256'h0c0c0a0a0b0d0c0b08000202080c0d0b0a010204030202020303030301080c0d;
    encBuf[5020] = 256'h0e0b0b0802050302080b0c09020504020101010405040202000000000000090b;
    encBuf[5021] = 256'h0c0c0a0a090001020303000b0d0c0a080102010808000202090e0f0c0b090003;
    encBuf[5022] = 256'h02020000010407050302020109090b0b0c0b0c0b0c0b0c0a0908010204030200;
    encBuf[5023] = 256'h08090a0b0c0c0c0a08030604030201080002050303000a0c0c0b0a0808020204;
    encBuf[5024] = 256'h0403030108090a0801030403040202020809080207060301080a0a0105060402;
    encBuf[5025] = 256'h0200000000080008010406050202090a0d0b0c0a090900010204020101020204;
    encBuf[5026] = 256'h0302000c0d0b0b09080808080102060302080a0b0c0a08080000080101090b0f;
    encBuf[5027] = 256'h0c0b080000080b0e0b0802040200090b0901060301090d0b0b0a080808090103;
    encBuf[5028] = 256'h070302000a0c0a080303030a0f0d0c0b090000010108080a0002060604020208;
    encBuf[5029] = 256'h0a0b0c0a090a0b0e0b0a010505030300080909080800090b0d0b0b0803050402;
    encBuf[5030] = 256'h01080a0b0b0a090800000103050402080c0f0c0b0908010301000a0b0a010305;
    encBuf[5031] = 256'h0300090a0901040402080a0c0b08010302080d0e0b0a000305030109090a0102;
    encBuf[5032] = 256'h04000c0e0c0a090802020202020203050201080b0f0c0c0b0b0a080001020101;
    encBuf[5033] = 256'h0203060404030108090b0b0b080103040400080b0d0b0c0a0b0d0b0c09080104;
    encBuf[5034] = 256'h0403030202030200090b0c0b0a0a0a0d0c0b0900010101080900020504020202;
    encBuf[5035] = 256'h030602000b0f0c0a09080100090a0b0a010305040304030201090a0a00050402;
    encBuf[5036] = 256'h000b0b0a010404000a0b0b010604010a0e0b0b08020403020008000808090b0e;
    encBuf[5037] = 256'h0b0c0a090800020202080b0d0a08020602000a0c090307050200090a0c090900;
    encBuf[5038] = 256'h0008090808010303030101000203040108090b0c0a0c0c0d0c0b0d0b0c0b0a08;
    encBuf[5039] = 256'h0204030403020403040202080a0b0a080303010c0e0c09000203020108080405;
    encBuf[5040] = 256'h040301080a090808080b0c0a090000090f0d0c0a090001020203050404030201;
    encBuf[5041] = 256'h090a0a0a0800030404020201000001010201090d0d0c0a0a0a0a090802060503;
    encBuf[5042] = 256'h03010809090000090e0f0c0b090802020301080800020405020101000800080a;
    encBuf[5043] = 256'h0d0c0b0a0801020100080801050404010108090a0c0d0c0c0a09000203040202;
    encBuf[5044] = 256'h0000080c0c0c0c0a0908000808080102050301090a0b0a010505020200000103;
    encBuf[5045] = 256'h050303080b0f0b0b0900030203020204040401080d0e0c0b0b0800020301080a;
    encBuf[5046] = 256'h0b0a01030501090c0d0a080202030200010307030100090b0a0800000a0d0c0b;
    encBuf[5047] = 256'h0a0900010203070304020809090900000a0f0d0b0a080808090b0a0207060402;
    encBuf[5048] = 256'h02000009080a0a0a0a0a080008080000030502090e0e0b0b0900010008000004;
    encBuf[5049] = 256'h06030401080a090a0808090b0d0d0a09000205030302080a0b0a0a09080a0d0d;
    encBuf[5050] = 256'h0b09010504020008090002050402000a0d0a0a080101080c0c0c090802030300;
    encBuf[5051] = 256'h090a0a00040402000a0d0b0b0900010101000801030704030200090909080101;
    encBuf[5052] = 256'h00090901060503010a0e0d0a0a080002020203040503030200090b0b0c0b0d0d;
    encBuf[5053] = 256'h0b0a09010404040101080008000008090b0a080004040503030201090a0c0b0b;
    encBuf[5054] = 256'h0a0a0b0a0a01060402000b0f0c0a09010204020200000a090a00010404030009;
    encBuf[5055] = 256'h0a0a08020302080d0c0a0001010a0f0d0b0901040201090d0b0b000305040200;
    encBuf[5056] = 256'h090b0b0900020503010008000304030a0f0f0b0a0801030301080a0a08050504;
    encBuf[5057] = 256'h0100090a0a090102020100010307040202000b0c0d0a0a090809080a0a090003;
    encBuf[5058] = 256'h06030201080900020303000b0d0a0004040400090a0c09000102020307050403;
    encBuf[5059] = 256'h02000a0c0b0b0b0b0c0b0a09000403030201010102080a0e0b0a000305020109;
    encBuf[5060] = 256'h0b0c0b0c0d0b0b0a00040403030304040303080b0f0c0b090a08090808020203;
    encBuf[5061] = 256'h01090b0901060403010a0c0c0909000101010202010a0f0c0c09000103030302;
    encBuf[5062] = 256'h02030201080d0d0b0900020201080a0b0a0b0a0b0c0c0b0b0b09090001020404;
    encBuf[5063] = 256'h0404040202080b0c0c0a0a09090a0b080407060301090d0c0a09010404020108;
    encBuf[5064] = 256'h0909090000000000020303080e0e0c0a0801040202000a0e0b0b0a0800010203;
    encBuf[5065] = 256'h0202020108090a0a08080a0d0f0b0a08020604040201010108090a0c0b0a0900;
    encBuf[5066] = 256'h0002030202080b0f0c0a0a0a090a0a090207060301080c0c0b0a090900080103;
    encBuf[5067] = 256'h07030402010808080000080a0d0c0a0900020302000008090c0d0d0a0a010306;
    encBuf[5068] = 256'h030201000108090c0e0b0b0900020100090b0802070603010108090a09090800;
    encBuf[5069] = 256'h0108080b0c0b08020402000a0b0903070301080a09010504010a0e0d0a0a0801;
    encBuf[5070] = 256'h0303030302000a0b0c0b080801000808030706040200090c0c0b0a0909090b0b;
    encBuf[5071] = 256'h0901070503040100080809080100000008000307030401090a0c0b0a0a0c0d0c;
    encBuf[5072] = 256'h0a0a0001030301000002020402080a0d0a0802040302090a090005040302080b;
    encBuf[5073] = 256'h0a080406040201090a0a0b080002080a0e0c0b090000010a0b0d0a0104040402;
    encBuf[5074] = 256'h010001000100000008090b0f0c0c0a0802040402010101010201090d0d0b0a08;
    encBuf[5075] = 256'h010301000a0a0a0104030201080b0c0c0c0a0a00030402030101020200090e0c;
    encBuf[5076] = 256'h0b0a0a0a0d0e0c0b0a080203050302030304040302000a0e0c0c0a0a00010303;
    encBuf[5077] = 256'h0201080808010201090f0d0c0c0a0a09090908020405050203010008090a0908;
    encBuf[5078] = 256'h09090a0b0a0802050402010909090002030108090a080202090f0f0f0a0a0801;
    encBuf[5079] = 256'h02030200000909080000090b0f0b0a0001050402030101020100080b0d0c0908;
    encBuf[5080] = 256'h02030200090c0b0a000304030301090b0d0b090900090e0e0c0b0b0a0b0b0c0a;
    encBuf[5081] = 256'h090205050303010100000200000b0d0c0b08000303010a0c0a0004060302000b;
    encBuf[5082] = 256'h0d0a08010204020100000003040402080d0e0d0b0b0a09080800010206040403;
    encBuf[5083] = 256'h020100080000080c0c0d0b0a080203050101090a090900030305020302020108;
    encBuf[5084] = 256'h0b0e0c0b0a0900020101080a0b0b0b0a0a0a0b0b0c0b08050706030303020100;
    encBuf[5085] = 256'h020201090e0e0c0b0b0909010103040301010009090b0a0a0a00020605030200;
    encBuf[5086] = 256'h090a0b0a0a0a0c0d0d0a0a08000102040504040200080a0a0a0001000a0d0c0a;
    encBuf[5087] = 256'h0a000000010204040401080a0b090206030308090b0a0101010b0f0e0b0a0808;
    encBuf[5088] = 256'h020202040201010103060404020100000800090b0f0d0b0a0901010200080809;
    encBuf[5089] = 256'h080203060304020108080a0a0b0c0b0d0a0a0802040301000808010102000104;
    encBuf[5090] = 256'h07070302010a0b0d090800020100090809010108090e0c0a0a08000000090b0b;
    encBuf[5091] = 256'h08030707020108090a0a09080000080000020201010809000205050402020001;
    encBuf[5092] = 256'h0002040302090f0e0c0b0b090908000800080000010203050404030304020009;
    encBuf[5093] = 256'h0b0d0a0a0800000b0f0d0c0a0a08010101000002050504020300080a090a0808;
    encBuf[5094] = 256'h08090a090a0800080b0f0f0c0b0b090803050304020100080a0b0c0a0a000304;
    encBuf[5095] = 256'h040201010000000a0c0e0b0c0a090001030503020108090a0b0b0b0b0d0b0a09;
    encBuf[5096] = 256'h0205030301000a09090908080a0b0a00060605030402080a0e0c0b0a0a0a0a0b;
    encBuf[5097] = 256'h0a0a000505040302010205030402000a0c0b0a0808080c0d0b0b090002030304;
    encBuf[5098] = 256'h03030402010000080a0c0e0c0b0900020303000a0908030502000b0d0a000001;
    encBuf[5099] = 256'h0a0d0d0a00020503030202010200090a0c090808090c0c0a08050403010a0b0b;
    encBuf[5100] = 256'h09010401080b0a090102080e0e0b0b0808000a0d0c0a09020304030304040202;
    encBuf[5101] = 256'h02010204050301000a0e0b0b0c0b0b0d0b0b0a00020403030403030502020009;
    encBuf[5102] = 256'h0c0c0b0b0b09080101020301010204050403020109090a090908090b0e0b0a08;
    encBuf[5103] = 256'h02050302010001030502010a0d0c0a0803040301080b0c0b0b0b0d0d0c0b0c0b;
    encBuf[5104] = 256'h0a0800020505040303020000090a0a0b0c0a0a0800030404040304030302080b;
    encBuf[5105] = 256'h0e0b0b09080009090b0c09080202080a0e0a0903050303080a0c0b0a09080a0d;
    encBuf[5106] = 256'h0c0b09040705030201090b0b0b0a000100080b0b0903070703020109090b0908;
    encBuf[5107] = 256'h0000090c0c0a08000302020809000103040100090a0a0a080105040302090f0c;
    encBuf[5108] = 256'h0a0902050302000909010403020a0f0b0b080001080a0b0a020502080d0d0b08;
    encBuf[5109] = 256'h020304020102050503000a0d0d0b090900010008080008010202030503050202;
    encBuf[5110] = 256'h02010000090b0c0d0c0c0b0b0a09080103030202010403060202080a0d0b0b09;
    encBuf[5111] = 256'h09090b0d0c0a0901040504030200090b0d0b0909010203030201020000080809;
    encBuf[5112] = 256'h00020404030200090d0b0d0b0b0a000307060304030201090c0c0c0c0b0b0c0a;
    encBuf[5113] = 256'h0a09000204040402020302030201090d0c0d0a0a0a0800000103030302000909;
    encBuf[5114] = 256'h08010100090d0b0803060402080b0d0c0a090909080801030403020109090a0a;
    encBuf[5115] = 256'h000204050302000a0b0b080203000f0f0d0b0908020304030403040302000b0e;
    encBuf[5116] = 256'h0b0c0a0908010204030301080a0b0c0a090a08080103040301090a0c0d0c0c0b;
    encBuf[5117] = 256'h0b0802040502010809080204030200090a0804050401000a0a0a010202000c0e;
    encBuf[5118] = 256'h0c0b0b09080102020200010205050300090d0b0b08010401000a0a0c090a0b0c;
    encBuf[5119] = 256'h0d0b0a090802040604040202000009080808090b0d0a0002060300080b0b0a00;
    encBuf[5120] = 256'h0302080e0d0a000206020208090b0a09090b0e0b0b0801060403020201010000;
    encBuf[5121] = 256'h0808000101020300080a0b0d0c0c0d0c0c0b0a08000303020200000204040302;
    encBuf[5122] = 256'h090c0d0b0c0a0a0a0a08020305040302030202020100090d0b0c090003040302;
    encBuf[5123] = 256'h080b0f0c0b090900010203050305030100090b0b0a090808090c0b0b0b0c0d0c;
    encBuf[5124] = 256'h0b0a0908080a0d0a0903070502020000010306030200090c0b0a090808000809;
    encBuf[5125] = 256'h0809090a0d0c0c0c0a0900030603020200080a0a0a0c0c0b0b08010604040301;
    encBuf[5126] = 256'h01000001030302080c0d0b0b08010102090d0c0c0a0908080008010307060202;
    encBuf[5127] = 256'h08080a0a0908090a0e0c0b0b0800030304010108080909000102040200080901;
    encBuf[5128] = 256'h03060301090a0b0901030201080804070303080c0c0b0b09090a0c0d0a0a0909;
    encBuf[5129] = 256'h08090a0a0d0b0c0901060604040202020200080b0f0d0b0a0908010101080800;
    encBuf[5130] = 256'h04050302000a0b0b0a000102010008010103050202080c0f0c0c0b0900010201;
    encBuf[5131] = 256'h01010104040202080a0b0a000101090a0c000407040308090c0b0a0003030301;
    encBuf[5132] = 256'h090a0a090a0d0d0d0c0a0a08010204030302010000010100090b0c0901070503;
    encBuf[5133] = 256'h030108090b0b0c0b0c0c0c0c0a09080002020403040302020000080101010108;
    encBuf[5134] = 256'h09080002010b0f0f0c0a0908010202020202030302080d0f0c0b0b0900010404;
    encBuf[5135] = 256'h0202020102020101080d0d0b0c09080102000809090001020301080801030403;
    encBuf[5136] = 256'h010a0e0a0a00030502000a0d0b080307060100090c0a090101080a0c0c090105;
    encBuf[5137] = 256'h03030009090802040401080b0c0c0b0b0d0a0908030504030108090909090a0b;
    encBuf[5138] = 256'h0d0b080207050303020009080a0c0c0c0b0a0800010000080900010503040301;
    encBuf[5139] = 256'h010800090a0a0c0b0b0c0a090002040301090b0c090203040109080106040309;
    encBuf[5140] = 256'h0f0d0b0a00010201080a0a010604030200090a08010304020201000000000100;
    encBuf[5141] = 256'h0a0e0f0c0d0b0a0a080003040404020200000a0a0b0a09000304030301090b0e;
    encBuf[5142] = 256'h0c0b0a090102020100090800030502080a0d0b0b09080001030706020208090c;
    encBuf[5143] = 256'h0b0a09090a0c0a0802060403020202020301090c0e0c0b0b0b09010307040302;
    encBuf[5144] = 256'h0108090a0b0b0c0c0c0b090802040503020108090a0b0a0a0a0b0d0d0b0b0802;
    encBuf[5145] = 256'h0604040201000808000101090a0d0b0908000101080a09080204040202020009;
    encBuf[5146] = 256'h0b0d0c0a09080002030306030301080d0e0c0b0b090801020304020303030304;
    encBuf[5147] = 256'h0202010a0f0c0c0a0901010301000a0a0a0901040404040200090b0d0b090908;
    encBuf[5148] = 256'h0a0b0f0a090004030401080a0a08020303000a0b0a0207050302000008010108;
    encBuf[5149] = 256'h090d0c0b0c0a090900020504030301010101000b0f0f0b0b0908010302020102;
    encBuf[5150] = 256'h010100080b0b0c09080002020504060304020200080a0a0c0a0b0b0c0b0d0b0b;
    encBuf[5151] = 256'h09010405030301090b0b0a00020404020100080a0a0b0b0c0c0c0a0b08010503;
    encBuf[5152] = 256'h0302090a0b090204010a0f0c0a00040603020108090908090a0d0c0a0a000101;
    encBuf[5153] = 256'h000a0a0b0802060301080b0e0c0b090002040402010100010008090a0a080306;
    encBuf[5154] = 256'h03000b0d0c090801010a0b0b080407040100080a00020502010b0e0c0b090102;
    encBuf[5155] = 256'h03030100090b0b0c0b0a0a0a0a090805060504020200000800000a0c0c0b0900;
    encBuf[5156] = 256'h0202080c0e0b0a0801040503040201000a0b0c0b0b0909000809000000020202;
    encBuf[5157] = 256'h010305040301090d0c0b0a08090a0a0904070702020100090a0a0b0c0c0b0b09;
    encBuf[5158] = 256'h000204040303020100080b0a0a0800080a0e0c0a090203030208090007040401;
    encBuf[5159] = 256'h090c0d0a09000203020102010101080c0c0b090001000c0e0b0a010405030201;
    encBuf[5160] = 256'h01010000080a0c0c0b0c0a0a080004040301000a090802060301080a0c0b0b0a;
    encBuf[5161] = 256'h0a0c0c0b09020505020208090a09080205030301090d0c0c0a09000201010909;
    encBuf[5162] = 256'h0b0a0a090a090006070403030200080a0a0b0c0c0b0b0a080000020100010203;
    encBuf[5163] = 256'h060302000c0f0c0b0909010102000808030705030200090c0d0a0a0900010203;
    encBuf[5164] = 256'h050203030201090c0c0b0b080002010009090105050402000b0e0b0b0a000205;
    encBuf[5165] = 256'h020300000a0a0b09080102000b0f0c0a08010503040203040303000b0f0c0b0a;
    encBuf[5166] = 256'h090808090b0a08020405030101000002030403030208090d0c0d0b0b0b0a0800;
    encBuf[5167] = 256'h0307050302010a0c0d0a0a00000102010202030401000a0c0b0b0a0a0a090908;
    encBuf[5168] = 256'h0900000206050302080c0d0b0a0800080b0e0c0b080205040303010100010201;
    encBuf[5169] = 256'h00080c0c0c0b0a0a0900000103030503030300080b0c0b0c090a090a0a090006;
    encBuf[5170] = 256'h0605030401000a0d0c0b0a09080000010203050304020201020100090c0d0c0b;
    encBuf[5171] = 256'h0a0a0a09090909000103040304030201080b0a00040603000a0f0c0a09080000;
    encBuf[5172] = 256'h0809080407040301080a0c0a09000101080800020307020200090b0c0a0a0800;
    encBuf[5173] = 256'h08080a0c0b0900040401090c0b0802060402000a0a0a01020501080b0d0c0908;
    encBuf[5174] = 256'h00010809090802060402000a0c0c0a0102050301000908000200080d0d0b0a01;
    encBuf[5175] = 256'h04040201090909000202080a0f0b0b0a09000104050403030301080a0b0f0b0c;
    encBuf[5176] = 256'h0a0a09000203030202000008090b0d0c0b0901030404010008090808080a0d0d;
    encBuf[5177] = 256'h0b0c0a08020504030200080a0a0a08000101020306040302000b0f0d0b0a0b0a;
    encBuf[5178] = 256'h0808010206040403040100090a0b0b0c0a0b0a0a08020704030201080a0b0909;
    encBuf[5179] = 256'h0008090b0c0a0802040201090a0a0803050301090c0c0c0a0a0a0a0a0b0b0908;
    encBuf[5180] = 256'h01030504040303030503040201080a0b0b0b090808090b090107060503030108;
    encBuf[5181] = 256'h0b0f0b0d0a0a090800020403050302000a0c0b0c0901020303020009090b0b0b;
    encBuf[5182] = 256'h0c0c0a0a090a0a080106050403030300090c0d0c0b0a0103050403010008090a;
    encBuf[5183] = 256'h0b0d0b0c0a09000203040200080a080104060301010908080001000a0e0c0a09;
    encBuf[5184] = 256'h0003030208080803070303080c0d0c0b0a09080800010304030200090a0b0908;
    encBuf[5185] = 256'h08090c0c0a0105050302080a0a09010301080b0d0901040402000c0c0c0b0a0a;
    encBuf[5186] = 256'h0801030504030201020101080d0f0c0a0a00030303010008000203000c0f0c0b;
    encBuf[5187] = 256'h090002030402020303030301080c0d0c0b0c0a090803040301080c0b0b090203;
    encBuf[5188] = 256'h0401080b0b0b0002040201000901040302090f0c090004050202090a0c0b0a09;
    encBuf[5189] = 256'h0a0a0a080407070303030108090a0b0e0c0b0c0b090001020200000801040404;
    encBuf[5190] = 256'h020008090800030303000a0b0d0c0a0b0c0b0a0a0a0909080106060304010008;
    encBuf[5191] = 256'h08080100080b0f0a0a0001020108090900010201000003060402090e0d0b0a08;
    encBuf[5192] = 256'h00020108080103070503030200090a0b0c0b0909080809090b0c0a0801040403;
    encBuf[5193] = 256'h04020100080b0c0c0c0b0b0a0a0902040704030303020100080a0c0b0c090808;
    encBuf[5194] = 256'h080a0e0c0d0a0900010305030202010008000900080808090a0a0b09090a0d0d;
    encBuf[5195] = 256'h0d0c0b0a0a080802050504030403020108080b0c0c0a0909090a0b0e0b080205;
    encBuf[5196] = 256'h05020100090808020301090c0d0b0b0b0c0b0d0a080206040202010000010102;
    encBuf[5197] = 256'h080a0e0c0a0a08080102010201020000090b0b0d0a0a09030605040201080a09;
    encBuf[5198] = 256'h08000200090e0d0b0b09000101010101010405030301000909090101000a0c0d;
    encBuf[5199] = 256'h0a08020302090d0e0b0a000103040200080a0b0a0802040201090a0803070403;
    encBuf[5200] = 256'h02080a09090a0a0f0d0c0a09010202020008080207030300090d0b0a00020403;
    encBuf[5201] = 256'h030008090a090808080b0d0c0a080800090e0d0b0900030402080a0a00050604;
    encBuf[5202] = 256'h0402010009090b0a0b090a09090a0902040502090c0e0b0a0802030200090908;
    encBuf[5203] = 256'h040604040200080a0c0b0b0a00000108090a000306040200090c0b0a09000809;
    encBuf[5204] = 256'h09090105030401000909090800010406040301080c0c0b08010201080d0d0c0b;
    encBuf[5205] = 256'h0a09010304040302020201080a0b0e0a090900080800000202080e0e0b0b0901;
    encBuf[5206] = 256'h0202000000030603030200080002030100090b0b0e0d0d0b0b0901040301080b;
    encBuf[5207] = 256'h09030706030100090a090008090a0d0b0a0a0800020405040303000009080808;
    encBuf[5208] = 256'h090c0b0c0b0b0d0d0c0b0908010201020505060303010809090800090c0e0d0a;
    encBuf[5209] = 256'h090001030008090a0801040201090a0a00020301090d0a000407040203010200;
    encBuf[5210] = 256'h080b0d0e0b0b0b0a09090001030505030302010100080a0a0d0b0a0b09090909;
    encBuf[5211] = 256'h010206030301090a0b0b0a0a0d0e0c0b0802050403030100010102000a0e0d0b;
    encBuf[5212] = 256'h0b090909000002050604020300080a0b0c0b0a0a0a0908000203050303020201;
    encBuf[5213] = 256'h0000080b0c0c0b0b080103050302000000030403010b0f0f0b0a0a0808080102;
    encBuf[5214] = 256'h04050403030008090a0c0c0c0c0b0a090002020203030305030301000a0b0b09;
    encBuf[5215] = 256'h01020302090d0d0c09080102080c0f0c0b080205030301080900030403080d0c;
    encBuf[5216] = 256'h0c0a00010102080a0b0900030504020201000808090b0e0c0c0a090800020201;
    encBuf[5217] = 256'h0000020505040202090a0b0c0a090a0b0c0a000207030302080b0c0b0a0a0808;
    encBuf[5218] = 256'h090a0801040603030208000802040302000a0b0b00040403080e0e0c0b0b0908;
    encBuf[5219] = 256'h08010101000203070404030301090b0c0b0a0908090b0d0c0a09000202030203;
    encBuf[5220] = 256'h04050301080b0d0c09000101080b0d0b0801040503020100000000090b0d0c0a;
    encBuf[5221] = 256'h09010403040108090c0b0b0a09090a090802060504020201000808010101000b;
    encBuf[5222] = 256'h0d0e0b0b090800010009080002050402000a0a080206050301090b0d0b0a0908;
    encBuf[5223] = 256'h00000009090a090a090a0b0d0a090407060303020008090008000a0e0d0b0b09;
    encBuf[5224] = 256'h000304020100090000020200090c0b0b08030304080b0f0c0a08000202010001;
    encBuf[5225] = 256'h060704030301080c0c0c0a0b0b0a0909000104030304040203020208090b0b0b;
    encBuf[5226] = 256'h0a0a0b0b0a00020302090f0b090307060200090b0b080202000b0f0d09000403;
    encBuf[5227] = 256'h040100090908000008090a0b0900030301090d0d0b0a0801020301090b0d0901;
    encBuf[5228] = 256'h05050200090b0c0801030401090b0a0908000a0e0d0b09000305040302010009;
    encBuf[5229] = 256'h0c0d0c0b0a0908010101030503030301090a0b0b0b0c0c0b0a01040503030008;
    encBuf[5230] = 256'h080808080b0f0f0b0b0a0003050503030200090a0c0a0b0a0b0a090902040503;
    encBuf[5231] = 256'h0201000103060302090c0d0b0b0800020108080a090003040302000000040503;
    encBuf[5232] = 256'h01080d0c0a090001020200000204040302080d0e0c0a09080103020200010404;
    encBuf[5233] = 256'h02010b0f0e0a0a080100000000010405030300090a0a080000000a0a09010303;
    encBuf[5234] = 256'h090f0e0c0b0a090900030504040200000908080008090c0b09010403020b0f0b;
    encBuf[5235] = 256'h0c080001020808090004040401090c0c0b090003030302010001020403000c0e;
    encBuf[5236] = 256'h0c0b09080800080a080004050201090c0a08020503020009090103050301090c;
    encBuf[5237] = 256'h0d0c0b0b0b0a0800020303050304040302010a0c0d0a0b0b0a0b0a0902060503;
    encBuf[5238] = 256'h0201080800020202090c0f0b0c09080001010302020101080908080204020209;
    encBuf[5239] = 256'h0b0e0b0b0a09080908000307040403020200010008080c0e0c0c090802040303;
    encBuf[5240] = 256'h00000a090a0b0b0e0b0a0802060403020808090a080801010200090b0e0c0b0a;
    encBuf[5241] = 256'h08000101020504050302000c0d0b0a0002040301080a0b0b0a0a090c0c0a0901;
    encBuf[5242] = 256'h0704030201080a09080800090a0c0c0a080801040404040200090d0d0b0b0b0a;
    encBuf[5243] = 256'h090800030505030302080a0b0b0a0901020403040200080a0d0c0d0c0b0b0a08;
    encBuf[5244] = 256'h020504030201080909080808080a09090004060503030300090d0c0c0b0a0a0a;
    encBuf[5245] = 256'h0908010306040302010008090909090a0a08030504020109090c0a0c0b0c0b0a;
    encBuf[5246] = 256'h08030403010809000506040301080b0b0c0a0c0b0b0a00070504020100090b0a;
    encBuf[5247] = 256'h0b0b0b0b0b0a0902060402020108080101030301080c0c0b080002000a0d0d0b;
    encBuf[5248] = 256'h0900020302080a0b0a020705030108090b0909000108090801050602010b0f0d;
    encBuf[5249] = 256'h0b0a0800010102020304040301090a0c0b0a090800080001020403040101080b;
    encBuf[5250] = 256'h0c0d0b0c090a09090a08020605050303020108090d0b0d0c0a09000001020102;
    encBuf[5251] = 256'h0203040201090c0c0b0b09000102030504030201090c0c0c0a0801020302000a;
    encBuf[5252] = 256'h0d0a090900090b0c09020606030202000008090b0d0d0b0a0900030403020201;
    encBuf[5253] = 256'h0008080a0b0b090005050201000a0a0b0b0b0c0d0c0c0b0a0800030505030402;
    encBuf[5254] = 256'h03020100080a0a0b0b0c0c0c0a0b090801010100000205040402080a0c0c0a09;
    encBuf[5255] = 256'h08000201020403030301000909010302080e0f0b0b0900000008090802040302;
    encBuf[5256] = 256'h0a0c0b0900020a0f0f0b0a0804040402020203030301090f0c0c0a0909080808;
    encBuf[5257] = 256'h0001020100090c0a0900050404030403030301080b0d0c0a0b090b0b0c0b0c0a;
    encBuf[5258] = 256'h090808010406050304030108090a09080800090b0d0d0a0a0808000100010103;
    encBuf[5259] = 256'h03040302030203030302090d0f0c0c0a0a000203030301080a0d0c0b0a0a0104;
    encBuf[5260] = 256'h0504030302010108090a0b0c0b0b0b0d0b0d0b0908010100090a010606040302;
    encBuf[5261] = 256'h010808080100080b0d0c0b0a0a09090a0908020604020200090c0c0b09080306;
    encBuf[5262] = 256'h040202080a0a0b080808090a0d0a090003040201080800020403010a0d0c0902;
    encBuf[5263] = 256'h060403000b0e0d0b0a0908010304030503030100090c0b0b090900080a0b0c0b;
    encBuf[5264] = 256'h0a0002040303020404040302000a0c0c0a09080100000809000104050202080a;
    encBuf[5265] = 256'h0c0b0a09090008090a0b090205060303030203050403010b0f0c0a0900020108;
    encBuf[5266] = 256'h0c0c0a09010304020008080800010001020405030400080a0b0a0b0a0d0e0b0d;
    encBuf[5267] = 256'h0a0a0808000102060305020200090908080000000a0b0e0b0b0a080001020100;
    encBuf[5268] = 256'h090909090b0f0c0c0900050504020201010000000a0c0e0b0b0b090800030404;
    encBuf[5269] = 256'h0202080b0c0b0a0900000800020706030301090a0b0b09090a0c0b0b08010303;
    encBuf[5270] = 256'h080a0c0a0901030604040303020101010303030a0f0f0d0b0909000002020305;
    encBuf[5271] = 256'h03020208090b0d0a0a09090800010101000802040604030200080a0c0c0b0c0a;
    encBuf[5272] = 256'h090204050301080a0c0a0901040202080a0c0a0a09090c0c0a0904060302080c;
    encBuf[5273] = 256'h0d0a00030703020108090809080b0c0d0b0b080104030302080a0a0908000000;
    encBuf[5274] = 256'h090b0a000407040301080a0b0a090001090c0c0a080204030100090a0a0b0c0c;
    encBuf[5275] = 256'h0b0a08040603030301000a0d0d0b0c09010202020809000207030300090a0b00;
    encBuf[5276] = 256'h00080c0e0c0a00020402000b0c0c0a090801010205040403030100080a0d0c0c;
    encBuf[5277] = 256'h0b0a09000102020503060302010a0c0e0b0a090800000101030405030200090b;
    encBuf[5278] = 256'h0b0b0b080908090b090004060401080b0e0a0801040302010808010102000d0d;
    encBuf[5279] = 256'h0d0a0a000102020108010205040202080b0b0c0908000001090a0b0d0b0b0c0b;
    encBuf[5280] = 256'h0c0a0902050604030202010100000000080c0d0d0c0a0a080002020100000900;
    encBuf[5281] = 256'h000000000808010406030403010008090800080b0f0e0b0b0908000201080908;
    encBuf[5282] = 256'h010307020208090909080101080a09000407030208090b0b090000010909090a;
    encBuf[5283] = 256'h080002040402010d0f0b0b090002000b0e0b0005050400080c0a090003040201;
    encBuf[5284] = 256'h080801020302090d0d0b0c0b0a0b0a080205040302040305030201090b0a0a00;
    encBuf[5285] = 256'h090c0f0e0b0a0a000102030202030304020108090a08080800090a0c0d0c0b0a;
    encBuf[5286] = 256'h010504040100090a0908090b0f0c0b0802070403020100080800090b0d0d0c0a;
    encBuf[5287] = 256'h0a09080000020204040303030201000a0d0b0b0b0a0808080801020403030009;
    encBuf[5288] = 256'h0b0a09010108090a080407040300090a0b080103020a0d0c0a000302080f0e0b;
    encBuf[5289] = 256'h0b09010306020100090a09080002020008090a00020502000b0b080707040301;
    encBuf[5290] = 256'h080a0b0b0a0800090d0c0b09010203080b0e0a09010202080b0a000707040201;
    encBuf[5291] = 256'h08090b0c0a0a090909090801020505030201080a0a0a0a0808090a0b00050705;
    encBuf[5292] = 256'h030100090b0b0b0a090a0c0b0c0a090001020204020302020000090b0e0a0a00;
    encBuf[5293] = 256'h04050402000a0b0c08000202080a0b0806070304010008080000080b0e0c0a0a;
    encBuf[5294] = 256'h080008090b0e0b0908020305030202020203020302000a0e0d0c0b0b09090000;
    encBuf[5295] = 256'h03030503030100090a000305040200000001030301090c0c0b0a0c0c0f0c0c0a;
    encBuf[5296] = 256'h0b090802040402020108080801000200080909010202080f0d0c0a0802030301;
    encBuf[5297] = 256'h0809080406050302010008090a090a0b0b0d0c0b0b0a09080809090b09010505;
    encBuf[5298] = 256'h030301090a0a090900090b0e0d0b0a02070503030100090908080008090a0a00;
    encBuf[5299] = 256'h0407040201080b0b0a0a08090a0c0c0b090000000a0d0c0b0900020303030103;
    encBuf[5300] = 256'h04040401000b0d0b0b08000008090b0801070703040402020102010201080c0e;
    encBuf[5301] = 256'h0c0b0b0a0909090c0a0a000405040201080908090808090b0c0c0b0a09000104;
    encBuf[5302] = 256'h03030201020405040303010808080000090c0d0c0a000205030100090a0a0a0a;
    encBuf[5303] = 256'h0a0d0b0a0902040401090d0e0b0b0a0900000809090802070504030202000000;
    encBuf[5304] = 256'h0008090b0d0b0c090003040302090a0d0a000206020208090a09000101090c0e;
    encBuf[5305] = 256'h0b0a090809090d0c0b0b09020405030100090a08010305030301020403050201;
    encBuf[5306] = 256'h090b0d0a0a080009090a0a00020402000a090003050401000b0e0c0c0c0b0b0a;
    encBuf[5307] = 256'h0a080809080800030504040302030304030302090b0d0a0003050301000a0a08;
    encBuf[5308] = 256'h010203010b0e0c0c090801040303000a0d0d0b0d0a0c0b0c0a0a000105030502;
    encBuf[5309] = 256'h020100010808080a0a0a0a090a0909000003040405040405020300080a0a0901;
    encBuf[5310] = 256'h0202010a0e0d0b0c0c0a0a090909080009080900020405030302020202020009;
    encBuf[5311] = 256'h0c0b0a02060402010a0d0a0a0002030301010102050503030200080b0c0a0901;
    encBuf[5312] = 256'h01010a0f0e0c0c0b0b0b0b0a0a09000405040303020102030202090d0d0d0a0a;
    encBuf[5313] = 256'h08010205030303030201080a0b0b0a08010201080c0c0c0a0b090b0b0d0c0a0b;
    encBuf[5314] = 256'h0a0a0a090001030503030108080900050604040200090b0e0a09010306020202;
    encBuf[5315] = 256'h00000100000809090a090a0c0c0b0b09010303000c0f0c0b0b0a090900010203;
    encBuf[5316] = 256'h040300090c0b0a0207050302000b0e0b0b080204030201080800030604020201;
    encBuf[5317] = 256'h01020302080c0e0d0b0b090a09090a0a09090203050403030401000a0d0c0b0b;
    encBuf[5318] = 256'h0808010100000800010304030403070305030101080a0a0909090a0b0d0b0c0a;
    encBuf[5319] = 256'h0a0808010306030300090d0c0b090800000101020102080a0f0d0b0b0c0a0a09;
    encBuf[5320] = 256'h08010307050304030302000009090a0908000800080a0a0d0b0c0b0a0a0a0909;
    encBuf[5321] = 256'h0b0c0d0c09080305050201080909090008080a0e0b0c0a090808010205050304;
    encBuf[5322] = 256'h0304020201010800000101000e0e0d0b0a0801020301090a0b09010304010109;
    encBuf[5323] = 256'h090909090a0d0b0c0a000205040201080b0d0b08020505020108090b0a000104;
    encBuf[5324] = 256'h020201010001010008090c0c0c0b0d0b0b0b0802070404030100080a0a0c0c0d;
    encBuf[5325] = 256'h0c0b0b09000202010008080104060304030302010202020100090d0e0c0c0a09;
    encBuf[5326] = 256'h090008080908020505040201080a090a08090a0a0c0b0a090100000a0c0c0a08;
    encBuf[5327] = 256'h02070503030201000009090c0c0b0b0900020200080900040705030101090a0b;
    encBuf[5328] = 256'h0b0b0c0b0b0a090104050302000a0b0c0b0a0909080a0b0e0b09000506040303;
    encBuf[5329] = 256'h0108090800000100090a0a080203000e0f0d0b0909010303040203030301000a;
    encBuf[5330] = 256'h0d0b0b0b0b0c0c0b09080002000808000306040201010003050503020108090b;
    encBuf[5331] = 256'h0c0c0c0b0b0b0a0a00020503040108080003060402080a0c0a08010303080b0e;
    encBuf[5332] = 256'h0b0b090a0b0d0b0c0a0803050404020008090908020405020108090002040300;
    encBuf[5333] = 256'h0a0f0d0a090908090a0b0a0104060402010800080808090a0c0c0b0908020203;
    encBuf[5334] = 256'h0208080900020603040100080a0b0a0909090a080004050401080b0e0a090001;
    encBuf[5335] = 256'h01090c0b0a01060502020102020402010a0f0d0b0b0a0a090808010305040202;
    encBuf[5336] = 256'h0008090008080a0a0803070500090d0b0005060302090b0e0a09000001000808;
    encBuf[5337] = 256'h00000000090a0c0901050503020a0f0c0b0a0104050301080a0b0b0900010305;
    encBuf[5338] = 256'h02040201090d0e0b0b0901050402000a0b0c0900020304020108090b0b0d0b09;
    encBuf[5339] = 256'h0004050402010a0d0d0a0a000204040201000a0c0b0b09000304050201080a0b;
    encBuf[5340] = 256'h0c0b09080103040302000a0c0c0b09000306040201090b0c0a0a080000000001;
    encBuf[5341] = 256'h020302000c0c0b0803070201080b0c0901030401000a0b09000301090f0c0b09;
    encBuf[5342] = 256'h00030201000a0900040603030200080a09090a0a0e0c0b0b0901020302000800;
    encBuf[5343] = 256'h01040304010809090b0b0b0b0b0002070403030100080a0a0b0d0a0b09000101;
    encBuf[5344] = 256'h0100080407040402080a0e0c0a0a0908080800010205030301090b0d0a010604;
    encBuf[5345] = 256'h0401000a0a0b0908010108080a0a0808080a0d0e0b0b090307050201000a0b0b;
    encBuf[5346] = 256'h0a0001040202020108090c0c0b0b0801040303020100090d0c0c0b0801040302;
    encBuf[5347] = 256'h000a0b0b0a0001020203040402000a0d0a010606030301090c0c0c0b0b0b0a0a;
    encBuf[5348] = 256'h080204050303030101000808090a0b0e0b0a0a08020403020200000808020404;
    encBuf[5349] = 256'h04000b0f0e0b0a090104030302020008000a0b0e0b0c090104030401080b0b0b;
    encBuf[5350] = 256'h08030603020108090a0c0c0b0d0a0a0901020304020302030302000a0c0b0803;
    encBuf[5351] = 256'h0403090e0d0a090105030200090c0b0b0b0909090909010307040302000a0d0a;
    encBuf[5352] = 256'h0901040301090c0c0a0004030302000908000202000b0f0b0c09080102080c0e;
    encBuf[5353] = 256'h0c0b090802050303020202030203000a0d0c0b0908010101090a0c0b0b0c0a08;
    encBuf[5354] = 256'h00030704030200090c0b0b0a090809080206040401000a0a090002040201090a;
    encBuf[5355] = 256'h0a0b0d0c0b0c0a01040603030200090a0d0b0d0b0b0b08010405030203020200;
    encBuf[5356] = 256'h080a0b0a0a000202090d0d0a0a080000090b0b0a00040403030008090b0c0901;
    encBuf[5357] = 256'h050604030201020102080a0f0d0b0b0900010201080a0b0a0801030506040301;
    encBuf[5358] = 256'h080b0f0c0a0a08000102030504030301080a0b0a080800090b0c0c0b0d0a0a00;
    encBuf[5359] = 256'h01040302080b0d0a0802050403020101010100090a0b0d0b09090008080a0c0b;
    encBuf[5360] = 256'h0a01040403080d0f0b0b0a010503040301010100000a0c0d0a0901040201080a;
    encBuf[5361] = 256'h0b0a000403030100090909080a0a0c0b0c0b0d0b0d0c0a0a0802040404030202;
    encBuf[5362] = 256'h080a0a0c0a000306040304020108080a0b0b0b0b0c0d0c0c0c0b0a0908010406;
    encBuf[5363] = 256'h0403030201090a0a090909090b0c0b0b0a010204020102020503010a0f0e0b0a;
    encBuf[5364] = 256'h090003040304020101000008090808080a0b0c0c0b0b0b0c0a09020605040302;
    encBuf[5365] = 256'h0208090c0b0d0a0a090909090908020505030200080800020202000a0b0b0003;
    encBuf[5366] = 256'h07030401080b0d0d0b0a0b0a0a0c0b0b0902070504020201080008080009090a;
    encBuf[5367] = 256'h0a0a090a0b0e0c0b0a0801020202020305040201080a0a090900080808010304;
    encBuf[5368] = 256'h040303040302000c0f0c0a0900020200090a0b0004060301090c0d0b0a0a0a0b;
    encBuf[5369] = 256'h0c0b0a0802060404030202010100020303030301080a0d0d0e0c0b0c0b090802;
    encBuf[5370] = 256'h0204020100080001020203010800000303020a0e0d0a0900080a0d0d0a090001;
    encBuf[5371] = 256'h0200090a0901070405030100090d0b0b0a000303030200000102030200090005;
    encBuf[5372] = 256'h0502080e0e0c0a080101020008090909090c0d0b090206040100090c09000204;
    encBuf[5373] = 256'h040202010008080a0a0b0b090808090c0e0b0c09080104040303010008000001;
    encBuf[5374] = 256'h080a0f0c0a0a09000008090908020605020201000800010201090d0d0b0c0a0a;
    encBuf[5375] = 256'h080801030503030108080802020202090900030503080f0d0c0a080103030208;
    encBuf[5376] = 256'h0b0d0b0a09090a0c0b090107040200090b0a0004050302000a09090103020109;
    encBuf[5377] = 256'h0b0b09000001080b0c0b0b0c0c0c0b080207060302080a0c0d0a0a0a09080801;
    encBuf[5378] = 256'h030302080c0b080607050201080a0b0a0a0a0a0a0b0802060401010809000103;
    encBuf[5379] = 256'h040101080909090808080a0d0d0d0c0a080104030401000a0b0c0b0b0a0a0801;
    encBuf[5380] = 256'h0102040404040200080a0b0801050303000809010403010a0f0d090003050401;
    encBuf[5381] = 256'h080c0e0b0c090901020304020108090a0b090103060201090a0c090801030202;
    encBuf[5382] = 256'h02040202090e0d0c0a09000008090b0c09010405040303020108090a0b0a0800;
    encBuf[5383] = 256'h01010a0d0d0b0a080306040303080c0e0c0b0909000100000800010305030303;
    encBuf[5384] = 256'h0304040301090b0f0a0a0800000008090808000000000000000a0f0d0c0b0900;
    encBuf[5385] = 256'h020402020008080801030703040200090b0c0a090808090a0b0a0908090a0b0a;
    encBuf[5386] = 256'h0507060202080809090808090a0c0a08010202080800040704020200090a0a0b;
    encBuf[5387] = 256'h0a0b0b0e0c0c0a0b09000000080900020605030202030504030200090a0a0908;
    encBuf[5388] = 256'h090c0e0b0b0a080008000900000001000808000304040108080a0b0b0b010707;
    encBuf[5389] = 256'h06030100090b0a090900090b0d0c0b0b0b0b0a00030705040302020100080909;
    encBuf[5390] = 256'h090a0b0d0d0b0a08020403030108090000030301090e0d0c0b0b0a0b0a090001;
    encBuf[5391] = 256'h0204030101010307060404020200000a0b0d0b0b090800010200090909090801;
    encBuf[5392] = 256'h020301090e0f0b0c0a080103050203020302010000090a090a0b0c0c0b090003;
    encBuf[5393] = 256'h0402000a0c0b0900000100000a0f0d0d0b0a080405040202010102020201080a;
    encBuf[5394] = 256'h0a0b0b0d0d0b0c0a0908000800010100080a0e0b0a080202000b0f0d09000506;
    encBuf[5395] = 256'h04030201000908080000080b0c0b0b09090a0d0b0b0a000302000a0a0a010505;
    encBuf[5396] = 256'h0201080b0d0a0a00040504030301000008010205030302080c0e0e0c0b0b0b08;
    encBuf[5397] = 256'h000101020102020404040203020201000b0f0b0b090801010101000202030401;
    encBuf[5398] = 256'h090c0e0c0b0c0a0a090908010204040303010001040404020108080a0a090a0a;
    encBuf[5399] = 256'h0a08000008090c0b0b000102000c0f0e0c0b0c09090102030201020406050302;
    encBuf[5400] = 256'h010a0b0b0a000202010a0b0b0a00080a0e0d0b0a0a0800080009080103070604;
    encBuf[5401] = 256'h03030208080b0a0a080000090b0d0b09000202090c0e0a09000101090d0c0908;
    encBuf[5402] = 256'h010301080a0b0a02070704040303010009090b0a0c0c0b0d0a09090000010203;
    encBuf[5403] = 256'h04020301080a0a0c0c0d0b0c0a09020404040302030303040100090a0d0b0c0c;
    encBuf[5404] = 256'h0c0b0b0a0908010103030403050303030201000a0c0d0b0a0b09080204050402;
    encBuf[5405] = 256'h000808090800000a0d0d0b0b0a090a0a0a080105040302020102020503030402;
    encBuf[5406] = 256'h01080a0c0c0b0a0b0b0a090004060303010809090a0a0c0e0b0c0a080008090c;
    encBuf[5407] = 256'h0d0b0a00050504030302010000000000010000080a0d0f0c0b0b0a0800010200;
    encBuf[5408] = 256'h08080a0801020403030201000102050405030301010800000101000a0d0d0b0a;
    encBuf[5409] = 256'h0b0d0e0c0c0b0b09000002010102050504040301010809090a0a0a0b090a0808;
    encBuf[5410] = 256'h0802030504040200080b0d0b0c0b0a0a0a0a0a0b0b0c0b0a0804060503050202;
    encBuf[5411] = 256'h020101000001020301080d0e0c0a0b09090809080808080009090a0901020403;
    encBuf[5412] = 256'h02010101050605040304010100080a09080908080a0c0e0c0c0b0b0b09090800;
    encBuf[5413] = 256'h01010203030403050404050302020009090a0b0a0b0b0a090a0808080000000b;
    encBuf[5414] = 256'h0f0e0c0a0a0001040200090b0d0b0908030505030502020101010101080b0c0c;
    encBuf[5415] = 256'h0c0a0b0c0b0b0b09010304040101010102030400080b0e0a0a08000102030404;
    encBuf[5416] = 256'h030302000800010103080b0f0f0c0b0c0a0a0a09090001020404040304030503;
    encBuf[5417] = 256'h0202000a0c0c0b0b0b0a090901020304030200090a0a090b0d0d0d0b0a0a0801;
    encBuf[5418] = 256'h0304040404030203010001010100080a0e0c0c0a0b0b0b0b0a09000205040203;
    encBuf[5419] = 256'h0202030302020a0e0d0c0b0a080002030403030503020101080908080108090e;
    encBuf[5420] = 256'h0e0c0c0c0a0a0900010303040303020101000001020202090c0d0c0b09080203;
    encBuf[5421] = 256'h060303040200000a0d0c0c0c0b0b0a0800000100080001030705040201010809;
    encBuf[5422] = 256'h090908080800000101000b0d0d0b0b0a0104040301080b0d0b0b080001080b0d;
    encBuf[5423] = 256'h0c0b0902040602030101010305040303010108090c0d0d0c0c0a090800000101;
    encBuf[5424] = 256'h00000002020303030208090b0b0d090900010406050404020008090c0a0a0909;
    encBuf[5425] = 256'h090a0b0c0b0a0a0b0c0b0b080405050403020201000009090908090008080a09;
    encBuf[5426] = 256'h090103040201080b0c0b0c0d0c0c0c0b0b0a0a09080001020504030404020403;
    encBuf[5427] = 256'h0303040202010008090a0e0c0d0b0c0a09090909090909000204040303030202;
    encBuf[5428] = 256'h0202020100010103040401000c0d0b0a0006050303000a0e0c0c0b0b0b0b0b0a;
    encBuf[5429] = 256'h080103040603050303030201000809090b0d0b0c0b0a0a080001020404030200;
    encBuf[5430] = 256'h090c0c0b0b0c0a0c0a0a09010305040304020303040203020108080b0d0c0d0b;
    encBuf[5431] = 256'h0c0b0b09090001010101010204040403020108090a0b0b0b0a0b0a0901040603;
    encBuf[5432] = 256'h05040203040201000a0d0c0c0c0b0b0a0a09090a080102060403040201020101;
    encBuf[5433] = 256'h010101080a0c0b0c090908080101040303020a0f0c0d0a0a0a090a0b0a0b0c03;
    encBuf[5434] = 256'h0707000000000800080008000800080008000800080008080008000008000008;
    encBuf[5435] = 256'h0000090008080108080008080008000000020100090d0a080a01030908010a00;
    encBuf[5436] = 256'h010901020004080007010803000b080a0c080b0a090d0a090902000903020407;
    encBuf[5437] = 256'h0100000009010809080b0e0b0b0105020000090103020000080f0a0801000202;
    encBuf[5438] = 256'h0008090b0b0801000b08020201010003090f090808000000080900010901010a;
    encBuf[5439] = 256'h090304020308000403010808080e0c090909080a0a080102010405030803000b;


    decBuf[0] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[1] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[2] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[3] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[4] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[5] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[6] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[7] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[8] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[9] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[10] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[11] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[12] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[13] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[14] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[15] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[16] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[17] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[18] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[19] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[20] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[21] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[22] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[23] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[24] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[25] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[26] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[27] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[28] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[29] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[30] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[31] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[32] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[33] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[34] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[35] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[36] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[37] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[38] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[39] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[40] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[41] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[42] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[43] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[44] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[45] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[46] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[47] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[48] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[49] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[50] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[51] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[52] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[53] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[54] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[55] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[56] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[57] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[58] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[59] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[60] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[61] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[62] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[63] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[64] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[65] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[66] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[67] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[68] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[69] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[70] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[71] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[72] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[73] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[74] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[75] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[76] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[77] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[78] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[79] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[80] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[81] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[82] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[83] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[84] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[85] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[86] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[87] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[88] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[89] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[90] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[91] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[92] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[93] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[94] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[95] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[96] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[97] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[98] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[99] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[100] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[101] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[102] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[103] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[104] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[105] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[106] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[107] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[108] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[109] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[110] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[111] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[112] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[113] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[114] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[115] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[116] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[117] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[118] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[119] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[120] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[121] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[122] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[123] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[124] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[125] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[126] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[127] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[128] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[129] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[130] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[131] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[132] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[133] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[134] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[135] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[136] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[137] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[138] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[139] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[140] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[141] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[142] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[143] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[144] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[145] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[146] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[147] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[148] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[149] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[150] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[151] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[152] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[153] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[154] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[155] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[156] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[157] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[158] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[159] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[160] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[161] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[162] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[163] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[164] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[165] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[166] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[167] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[168] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[169] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[170] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[171] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[172] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[173] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[174] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[175] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[176] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[177] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[178] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[179] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[180] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[181] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[182] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[183] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[184] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[185] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[186] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[187] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[188] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[189] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[190] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[191] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[192] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[193] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[194] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[195] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[196] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[197] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[198] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[199] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[200] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[201] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[202] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[203] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[204] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[205] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[206] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[207] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[208] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[209] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[210] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[211] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[212] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[213] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[214] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[215] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[216] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[217] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[218] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[219] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[220] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[221] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[222] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[223] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[224] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[225] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[226] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[227] = 256'h010000000100feff010000000100000001000000010000000100000001000000;
    decBuf[228] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[229] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[230] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[231] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[232] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[233] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[234] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[235] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[236] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[237] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[238] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[239] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[240] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[241] = 256'h0100000001000000ffff00000100000001000000010000000100000001000000;
    decBuf[242] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[243] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[244] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[245] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[246] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[247] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[248] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[249] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[250] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[251] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[252] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[253] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[254] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[255] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[256] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[257] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[258] = 256'h0100000001000000010000000100020001000000010000000100feff01000000;
    decBuf[259] = 256'h0100000001000000ffff00000100000001000000fffffeff0100000001000000;
    decBuf[260] = 256'h01000000010000000100feff010000000100000001000000010000000100feff;
    decBuf[261] = 256'h0100000001000000010000000100feff01000000fffffeff0100000001000000;
    decBuf[262] = 256'h0100feff01000000010000000100000001000000010000000100000001000000;
    decBuf[263] = 256'h01000000010002000100000001000200ffff0000010000000100000001000000;
    decBuf[264] = 256'h0100000001000000010000000100000001000000fffffeff01000200ffff0000;
    decBuf[265] = 256'h01000000ffff000001000200ffff000001000000ffff00000100000001000000;
    decBuf[266] = 256'h01000000010000000100000001000000ffff0000010000000100000001000000;
    decBuf[267] = 256'h01000000ffff00000100000001000200ffff0000010000000100000001000000;
    decBuf[268] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[269] = 256'h010000000100000001000000fffffeff010002000100feffffff000001000000;
    decBuf[270] = 256'h010000000100feff0100000001000000010000000100feff0100020001000000;
    decBuf[271] = 256'h0100000001000000010000000100000001000000010000000100000001000200;
    decBuf[272] = 256'hfffffeff01000000ffff00000100000001000000010000000100000001000000;
    decBuf[273] = 256'h0100feff0100020001000000010000000100feff0100020001000000ffff0200;
    decBuf[274] = 256'h01000000010000000100000001000200ffff0000010000000100000001000000;
    decBuf[275] = 256'h01000000010000000100000001000000010000000100000001000200ffff0000;
    decBuf[276] = 256'h01000000010000000100000001000000010000000100000001000000ffff0000;
    decBuf[277] = 256'h01000000010000000100feffffff000001000000010000000100000001000000;
    decBuf[278] = 256'h0100000001000000ffff000001000000010000000100000001000200ffff0000;
    decBuf[279] = 256'h01000000010000000100000001000200fffffeff01000000fffffeff01000000;
    decBuf[280] = 256'h01000000010000000100feff01000200ffff0000010000000100000001000000;
    decBuf[281] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[282] = 256'h01000000010000000100feff0100000001000000010000000100000001000000;
    decBuf[283] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[284] = 256'h01000000010000000100000001000000ffff0000010000000100000001000000;
    decBuf[285] = 256'h0100000001000000010000000100000001000000010002000100000001000000;
    decBuf[286] = 256'h010000000100000001000200ffff000001000200fffffeff0100000001000000;
    decBuf[287] = 256'h010000000100000001000000fffffeff01000000010000000100000001000000;
    decBuf[288] = 256'h0100000001000200010000000100000001000000010000000100000001000000;
    decBuf[289] = 256'h01000000010000000100feff010000000100feff010000000100feff01000000;
    decBuf[290] = 256'h0100000001000000010000000100feff0100020001000000ffff000001000000;
    decBuf[291] = 256'h0100000001000200ffff000001000000ffff000001000200ffff0200fffffeff;
    decBuf[292] = 256'h01000000010000000100000001000000ffff0000010000000100000001000000;
    decBuf[293] = 256'h0100feffffff00000100000001000000010000000100000001000000fffffeff;
    decBuf[294] = 256'h01000200ffff00000100000001000000fffffeff01000200ffff00000100feff;
    decBuf[295] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[296] = 256'h010000000100feff010000000100000001000000010000000100000001000200;
    decBuf[297] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[298] = 256'hffff000001000000010002000100000001000000010000000100000001000200;
    decBuf[299] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[300] = 256'h010000000100000001000000fffffeff01000200fffffefffffffeff01000000;
    decBuf[301] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[302] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[303] = 256'h010000000100feffffff000001000000ffff0000010000000100000001000000;
    decBuf[304] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[305] = 256'h0100feff01000200010000000100000001000000010000000100000001000200;
    decBuf[306] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[307] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[308] = 256'h010000000100020001000000ffff000001000000010000000100000001000000;
    decBuf[309] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[310] = 256'h0100000001000000010000000100000001000200ffff00000100000001000000;
    decBuf[311] = 256'h01000000010000000100000001000000010000000100feffffff00000100feff;
    decBuf[312] = 256'hffff00000100000001000000010000000100feff010000000100000001000200;
    decBuf[313] = 256'h010000000100000001000000010000000100000001000200ffff00000100feff;
    decBuf[314] = 256'hffff000001000000010000000100000001000000010000000100000001000000;
    decBuf[315] = 256'h0100000001000000010000000100feff01000000fffffeff01000200fffffeff;
    decBuf[316] = 256'h01000000010000000100000001000000010000000100000001000200fffffeff;
    decBuf[317] = 256'hffff000001000000010000000100feffffff00000100000001000200ffff0000;
    decBuf[318] = 256'h010000000100000001000000010000000100000001000000010000000100feff;
    decBuf[319] = 256'h0100000001000000010000000100000001000000010000000100000001000000;
    decBuf[320] = 256'h01000200ffff0000010000000100000001000000010000000100000001000000;
    decBuf[321] = 256'h0100000001000200ffff0000010000000100000001000200ffff00000100feff;
    decBuf[322] = 256'h01000000010000000100000001000000fffffeff0100feff01000200ffff0000;
    decBuf[323] = 256'h01000000fffffefffffffeffffff00000100000001000200fffffeff01000200;
    decBuf[324] = 256'hfffffeff01000000010000000100000001000200fffffeff0100000001000000;
    decBuf[325] = 256'h01000000010000000100feffffff00000100000001000200010000000100feff;
    decBuf[326] = 256'h01000000ffff000001000000010000000100feff01000200ffff000001000200;
    decBuf[327] = 256'h01000000ffff000001000200ffff00000100feffffff00000100000001000000;
    decBuf[328] = 256'h010000000100000001000000010000000100feff01000200fffffeff01000000;
    decBuf[329] = 256'h0100000001000000010000000100000001000200ffff00000100000001000000;
    decBuf[330] = 256'h01000000010000000100000001000000010000000100feffffff000001000000;
    decBuf[331] = 256'h01000000fffffeff010000000100feffffff0000010000000100000001000000;
    decBuf[332] = 256'h0100000001000200fffffefffffffefffcfffbff01000c0018001300ffffeaff;
    decBuf[333] = 256'hf8ffffffecffdeffeffffeff0400100018000b00f4fff1fffaff01000d000f00;
    decBuf[334] = 256'h0d0008000a000b000f001b0028002d0029001500fdff0d002d002800eeffd6ff;
    decBuf[335] = 256'hddfff2ffdffffbff29002f001f00240032002d0012000800050007000f000800;
    decBuf[336] = 256'hf9fff3fff9fffdfff9ffe7ffcdffc2ffd2ffd5ffbdffcdfff8ff24001e002e00;
    decBuf[337] = 256'h45001600c5ffbaffecff0700deffb8ffa4ffb6ffc7ffe1ffe6ffeaffeeffe3ff;
    decBuf[338] = 256'hdaffe2fffaff160031002700f8ffacffcafff8ff1100450083005a0007002800;
    decBuf[339] = 256'h6e002e00b3ff59ffabfff4ff1c0029001e0000000900110009000300f0ffc8ff;    
    decBuf[340] = 256'h9aff94ff8eff94ffd9ff5b00250015005f00370099ffafff5f00e9ff51ff7800;
    decBuf[341] = 256'hef023d08830ad309730ae1095d09e4085209b5095b09ad09f809b40976093e09;
    decBuf[342] = 256'ha5081a089b0775070c07ed0643075d0716072b073f07e6065306f10598054705;
    decBuf[343] = 256'h5505e905720684067406470604062906600692068906a106c706ce0606077707;
    decBuf[344] = 256'h4a081309ca09410a2b0af009de09ef09e0093d0ac30a400bd20b340c460c360c;
    decBuf[345] = 256'h620c700c330ce60bc80b880b3e0b480b9a0bbb0bb10bba0ba10b4f0b020bbc0a;
    decBuf[346] = 256'h6a0af109c009940951092c0937092d09ee08b4087f08180876073507fa06e806;
    decBuf[347] = 256'hf906250732073e0749076707700779078f078807690763077d079407cb073c08;
    decBuf[348] = 256'hae08f7085509c209ee09fc09200a150a0b0a140a3e0a810ad30a360b790b9d0b;
    decBuf[349] = 256'h920b880b490bfe0ae00ad70acf0ad60add0acb0aa30a750a3d0a080ad809b909;
    decBuf[350] = 256'h9209630938091009e208b6088f0861081008c30769072c0721073f075a077307;
    decBuf[351] = 256'h6c0757072b07ed06d506cd06e206010728075707760787079607a407b907d407;
    decBuf[352] = 256'hed07fc0711081e082e08410854086008620864086208640871088b089f089b08;
    decBuf[353] = 256'h85085a08fd0784071207c906bb06af06a4069a066d062206c8055b05f4049604;
    decBuf[354] = 256'h5a0439042f0426040d040504f103de03cd03b3039c0376034803290318032703;
    decBuf[355] = 256'h51038303a603b903be03a5039703a303c60302043c048004c004d804e004e704;
    decBuf[356] = 256'h060539057605b005d605ea05f105e005d005c205ad058a0557050c05b2045d04;
    decBuf[357] = 256'h2604f403d903af036c0307038f021d0299013f010e01e200ba00960049001700;
    decBuf[358] = 256'hc5ff78ff46ff06ffdcfe99fe6bfe42fe1dfe08fe02fefcfde2fdb9fd86fd56fd;
    decBuf[359] = 256'h37fd3cfd56fd92fddcfd22fe75feacfedefe0bff34ff69ffb5fffbff4d009a00;
    decBuf[360] = 256'he000fb000301fc00e700d400c400be00b1009b00780046001500ddffa9ff86ff;
    decBuf[361] = 256'h67ff4bff27ff07ffe9fecefeaefe88fe50fefdfd9afd3dfdcffca3fc60fc54fc;
    decBuf[362] = 256'h33fc01fcaffb62fb1cfbdcfab3fa8dfa6bfa3ffa0dfaddf9caf9c4f9def907fa;
    decBuf[363] = 256'h3afa6afa89fa9afa9ffa9bfa97fa9afabafae9fa21fb73fbc0fbf2fb20fc39fc;
    decBuf[364] = 256'h31fc0ffcd7fba2fb80fb6dfb7efb98fbaffbaafb97fb63fb2efbfefac6faaffa;
    decBuf[365] = 256'ha8faa2fa91fa82fa61fa33faeef9aef974f94ff948f94ef95ff95af943f903f9;
    decBuf[366] = 256'hb1f84ef8f0f7b4f793f7b1f7def739f88ef8c5f8bbf88df843f8e9f7acf78bf7;
    decBuf[367] = 256'hbdf722f89af80cf973f99bf98ff96ef928f9fbf8f2f809f939f97ef9bef9f7f9;
    decBuf[368] = 256'h2cfa40fa3afa1efae6f9b1f981f955f939f93ef930f924f9f9f8b0f856f819f8;
    decBuf[369] = 256'hccf7aef7b7f7aff7a8f778f733f7cef671f634f6fdf5f3f5fcf515f62cf640f6;
    decBuf[370] = 256'h53f64df61ff6daf5adf573f55df57ff5abf5f4f53af67af692f6a9f6a2f6a8f6;
    decBuf[371] = 256'hb9f6c9f6e9f618f750f793f7e6f71df84ff88ef897f8adf8c2f8e1f814f952f9;
    decBuf[372] = 256'h7bf991f998f985f95ef93af91af90df909f9f8f8e8f8daf8b8f897f879f847f8;
    decBuf[373] = 256'h09f8cff77df730f712f709f701f717f710f7f1f6bef680f647f621f60df6faf5;
    decBuf[374] = 256'hfff5e6f5cff5c2f5a7f5a3f5b3f5bcf5d8f5fbf512f630f65bf682f6b0f6e9f6;
    decBuf[375] = 256'hfff62ff75bf782f7bbf70df844f88af8caf8e3f8eaf8f1f8ebf8daf8dff8dbf8;
    decBuf[376] = 256'hdff8faf819f948f974f990f99ff99bf97df96af966f95df965f978f971f959f9;
    decBuf[377] = 256'h37f9fbf8c1f89cf879f84df831f8f9f7c4f794f775f764f769f765f769f76df7;
    decBuf[378] = 256'h5bf758f772f792f7c9f7fdf72df84df874f898f8c2f8f4f824f944f96bf97af9;
    decBuf[379] = 256'h91f9b8f9e6f912fa4ffa79fa8ffa96fa90fa95faa5fab3fab7fac3fab8faaffa;
    decBuf[380] = 256'hb7fabffae3fa11fb30fb41fb46fb26fb08fbf5fae3fad4facbfaa4fa7cfa4efa;
    decBuf[381] = 256'h16fafff9ebf9d8f9c7f9adf984f95cf943f935f939f94df965f987f9b1f9d8f9;
    decBuf[382] = 256'h07fa3ffa73fab1fadafa00fb30fb68fb9dfbe8fb2efc5cfc75fc7cfc83fc96fc;
    decBuf[383] = 256'hbdfcf6fc39fd79fdb3fdd8fdedfde7fde1fddcfdcefdcafdbefdb4fdaafda7fd;
    decBuf[384] = 256'haafdb1fdb8fdb2fd97fd74fd38fdeefcbcfca1fc88fc8ffc89fc82fc7dfc59fc;
    decBuf[385] = 256'h2ffc08fceefbd7fbd3fbcffbcbfbd5fbd2fbd5fbd7fbddfbeffb0efc34fc6dfc;
    decBuf[386] = 256'hb0fcf0fc3afd80fdc0fdfafd2ffe5ffea3fed1fefafe2fff51ff70ff8dffbbff;
    decBuf[387] = 256'hf3ff270065009f00c500cb00d200b600a6008f007a006600550045003d003500;
    decBuf[388] = 256'h320039003b00390027000400cbff88ff48ff0effdafed3fed9fe00ff2eff5aff;
    decBuf[389] = 256'h76ff71ff5aff34fff1feb1fe88fe63fe5cfe6efea1feedfe47ff9cffe9ff1b00;
    decBuf[390] = 256'h36003e0046004d005f009200d0002b017f01e201250231023c02320229022102;
    decBuf[391] = 256'h29023d025c02790288028d028002740271027a028802a502c002d202db02d802;
    decBuf[392] = 256'hc602b10297027e027502780285029602a0029a028002550223020002ee01f301;
    decBuf[393] = 256'h170253028d02b202d502db02e102d102ba02b602c202d30202034e03a8031504;
    decBuf[394] = 256'h5e04870493045c041604c4038d0383039e03d8030c044a0473047b0474045504;
    decBuf[395] = 256'h2d04ff03e003b903a903a503a903c403e303f9031404330440044c0448043204;
    decBuf[396] = 256'h18040004de03d003dc03e80308042e043d04540461046504760486049a04b704;
    decBuf[397] = 256'hd204eb040d0537056905b505fb053b0675068b06920698069306a206cc06f306;
    decBuf[398] = 256'h1707400751074c073e072107f606cf06a00681067c0681068f06a406af069e06;
    decBuf[399] = 256'h7c063f06f505af058205690552053e052b0531052b051e0522051605fe04e804;
    decBuf[400] = 256'hbd049104750465046104650469045e045b04580456047504a304cf0402051605;
    decBuf[401] = 256'h10050b05f104da04e70409054605a005f50542069c06d906e406ee06c0069706;
    decBuf[402] = 256'h80066c067f06b106e1060d0734073a072c0727071c07110714070c07ef06dc06;
    decBuf[403] = 256'hbc06a706ab06ae06b106b406a2067e0665063b061406fa05da05bc05a1057a05;
    decBuf[404] = 256'h6105530557055b056c05630549052a05fb04c304ac048a0477047d0477046004;
    decBuf[405] = 256'h5c0450043f043604270410040604f203e003e703f103fb030b040d0403040204;
    decBuf[406] = 256'hf903f503ff03fb03ec03da03c003a1039c03a803c703ff033304560468045704;
    decBuf[407] = 256'h34041304ed03de03eb0301041c04490469046e047e04700463045f0455045104;
    decBuf[408] = 256'h5a0462046e04810489048b049a04a004a504b704c304c504cb04bf04a7048004;
    decBuf[409] = 256'h52040d04e003b603a003a703ad03be03cd03bf0388034503ce025c021202ea01;
    decBuf[410] = 256'hc601e70105022002390232020102c90186013401fd00df00c300dc00f200f900;
    decBuf[411] = 256'h0c01fb00d700ae007b004b0045003f0044005b00680074007e008e009c00b900;
    decBuf[412] = 256'hd400f4001a0134014b016001730185019b01af01c101d701eb01fd0112022102;
    decBuf[413] = 256'h290222020e02f701e101cd01c001bd01bb01b901bb01b601a9019c018a017501;
    decBuf[414] = 256'h6101490133011f010801f200d200ac00920072005d0051004e003e002400feff;
    decBuf[415] = 256'hc5ff82ff54ff2bff14ff1bff21ff32ff37ff2aff0cffe1febafea0fe89fe7cfe;
    decBuf[416] = 256'h78fe83fe93fea7feb4febbfeb5fea3fe88fe70fe67fe6ffe82fe9cfeb4febefe;
    decBuf[417] = 256'haffe98fe7bfe68fe5efe61fe69fe7cfe91fe9afe9cfe95fe86fe74fe64fe5dfe;
    decBuf[418] = 256'h5ffe76fe98fecbfefbfe1bff37ff3cff25ff10fffcfef2fe08ff33ff5eff86ff;
    decBuf[419] = 256'h9fffa4ff8fff6cff4cff3fff43ff54ff77ff8effa3ff9fff95ff85ff77ff6fff;
    decBuf[420] = 256'h68ff65ff5bff4cff3dff27ff07ffe9fecefea1fe75fe4efe2afe13fe0efe12fe;
    decBuf[421] = 256'h16fe0cfee1fd9dfd4afdfdfccbfcb0fcb8fcedfc0ffd22fd28fd18fdf8fcd2fc;
    decBuf[422] = 256'haefc97fc8afc95fca7fcd0fc02fd32fd5efd7afd7ffd7bfd6efd62fd6dfd8ffd;
    decBuf[423] = 256'hb9fdebfd29fe53fe78fe9afeadfed5feeefe0fff35ff4eff5cff61ff64ff68ff;
    decBuf[424] = 256'h71ff7aff82ff89ff8bff85ff7cff71ff5aff38ff0effdcfeb9fea7fea1fea6fe;
    decBuf[425] = 256'hc7fed3fedffed4feacfe79fe49fe11fefafde6fdecfd08fe22fe30fe2bfe18fe;
    decBuf[426] = 256'he3fdaffd71fd48fd31fd2afd3dfd65fd88fda0fdacfdb0fd9ffd8ffd81fd74fd;
    decBuf[427] = 256'h7bfd8afda0fdbffdddfdf0fdfbfd04fefcfdf9fdf2fdebfdedfdeffdeefdeffd;
    decBuf[428] = 256'heefde0fdd0fdc1fdabfda3fda0fd9efda4fdaafda1fd96fd88fd72fd68fd6bfd;
    decBuf[429] = 256'h7efda1fddafdfffd21fe34fe2ffe1ffe11fefcfd08fe19fe3cfe65fe8dfea6fe;
    decBuf[430] = 256'hb4feb8fea5fe8cfe7dfe7afe8cfeb0fee8fe1dff4dff6cff72ff6dff56ff49ff;
    decBuf[431] = 256'h35ff2bff28ff2bff28ff2aff24ff12fffdfed7fea9fe7dfe56fe47fe42fe4ffe;
    decBuf[432] = 256'h53fe56fe40fe15feddfd99fd6cfd53fd4cfd52fd65fd60fd46fd26fdfffcd1fc;
    decBuf[433] = 256'hbefcaefca8fcb6fcc3fcdefcfefc24fd48fd68fd7dfd81fd7efd81fd95fdbcfd;
    decBuf[434] = 256'hfafd45fe77feb6fecffed7fedefee4fee9fef9fefdfe0aff16ff20ff36ff56ff;
    decBuf[435] = 256'h74ff8fffa7ffa4ff9bff8eff79ff6bff72ff7eff96ffacffc0ffcdffcfffcdff;
    decBuf[436] = 256'hc3ffb0ff8eff64ff31fff4fecafeb4fe9ffea5feabfea6fea1fe8cfe71fe58fe;
    decBuf[437] = 256'h43fe2efe1cfe15fe17fe25fe3cfe5efe7ffea5febefeccfed1fecdfec2feb3fe;
    decBuf[438] = 256'ha4fe9cfe95fe97fea1feb8fecefee8fe07ff14ff10ff06ffeafecefebdfeb4fe;
    decBuf[439] = 256'hc2fedffe02ff2bff47ff57ff52ff3dff22fffbfed7feb7feaafeaefec7fee9fe;
    decBuf[440] = 256'h13ff24ff33ff38ff22ff07fff6fee0feddfeeafe04ff32ff6aff9effc1ffe0ff;
    decBuf[441] = 256'he6ffe1ffd3ffbdffbaffc4ffd4fff3ff11002c003e004d005600590064006f00;
    decBuf[442] = 256'h81008d0098009e009800900083007a007200730077007b007c0071005b002c00;
    decBuf[443] = 256'he0ff9aff48ff11fff3fed8fee0fef7fe19ff2cff26ff0cffe3feb0fe80fe54fe;
    decBuf[444] = 256'h43fe53fe73fea2fedafe00ff07ff0dfffcfee2fed4fed0fee4fe03ff32ff6aff;
    decBuf[445] = 256'h90ffb2ffd1ffccffd1ffd5ffebff0d004a009400da0007012001280121011b01;
    decBuf[446] = 256'h2b0145016f01a101c401e301dd01b90199016a014b012f0120011b011f011b01;
    decBuf[447] = 256'h11010101e700c1009d0073004c003d0038004d00700090009d008a0063002b00;
    decBuf[448] = 256'hf6ffc6ffc0ffc6ffeaff0a001f00230019000300e3ffd6ffd2ffebff1a005800;
    decBuf[449] = 256'h9100c600f600fc000201f300ee00f2000d0134016c01a101d101e401de01c401;
    decBuf[450] = 256'h9b0173015a0143013e01520163017f018b018e0185016b01530137012b012001;
    decBuf[451] = 256'h240126012401260120011e01200128013801470155015a015f015b0154014901;
    decBuf[452] = 256'h38012901230125013d016b01a301e70114021c0224020202e201d101e1010102;
    decBuf[453] = 256'h30027502a202cc02e202db02c802b8029e0287027a0267025c025f025c026402;
    decBuf[454] = 256'h6b0261024f022b02fd01c5019f017d016a0165015f015b015701430132012201;
    decBuf[455] = 256'h0e010101f500ef00ed00eb00f000fa0009011f013901590176019201aa01ba01;
    decBuf[456] = 256'hc801d501dc01e301ed01f201fa0105021102230242025f027b0293029c029f02;
    decBuf[457] = 256'h97028c0285029302aa02cc02f6021d0337034e034a033e031f03e702b3027502;
    decBuf[458] = 256'h3b021602010214021a021f020802d90188012501e200a50084008e0097009f00;
    decBuf[459] = 256'ha700bc00c200de00f8000f0113010f010501f500f200fa000b0126013a013d01;
    decBuf[460] = 256'h3a012c012e013a0151016e0189018c018901860184019401b401f0012a025e02;
    decBuf[461] = 256'h810287028d02730265025802550258025b02640266025f0248022602f301b501;
    decBuf[462] = 256'h7b0138010a01e100d900d200d900c800ae00840052002f001000fffffaff0800;
    decBuf[463] = 256'h1500200032003b003e0046004d0054006200710084009700ac00bb00cd00d900;
    decBuf[464] = 256'he300e900f6000801260144016f019601b001c701d401d001c501bc01b301b101;
    decBuf[465] = 256'hb801c201c801c301ab018401600137011b010b01fd00f100dd00c500a2008200;
    decBuf[466] = 256'h5c0042002b000d00faffe8ffd9ffc5ffbdffb6ffafffadffa8ffa3ffa2ffa3ff;
    decBuf[467] = 256'hacffbdffd2ffecff0b0021003c00540064007e008f00a500b900d100da00e900;
    decBuf[468] = 256'hfb0002011101230134014701590160016701610154013f012b010e01fb00e900;
    decBuf[469] = 256'hda00cb00c400b800a50088005d003600fdffc9ffa6ff87ff76ff5dff4fff3aff;
    decBuf[470] = 256'h26ff1cff0cff09ff07ff04fffefef8feecfee3fee8fef7fe11ff31ff4eff69ff;
    decBuf[471] = 256'h7bff84ff98ffabffbbffd3ffe9fff7ff040010001b003100500077009a00bb00;
    decBuf[472] = 256'hd000dc00df00e200e500ed00f900ff0005010401fb00f100df00ce00b7009b00;
    decBuf[473] = 256'h780045001500ddffa8ff78ff59ff32ff18fff8fedafeb7fe97fe81fe66fe55fe;
    decBuf[474] = 256'h4bfe43fe45fe51fe64fe86fea7fecdfef1fefffe0cff0fff05ff02fff9fefcfe;
    decBuf[475] = 256'hfefe09ff17ff27ff3aff51ff61ff75ff82ff85ff87ff85ff7fff81ff89ff95ff;
    decBuf[476] = 256'hadffd4fff8ff210032004200460039001e000600e3ffbaff92ff6fff45ff29ff;
    decBuf[477] = 256'h19ff0cff07ff03fff9fef0fedbfecefec7fecefee0fefefe1cff30ff3aff3dff;
    decBuf[478] = 256'h3aff2dff26ff1bff15ff14ff0cff0dff09ff05ff02fffbfeeefed4feb4fe8efe;
    decBuf[479] = 256'h60fe41fe24fe15fe1afe2ffe4afe6afe7ffe92fe9dfea6fea9fea6fea4fe9efe;
    decBuf[480] = 256'h94fe8bfe86fe84fe8bfe9cfeb7fed2fef9fe1dff34ff52ff5dff68ff6bff6eff;
    decBuf[481] = 256'h70ff81ff90ffa6ffbaffd2ffdbffe9ffe7ffe4ffdeffd0ffb6ff9bff74ff50ff;
    decBuf[482] = 256'h27fff4fec4fe98fe65fe35fe0afeedfdcafdb2fda6fd9afd90fd80fd77fd7afd;
    decBuf[483] = 256'h7cfd87fd99fdaafdb4fdb6fdb1fda9fd9efd95fd93fd99fda8fdbffde2fd0bfe;
    decBuf[484] = 256'h3efe6efe9afec1fed1fed5fed1febefeb3feaafeb2fec5fedffefefe1cff28ff;
    decBuf[485] = 256'h32ff2fff21ff09ffe7feb4fe84fe3ffefffdc5fd82fd54fd2bfd06fdf1fcdefc;
    decBuf[486] = 256'hc2fcbdfca6fc99fc7efc6cfc50fc35fc16fc00fcedfbeafbf9fb19fc50fc94fc;
    decBuf[487] = 256'he6fc49fda6fdfbfd48fe8efecefef7fe0eff15ff0efffefeeefee0fee5fe00ff;
    decBuf[488] = 256'h26ff5fff84ffa6ffadff9cff6eff35fff2fea0fe69fe23fee3fdbafd94fd80fd;
    decBuf[489] = 256'h6dfd67fd58fd37fd09fdd0fc8dfc5ffc26fc00fcebfbd9fbbdfb99fb6ffb3cfb;
    decBuf[490] = 256'h0cfbe1fad0fadffaf6fa2dfb71fbb1fbfbfb2dfc5bfc84fca9fcbefcddfc10fd;
    decBuf[491] = 256'h4efd98fd06fe6dfecbfe08ff3fff5dff53ff2aff05ffc7fe8dfe4afe1cfef3fd;
    decBuf[492] = 256'hcdfdabfd98fd87fd78fd6afd4cfd31fd0bfde7fcc6fcbafcbdfccffcf8fc1ffd;
    decBuf[493] = 256'h39fd50fd43fd28fd01fdc9fc94fc64fc45fc29fc1afc1efc33fc4ffc6efc8cfc;
    decBuf[494] = 256'h97fc94fc78fc4dfc26fc0cfc08fc2efc70fcc3fc26fd83fdc0fdf7fd15fe30fe;
    decBuf[495] = 256'h38fe40fe39fe33fe2dfe1efe19fe15fe19fe23fe39fe53fe6cfe81fe96feadfe;
    decBuf[496] = 256'hc9fee4fef6fefffefcfeeafed5fec1febefec5fee1fe04ff24ff31ff35ff31ff;
    decBuf[497] = 256'h2eff37ff59ff95ffdfff39008e00c500e300fe0017013d018801ce0133027502;
    decBuf[498] = 256'h9a02a50287026b0253022d02190212020d02fd01ef01e301e701f1010d022802;
    decBuf[499] = 256'h410244024102390237024a027102c6021b037e03db031804390443041504cb03;
    decBuf[500] = 256'h71030403ba0277023b021a02fc01e001b7018201520127011601fc00e500bf00;
    decBuf[501] = 256'h7200f9ff67ffddfe84fe53fe62fe8afeaefecffed9fed0fea7fe72fe5efe58fe;
    decBuf[502] = 256'h52fe57fe49fe34fe19fe0efe24fe4ffeadfe76ff3f00c2003801a40107023c02;
    decBuf[503] = 256'h6d02b702df0203030e03dc029c0252020c02f10109023e02a5020c034f038c03;
    decBuf[504] = 256'h810363032303e902b502920273026d025e0250025d028002c5023303b8035904;
    decBuf[505] = 256'hc5040005ee04bd043804bb034a03e202850260023f02490265028e02e0022d03;
    decBuf[506] = 256'h8703f5033e044c0458044d042f0426041d044304580477049e04ae04bb04d104;
    decBuf[507] = 256'hdc04d904e804d404b70495044f04cd0350039d02c801380181003a0024005f00;
    decBuf[508] = 256'h0001ee01cb020704da044d05b605d505b9056a0552051205fe04ec04dc040805;
    decBuf[509] = 256'h30058505fe0590061a07bb075208b408ea08d908cb08a3087e083108ff07ad07;
    decBuf[510] = 256'h60070607c90692069c06ef0668071a08c10801093c09e3085108790776063c05;
    decBuf[511] = 256'h150409035a02bc019f01ba0160022203d90350043a04d803cc0226012dff51fd;
    decBuf[512] = 256'haafae5f84af73ff573f4b9f3a1f2a2f117f1f0ef16f07ff09bf1dbf3bff678f9;
    decBuf[513] = 256'ha6fceffd52feadfefffe4aff2601cd036608c70c0b13e018aa1c7d21df25b728;
    decBuf[514] = 256'h4e2bb72c492c1f2b5a29bf2774274028e82a802f6336ce3ca4427649364c0b4d;
    decBuf[515] = 256'h494cd8483543633c4d32e8285d206116ab0f2007940189fcc9f9f3f321ede0e4;
    decBuf[516] = 256'he4dad0ce71c327b637add8a16a9d63992b9847994e9cb9a28ea8e4b0a8b8bdc1;
    decBuf[517] = 256'h47cad3cfe3d64edd79e1c7e69aeb7df2e8f813029e0ad216f11e4729ac32373b;
    decBuf[518] = 256'hc340ca43b444df439941c63c2437523011284d203e19d212fd0c33096004feff;
    decBuf[519] = 256'hdffa4bf33bec25e210d6b1ca5bc0f5b6faab98a4339b8a9736943393f4951e9a;
    decBuf[520] = 256'he89dbba21da719aba7ac10aea2ad06ae60aefbaf9cb280b631bc03c36ec99ad2;
    decBuf[521] = 256'h24dbe8e2f8e963f039f687fb98fd79ff2e01b2013a018302ad037205b107bd09;
    decBuf[522] = 256'h990bcd0c050d060c650a8b07450325fef2f771f05de7d3ded7d471cbe7c2ebb8;
    decBuf[523] = 256'he4b4caaeaeada7aa92abbcaa7eabceaa2eaa79a8eba673a6e0a60ba839ab13af;
    decBuf[524] = 256'hcdb538bc64c55fd0b5da1ae416ef78f62efd48039c06a209630c380d7e0f8f11;
    decBuf[525] = 256'h2f12c1124613ec10c80e100ce108080568012dfd0df8daf159ea45e1bbd8bfce;
    decBuf[526] = 256'h59c5cfbc43b733b09dab1da9d7a627a607a8bda94aaba4ad11ae75aecfaed9ad;
    decBuf[527] = 256'hf8acb4ace9ade2af56b382b855bdb7c1b3c541c7b9c726c835c625c5d3c41ec5;
    decBuf[528] = 256'h72c610cab0cddcd270da80e1c0e984f190f6d0fe9406a90fa41aee2771340f43;
    decBuf[529] = 256'hd250e860b76b8b75e87ac87f4e7e477a0e7982737c70bb6d3b6bf5682364405d;
    decBuf[530] = 256'h2a53154736359024c80c9ef679e229d0c1ba5dac84a4619de596dc981297b298;
    decBuf[531] = 256'h209d789e21a275a585acc6b4c2be85cd48db5eeb80fa4308eb1b0029a639c948;
    decBuf[532] = 256'h8c560e632d6b8f724679ef7c0b7e0d7f4d7c22785874246e4f6801636d5b5d54;
    decBuf[533] = 256'h1c4c5844443b4930f325de197f0e290414f8f5ef93e8dde1c3dba7daa5d98fda;
    decBuf[534] = 256'h65db2fdf40e1a2e57ae811eb5bee7ff070f2eaf42af735f911fbc1fcbafe9600;
    decBuf[535] = 256'hc202380414064907f107be073307b8058703e6006cfe88fbd0f80bf770f5bbf5;
    decBuf[536] = 256'h87f6b2f8e9fbc2ff6b048c07880b280f8211a513d014df15d6164c18a019cb1b;
    decBuf[537] = 256'h6c1ee62025233125fd253a26922561232b20761bd415020fc106fdfee9f55eed;
    decBuf[538] = 256'h9ae58fe024daf9d52fd21ed0fdcc47cbb1c838c8cbc72ec83ec97ecb1ece02d2;
    decBuf[539] = 256'haad64ddc1fe38ae90af11ffaa9026d0a7d11be194a1f5524eb28162d5c2f6d31;
    decBuf[540] = 256'h4d33df335b33e2329a31a82fe42d002b472819253f21a01d64194414720f100b;
    decBuf[541] = 256'hcd04a20054fbe2f701f629f3a4f23bf1cdf031f1d6f0cdf118f25cf215f3ddf2;
    decBuf[542] = 256'h10f33ef369f328f4a8f5d9f77afaa8fda7005f038e06b1086a0be30d23102e12;
    decBuf[543] = 256'h1a15d3174c1a8c1c971eeb1f2021c821c722af232e243a25a32502261f266825;
    decBuf[544] = 256'h33240f226f1f401c6718be135c0f3d0a6a0508010cfd63f842f569f2d3ef88ec;
    decBuf[545] = 256'h8ae90ae6c0e2e6de47dbedd8a4d741d79bd792d808dae4db10deb0e02ae30ee6;
    decBuf[546] = 256'hc7e8aaec4af0a3f27df613f96dfb91fd82ff470187039205e60696083e09d709;
    decBuf[547] = 256'h060adc091c0928080b071805b402d0ff17fde9f9eaf66bf311f1c9ef9eeedaec;
    decBuf[548] = 256'he3eb03eb27e9f2e7f9e51de46ce273e01fdf6fdd56dcf1da0ada8bd965d988d9;
    decBuf[549] = 256'h26dab6daa1db00dc8fdca9dcc1dcacdce6dc1cddcfddd4de0ee089e154e304e5;
    decBuf[550] = 256'h8de6bee8c9ea2ded6def0ef287f4c7f63df891f9c6fa6efba1fbcffba5fb32fb;
    decBuf[551] = 256'hcafa2bfa62f977f85af74ef6cef403f3d7f0a1eda3ea5ce660e2c0de76db9cd7;
    decBuf[552] = 256'h06d5acd23ed214d1b9d00cd1ecd1b8d2edd376d5dbd6d9d82dda58dc64de40e0;
    decBuf[553] = 256'h6be20ce53be814ecb4efeff3ebf782faccfdcb00bc02cc03c3040d05c9049503;
    decBuf[554] = 256'h0c0275fffbfc17fa5ff730f40df28dee33ec5ae8c3e588e18cddecd9a1d6c8d2;
    decBuf[555] = 256'h28cfcfcc86cb5cca01ca53ca34cb88ccb3ce29d005d2b5d33ed5a3d68bd706d9;
    decBuf[556] = 256'h6bdab0db7fddabdf21e1ede121e3e9e2b6e22be204e1abdf20dfa1de15df4ee0;
    decBuf[557] = 256'h1ee24ae480e77eea70ece9ee29f19ff203f5e7f72efc9403a90ca417ee240335;
    decBuf[558] = 256'h2644e9516b5eca69386e906fc870746d6968d363a85f5a5ae956c753a84ed549;
    decBuf[559] = 256'hb241b637a12bc2191c09a7f557e3b0d28ec3bab9cab02aafa4b0fcb116b86abb;
    decBuf[560] = 256'h7ac2e5c8bace08d49ddbb1e43bed6ff9cf04250fe81dab2b9b343a43fc50ec59;
    decBuf[561] = 256'h4b65a16f5776717c8d7d8f7ea47d7a792c74f86d7866685f2757634f5448e841;
    decBuf[562] = 256'h133c4135d52e00292e22ed192912190bae04d8fe8af919f638f4a6f334f59df6;
    decBuf[563] = 256'hc0f840fc9afe980151041506b0079108d508a007f7062c0501038b01affffffd;
    decBuf[564] = 256'h56fdbdfc32fc5cfc83fc60fc7ffc9cfc4efca8fb10fb60fae9f9fef9affa13fc;
    decBuf[565] = 256'h10ffc5036709b50ee8141319611e34231525ca265728d0286228382728263225;
    decBuf[566] = 256'h51248523cc22b321b420b61e521cca189d13cb0ee807a7ff1bfa07f1edea61e5;
    decBuf[567] = 256'h56e096dd6bd9a9d8f8d799d82ad9c1db1bde19e160e539e8e1ec43f13ff5dff8;
    decBuf[568] = 256'h0bfedd023f075f0c92126818321c042166256229f92b622df52c912c182a3327;
    decBuf[569] = 256'hb423781f7c1bdd1792146f12b60ff20d560ce10a8d095808cf066a05c9034002;
    decBuf[570] = 256'ha7011c019a01a70226045706f808710b560e0e1188132315031647168e15e614;
    decBuf[571] = 256'he7134512bc10f10e410db80b530ab20899070007d206a8061b07c9072808f108;
    decBuf[572] = 256'h74091a0add0afc0b560df70ef010cc12f81403176719a71b481e0c200321e321;
    decBuf[573] = 256'h9f216a20011e1d1bd616da12310e100b140774032a002bfdacf961f663f3aaf0;
    decBuf[574] = 256'h7ced7deafee6a4e45be331e2d6e1cde243e4a7e68be90bed64ef63f21bf5e0f6;
    decBuf[575] = 256'h20f92bfb8ffd2aff35018902be0367040005d10453049303e502c8016f002aff;
    decBuf[576] = 256'h5bfdaafb41f901f760f432f10eef56ecdce941e836e65ae425e30de274e145e1;
    decBuf[577] = 256'h6fe1e2e191e2f0e27fe39ae3e1e322e484e401e5b4e52ae6c2e6fde60fe7fee6;
    decBuf[578] = 256'hd2e674e638e617e695e518e544e408e38de18ee049dfcbdef1de5adf77e0d0e1;
    decBuf[579] = 256'h15e33ce495e57de6f8e7c3e973eb6cedd0ef6cf177f3cbf400f618f7b1f73cf8;
    decBuf[580] = 256'hbbf82ef9c5f866f89df77ef624f583f3faf1c9efbeede2eb3be9c1e681e476e2;
    decBuf[581] = 256'h9ae0eaded1dd38dd50dcd2dbf8db1bdc7adcb6dd31dffce028e3c9e542e827eb;
    decBuf[582] = 256'h18ed92ef2df1a3f2f7f32bf5b4f619f817fa6bfb1cfd34fecdfe58ffdafe1afe;
    decBuf[583] = 256'he0fc11fbe5f844f6cbf342f0e8edeaeaf8e8e9e7f2e612e646e58de474e375e2;
    decBuf[584] = 256'heae16be1f8e0d5e034e151e19fe116e282e233e368e48fe535e7bee8bde948ea;
    decBuf[585] = 256'h1eea5ee9dee713e663e4f9e1badfaeddd2db22da0ad90bd87fd7fed7bed8f8d9;
    decBuf[586] = 256'h73db3edd72defbdf60e148e2c3e3f4e595e8e3edb5f4f5fc29098814c624e933;
    decBuf[587] = 256'hac41c151915c7662d3677369f967f263d85d4c583c51a74c7c48b244df3f3d3a;
    decBuf[588] = 256'he731eb272719640bbcf76be5c5d4a3c5cfbbdfb2ffad85acddadf7b383b993c0;
    decBuf[589] = 256'hd3c85fce6fd5dadbb0e182e8c3f087f8a003f60d0a1a6925bf2fd43b33478951;
    decBuf[590] = 256'hee5a08619466a06b8a6c0a6a40660d60375ae1511d4a0941ef3a6335532ebe29;
    decBuf[591] = 256'h9325c921571ef519d5140310600a9606c401a3fecafb3cfac4f90cfbfefc77ff;
    decBuf[592] = 256'hb7015804d1066d08b708fb08c7075d051e0352ffa9fa48f64bf2a3ed82ea85e6;
    decBuf[593] = 256'hf8e48fe321e34ce410e6abe7b7e993eb43edccee31f0d2f1cbf32ff6b8f9f3fd;
    decBuf[594] = 256'h13034709c710d7176c1c42229027022ba22b342ca62a5c278223da1e781a7c16;
    decBuf[595] = 256'hdc12920fb80b1908ce04f50055fd29f856f3b4ed66e833e25ddc0fd73cd21bcf;
    decBuf[596] = 256'h42ccbecb36cc5ace12d1f6d495d8c1dd94e236e800ecd3f0f4f3f0f787fad2fd;
    decBuf[597] = 256'hf5ffae022705b008fa0baf101115541b7f1fcd243f281f2ab12a2429ca26f022;
    decBuf[598] = 256'h511f151b19177a132011fc0ed20dc20ccc0b810bb50a05097c07e504b601ddfd;
    decBuf[599] = 256'h3dfae3f7c0f55cf5b7f5f7f72dfb2bfeab01050428061a087408c6087c08b007;
    decBuf[600] = 256'h7b06f204270377015e002b00130137036d06460ae60d31112f14e816ac18ec1a;
    decBuf[601] = 256'h621cb61dea1e73207221fd21d022dd23d124ed25fa267a281329e4286927d224;
    decBuf[602] = 256'hef203d1bef15bc0fe6099804c5ff64fb67f7c8f36ef14bef59ed4aec53eb73ea;
    decBuf[603] = 256'ha7e972e8e9e684e53fe415e4d5e4e0e616eaf0ed98f2faf6f6fa96fed102aa05;
    decBuf[604] = 256'h41089a0abe0ce80df80e010e210dcd0b980a0f0910088507b3063f0606053603;
    decBuf[605] = 256'h8f0015fe8dfa42f744f48bf15dee39ec81e9bce77ce59ce4d0e389e432e5fde6;
    decBuf[606] = 256'h31e8bae953ea82ea03eaf7e803e8e6e673e6c4e526e5d0e44de4a7e366e353e3;
    decBuf[607] = 256'h88e33be4e1e4a4e5f2e57ce562e409e368e14fe01ce004e1d3e2ffe435e834eb;
    decBuf[608] = 256'h25ed9fef3af145f399f4cef576f60ff7e1f663f6a3f53af5dbf4bff40df584f5;
    decBuf[609] = 256'hc5f58af5e9f4a4f3a6f1caef9fed93eb2fe994e71ee642e40ee385e186e0fbdf;
    decBuf[610] = 256'h25e0e5e064e22fe45be666e8caea0aed80ee5cf00cf225f38af4cef5f5f602f8;
    decBuf[611] = 256'hf6f8d3f9d6fa10fce2fca2fd51fe31fedbfdf0fc55fbccf901f8d5f55ff493f3;
    decBuf[612] = 256'hdaf232f2fff173f1f5f082f08eef2fefd9ee56ee3eee29eeeeed71edffec7aec;
    decBuf[613] = 256'hd9eb6deb0bebd5ea06eb6debe6eb78ec50ede0ed2eee46eeaeedafec30eb65e9;
    decBuf[614] = 256'hbde6f9e4b9e218e054de5ddd7ddcb1db73dbcbdafeda2cdb02db75dbafdcd6dd;
    decBuf[615] = 256'hc9dfb5e234e67fe958edf8f033f577fb4c01260b3b179a22d832fa41ac53905f;
    decBuf[616] = 256'h606a3474fd755d74e3722d6ca363175e07579c50c64afc462942473bdb34062a;
    decBuf[617] = 256'hbc1ca60c84fdd2eb2cdb0acc47be57b5b8b332b5e8bb02c2c6c9dad264db28e3;
    decBuf[618] = 256'h38eaa3f079f64bfd8c05500d6416ef1eeb28ff341f3d694a5853785bce65846c;
    decBuf[619] = 256'h2d7049714b728b6fb5696764d35cbf53344b7043603ccb37f5312b2e1a2c392a;
    decBuf[620] = 256'h8428ed259423ba1f1b1cdf17e3134310da0e920dbc0ecc0f67117213c6148015;
    decBuf[621] = 256'hb8151f15da135f122e10620cc3089703c4fe22f950f2baed8fe9c5e515e574e4;
    decBuf[622] = 256'h2ae6c0e80becbff021f541fa13ff75037107110b5c0e5a111314f6179f1c4122;
    decBuf[623] = 256'h8f27c22d98336237d43a743be23a43370733e82d152932229c1dc7177912a60d;
    decBuf[624] = 256'h04083a0467ff46fc4af8aaf460f186ede7e99ce6c3e22ce0e1dc99db6eda14da;
    decBuf[625] = 256'h0bdb80dce4de6de2a9e6c8ebfcf127f675fb47002802dd036b05f2048504e804;
    decBuf[626] = 256'h43053a06af078b093c0ba50de50f5a11261264124c11810fd90cab09ac06bb04;
    decBuf[627] = 256'h4102ef01a4017002a5032e059306d807a709570be00cab0ed7104d121913d213;
    decBuf[628] = 256'h0a143d14c8144615a016e41760195f1a8d1aba19611863167713f70fad0cd308;
    decBuf[629] = 256'h2b04c9ffa9fad7f5b5f200f17cf0e5f12df31ff5e3f67ef88afadefb09fe1500;
    decBuf[630] = 256'h01038006cb09c90c4910a312a1159317c11ae51c6420be22e2240c26fd246123;
    decBuf[631] = 256'h2b20521cb21877149e11fe0da50b8109900716057b030502b100f8ff4fffeafd;
    decBuf[632] = 256'hecfb88f9a4f6ecf327f230f111f265f390f59cf778f931faf9f960f91bf8a0f6;
    decBuf[633] = 256'h3bf5f6f3cff229f130efccec8ceaece727e68ce4ace3f0e32de466e499e46ae4;
    decBuf[634] = 256'h94e407e5fce557e756e9baeb55ed60efb4f0e9f101f366f465f6c9f8adfb9efd;
    decBuf[635] = 256'h18006a001f0043fe9cfb6ef894f4f5f0aaedabeaf3e7c4e4c6e146defcdafdd7;
    decBuf[636] = 256'h45d580d38ad2a9d1ddd024d00bcf72ce44ce17cf0ad1f6d375d7b0dbaddf43e2;
    decBuf[637] = 256'h8ee58ce87eeaf7ec37ef42f196f2cbf393f3faf259f1d0ef6bee83edb0ec8aec;
    decBuf[638] = 256'h67ecc9ebc6ea46e97be750e544e368e1afe007e06edf3fdf15dfefdeccde2bdf;
    decBuf[639] = 256'hf4df14e1bae2b3e48fe63fe858e9f1e91fea49ea70ea92eab2eacfeab5ea3eea;
    decBuf[640] = 256'h7be9c4e8bfe711e7b2e622e608e6c1e5fee413e436e3c0e1c1e036e060e020e1;
    decBuf[641] = 256'h9fe26ae41be6a4e709e94deac8eb2ded72eeedef52f1ddf107f247f1c8effded;
    decBuf[642] = 256'h4dec53eaffe846e82ee795e6ade586e493e22fe04bddcbd990d5b7d20fceedca;
    decBuf[643] = 256'h15c87ec524c3dcc178c11ec170c150c2a4c3d9c462c6c7c7c5c929ccb2cfedd3;
    decBuf[644] = 256'h0dd940df16e56cedf8f20cfc9704930ea71a462909371e47415615600569e46d;
    decBuf[645] = 256'h5e6f576bae67ea5fd6564b4e8746783f0c398c317c2a3c2240182b0c8cfdc9ef;
    decBuf[646] = 256'hb4df91d0cfc24cb62daebfa967a810acd4b3e8bc73c56fcfd4d85fe123e937f2;
    decBuf[647] = 256'h51f84d02b30b3d14011c1525a02d6435743cdf425f4a6f510556305afa5daa5e;
    decBuf[648] = 256'hc95cf1593f546d4d0247823f6d365330c72abc25fc22272265211522f6236423;
    decBuf[649] = 256'hd6217d1fa31b0418c813cc0f3e0ed50c430da60d4c0dfa0c840b20093c06bc02;
    decBuf[650] = 256'h81fe84fadcf57af15aec88e7e6e198dc26d9c4d4ebd167d1dfd103d482d7aedc;
    decBuf[651] = 256'he2e262ea72f1b2f976018608f10e1c13e616581a791d762115255129702ee231;
    decBuf[652] = 256'h033595351135c631122d6f279d20321ab212a20b370561ff13faa1f63ff243ee;
    decBuf[653] = 256'ha4ea4ae826e635e470e2d5e05fdf0bde52ddaadcdddcc5ddebde92e08be2efe4;
    decBuf[654] = 256'hd3e752eb9dee52f3b3f7b0fb4fffa901f1025503fa025f017f00b3ff75ff8e00;
    decBuf[655] = 256'hf3014e043207ea09640ca40eaf10031238137013a313d113a713cd137c14d815;
    decBuf[656] = 256'h3318171b961ed222aa253827c0267725bf22db1e331a111715137f10340d100b;
    decBuf[657] = 256'h1f095a0764068305b7047a04d103d2023101a8ff77fd01fcadfaebfa74fc0bff;
    decBuf[658] = 256'hee028e06c90ac60e6512b0158919201c6a1f4423da2543278c28ef28e027e926;
    decBuf[659] = 256'h09263d2584244c24b323cb2250211f1f7e1c4f195116d112870f880c0909be05;
    decBuf[660] = 256'hc00207008efd97fce2fc36fee6ff4f02ea0360052c06ee05b6051d0535040b04;
    decBuf[661] = 256'he503c203e203c50377035f0349038403010473046404b6035202bbff8dfc8ef9;
    decBuf[662] = 256'hd6f611f51af4d0f314f451f46af569f651f7ccf831fa19fb94fc93fdc1fd97fd;
    decBuf[663] = 256'hd7fc58fb59fa14f941f81bf8f8f718f835f8b2f77df6aef4fef294f054eedfec;
    decBuf[664] = 256'h8beb56eacde868e7c7e5cee37ae2c0e188e121e266e3e1e446e62ee755e815e9;
    decBuf[665] = 256'hc3e9e0eaeceb6cedd1eeb9efe0f0ecf1e0f23cf4def5d7f73bfa7afcf0fd44ff;
    decBuf[666] = 256'h06ffeefd23fc7cf902f7c2f44df381f243f20bf2d8f1a9f1d7f064f0fbef9cef;
    decBuf[667] = 256'hb9ef07f04ef039f0feef5deff1eeb6eeeceedfef19f1e9f299f4b2f5b1f63cf7;
    decBuf[668] = 256'hbaf72df8dcf8b9f9bcfab0fb0ffcf2fba4fbfdfa91fa2ffa88fa3bfb40fc35fd;
    decBuf[669] = 256'h12fe68fe4efea8fd8ffccffbdbfafdf96ef9ebf845f8d9f74ff71af76bf7d2f7;
    decBuf[670] = 256'h80f856f9acf9c6f9aef9c0f8e3f7e0f632f6d3f5b6f5d0f5e8f5d3f549f585f4;
    decBuf[671] = 256'h65f30cf2c7f0a0efe0ee78ee19eefced7aed74ec3aeb14eabae8d2e754e747e6;
    decBuf[672] = 256'hdfe541e504e4dde21ee2e4e065e03fe0d6dff6df4ce032e04ae0b6e067e16ce2;
    decBuf[673] = 256'h31e4d8e652e9dbec16f112f5bbf99e00de08da12ef1e8e2d513bd34772564660;
    decBuf[674] = 256'h3669d66a506c4968a064145f04589951c34b75464240c138b1317129751f6013;
    decBuf[675] = 256'hc104fef6e9e619dc57ce67c588c00ebf65c07fc60bcc1fd5aadd6ee57eecbef4;
    decBuf[676] = 256'h4afa5a019b09270f3b18551e1926292d9433bf37913e2743fc484a4ebc511e56;
    decBuf[677] = 256'hd3575858ef56cb548550654b9246af3f44391935cb2f592c3829a6282b29a329;
    decBuf[678] = 256'h112a742a652925278424a1200a1ec01ac117d0150b1470126510010e780a2d07;
    decBuf[679] = 256'h790217fe1bfa72f511f114ed6ce80ae40ee06edc24d900d79dd6f7d6dbd95bdd;
    decBuf[680] = 256'h87e2bae83bf04bf78bff87093d10c818541e5f232026a028e62af72cd82eb031;
    decBuf[681] = 256'h3e33a73439340f339530c42b9025101e00179510150909049efdc8f7fef38df0;
    decBuf[682] = 256'h6bed93ea0eeaa5e812e976e9d0e923ea6deab1ea6beb13ec12ed57eed2efd1f0;
    decBuf[683] = 256'h5cf1daf101f224f2c2f28bf3aaf450f6d9f73ef926fa50fa2afa36f9d7f881f8;
    decBuf[684] = 256'h9bf8d0f99ffbcbfd6b009a03bd053d09880c860f0613501674189e19f919a619;
    decBuf[685] = 256'h5c19181955198e198d1ad11ba41cca1c1c1c411add1755140a11310d91095605;
    decBuf[686] = 256'h5901bafd7ff9a6f606f3acf089ee5eed04ed56eda1ed6deea2efbaf01ff21df4;
    decBuf[687] = 256'h81f60afa55fd2e01d705f808f40c9d11be14ba18511b9b1ebf20e92144224d21;
    decBuf[688] = 256'hac1e331caa186f147310dc0d910a9307da041603d600cbfeeffc3ffbb6f951f8;
    decBuf[689] = 256'h0cf791f52cf4e7f215f255f178f116f252f3cdf498f6cdf775f8a8f87af850f8;
    decBuf[690] = 256'hddf774f7d6f60df622f505f45ff2d6f00bef5bedd2ebd3ea48eac9e9f0e913ea;
    decBuf[691] = 256'hf3e910eac1e9aae9bfe9d3e950ea44eb7eeca5edfeee43f069f1c3f2abf37df4;
    decBuf[692] = 256'hf0f413f575f439f315f175eefbeb17e95ee69ae45ae24fe073de47dca6d9e2d7;
    decBuf[693] = 256'ha2d597d343d28ad1e1d048d0bdcf3fcf65cf42cfa1cfa4d0ded1add3d9d5e4d7;
    decBuf[694] = 256'hc0d970dbf9dcf8dd9adfb2e0b1e1f6e274e3e7e3c4e366e30fe3f5e20de379e3;
    decBuf[695] = 256'h78e427e5c5e58ee6dce6f4e635e721e733e764e755e748e723e77ee679e585e4;
    decBuf[696] = 256'h29e3e5e112e105e011dfb2de23dea0dd59dd18dd04dd5eddcfdd8fdeaedfbbe0;
    decBuf[697] = 256'hafe18de21ce3d3e3d8e4cde568e761e93deb69ed74efc8f078f291f32af458f4;
    decBuf[698] = 256'h2ef421f32df2d1f08def12ee13ed2becaceb86eb1debfeeae1ea93ea4beadfe9;
    decBuf[699] = 256'h07e93ee887e7b1e622e6d3e5ebe582e682e7bbe88beab7ecc2ee9ef04ef267f3;
    decBuf[700] = 256'h9af3c8f3f5f2e9f1aff034efcfed2deca5ea40e9fbe7d4e67be536e40fe369e1;
    decBuf[701] = 256'h70df0cddccda2bd8b2d572d3fcd130d16ed117d27cd3d6d516d8b7da30dd15e0;
    decBuf[702] = 256'h06e235e533e825ea53ed52f098f494f84fffba059010e61afb269a355c434c4c;
    decBuf[703] = 256'h6b54d958e05ca85b1c561051a54ad044fe3d9237bd316f2c3b26662094195311;
    decBuf[704] = 256'h570742fbe3ef99e217d6f7cd95c68ec256c1aac4b1c7f2cfb6d7c5de31e5b1ec;
    decBuf[705] = 256'hbcf127f8fdfd4b037e09540fa2147519171f65243829992db9328c37ed3b0d41;
    decBuf[706] = 256'he0450149b64a444ccb4b834a0347c842cc3e1a395035de31bd2e082d832cfc2c;
    decBuf[707] = 256'h442ea82e022f0c2e2b2dc72a3f27f4233f1fde1ae1163912d70ddb093205d100;
    decBuf[708] = 256'hd4fc2cf8caf3f1f05bee01ecdee925e7ace410e305e1b1dff8de30df2fe0e7e2;
    decBuf[709] = 256'hf4e7c7eceaf4aefcc2054d0e4918ff1e19256d28742b5e2c342df62d452da52c;
    decBuf[710] = 256'h132c8f2b162bce29dc2763257f22ff1ec41ac8162813dd0fdf0c260aad071206;
    decBuf[711] = 256'h9c04d0039203ca0363044b0572067f07730811092e09430826073305cf028f00;
    decBuf[712] = 256'h59fd5bfadbf681f483f191ef82ee8bedd6eda2eedfee88efbbef8cef62efd5ef;
    decBuf[713] = 256'h84f01ff2f9f478f8a4fd3805480c5e16c41f4e2812302237b83be33fa540f43f;
    decBuf[714] = 256'h143e3b3ba4385a355b32a32f292de92a74299827f0240d21641c0318e312100e;
    decBuf[715] = 256'hef0a1608890610067e06a807b808530ac90ba50d5e0e770faa0f7b0fa90ee90d;
    decBuf[716] = 256'h690c040bc0094508e0069b05740401046a044705f606190a170d9710e213e016;
    decBuf[717] = 256'h99195d1baf1bfa1b3e1c001ca91c421d861e56200622ff23db251027b827eb27;
    decBuf[718] = 256'h03278825bd239121f11ec21bc4184415fa11200e8a0b3f086504cf0184fe61fc;
    decBuf[719] = 256'h6ffaabf810f79af5cef490f4e8f3b5f3cdf2a6f1e6f038f097f099f1a4f345f6;
    decBuf[720] = 256'hbff8a3fb94fd59ff50009a00ceff15fffdfdfefc16fc43fb1dfb40fbdefb6dfc;
    decBuf[721] = 256'hf0fc67fd51fd3efd08fdd7fc70fc48fcf3fb90fb4dfbf8fa95fa38fab2f9a6f8;
    decBuf[722] = 256'h00f707f5a3f263f0c2ed49ebaee90de748e509e368e0eedd0adb19d909d8b7d7;
    decBuf[723] = 256'h02d8ced87eda77dcdbde1be1bbe380e5c0e7cbe91feb4bedc0ee24f164f305f6;
    decBuf[724] = 256'h7ef863fb54fd19ffb400ff00bb00010079fe14fd72fbe9f984f840f719f6bff4;
    decBuf[725] = 256'h1ef395f130f0ecee70ed0bec24eba8e9a9e865e792e6d2e56ae54ae567e51ee6;
    decBuf[726] = 256'hf3e6f6e730e9abeaaaebefec16ee22ef5cf083f143f2acf2cbf2aef2f8f122f1;
    decBuf[727] = 256'h59f0d6ef5fef75efb0efc2eff2ef3cf064f0d1f091f17cf2d8f379f592f6f7f7;
    decBuf[728] = 256'hdff809f97cf99ff9bff915faccfaa2fba4fc53fdb2fd22fdcefbd0f9e4f62cf4;
    decBuf[729] = 256'hfdf0ffed46eb82e9e6e7dbe5ffe34fe2c6e061df1cdef5dc36dc41dba6d91dd8;
    decBuf[730] = 256'h52d627d4b1d2e5d12cd164d163d204d46ed652d90adceedf8de3b9e88cedeef1;
    decBuf[731] = 256'h31f807fe55038809081118182e22432ea239ec466f53ce5e3066376a6f6b1b68;
    decBuf[732] = 256'h0b61cb58cf4eba429b3a45308e290421781b6814270c63044bf9f5ee8fe594da;
    decBuf[733] = 256'h3ed088c96ec31ac01cc1b2c587cb61d5c7dec2e924f18afa1403a008ab0d4112;
    decBuf[734] = 256'h6c16ba1b8d20ae23aa274a2ba42dec2ea53169330435a5376a39a93b1f3deb3d;
    decBuf[735] = 256'h293e803d813ce03a5739f237ae36db35b535a936c537b839943bc93ce23daf3d;
    decBuf[736] = 256'h0d3c3439b4358830552a7f24ad1d4217c10fb208710075f6bfef34e770df65da;
    decBuf[737] = 256'hcfd5a4d1e2d0d1ce71cf03d088d0e1d205d584d8c0dce0e113e893efa3f6e4fe;
    decBuf[738] = 256'he0084512d01a94229f27352cb52e772fc72ee62c0d2a6e263222591fb11a9017;
    decBuf[739] = 256'h70129d0d3c091c04aa0048fc6ff9e2f779f60bf66ff6c9f6c0f7a0f87cfab1fb;
    decBuf[740] = 256'haafd86ff3601300384043d0505056c04ca0261007dfd36f93af588ef3aea68e5;
    decBuf[741] = 256'h06e1e6db74d894d6ded45ad4c3d50cd7c4d9f3dcf1df71e3ace7ccec9ef141f7;
    decBuf[742] = 256'h8ffcc2029808e60d191444180e1c1f1e0020b5213021b8204b20e71fd81ee11d;
    decBuf[743] = 256'h6b1c8f1adf187516ed12a20fc90b2007be02c2fe23fbd8f7b4f5c3f368f3bbf3;
    decBuf[744] = 256'h30f584f6b9f742f9a7faecfb67fd66feaaffd10077020004cb05f7076d09490b;
    decBuf[745] = 256'h7e0c960d2f0e5e0e880eae0e8b0e2c0ed60d1f0dea0b6f0a0a09c6074b064c05;
    decBuf[746] = 256'h1d05f3041905c805a506a8075608f40884099e0987091a091b08e1061205e602;
    decBuf[747] = 256'hdb00fffe4ffd36fcd1fae9f9c2f81cf704f69ff4fdf2e5f1e6f0feef7fefc0ee;
    decBuf[748] = 256'h57ee77ee93ee4aef7ff0a6f14cf3d5f43af67ef7faf8f9f9e0fab3fb26fc49fc;
    decBuf[749] = 256'ha8fc8bfc71fc59fc18fcdefb84fbf2fa41fa6cf969f875f758f64bf5ccf367f2;
    decBuf[750] = 256'hc5f03def72edc1eb38ead3e8d5e6f9e4c5e3cbe177e0bedfa6de0dde81dd03dd;
    decBuf[751] = 256'h90dc27dcc8db39db1fdb07dbf1da05db17db06db33db40db64dbc7dbf0db14dc;
    decBuf[752] = 256'h35dc03dce8db00dc44dccddcf3ddc2df73e1dce377e583e7e7e982ebf8ecd4ee;
    decBuf[753] = 256'h08f021f1baf1e8f167f28df2b0f2d0f2b3f2fcf1f7f077efe0ec67ea27e8f1e4;
    decBuf[754] = 256'hcde215e050de10dc9bda47d912d8dad7a7d78fd80adad5db00de37e135e4b5e7;
    decBuf[755] = 256'hffea23eddbef55f2f0f3d0f414f5d7f42ef495f3adf2dbf1cef094ef6dee14ed;
    decBuf[756] = 256'hcfebfdeaf0e9fce81fe88fe70ce7c5e65ce70de842e9bdea88ec38ee31f00df2;
    decBuf[757] = 256'hbdf346f545f62df7acf7d2f769f7cbf6c8f58ff468f3c2f1a9f0aaefc2ee44ee;
    decBuf[758] = 256'hd1edaeed10ed46ec5bebffe9bbe894e787e61fe6c0e5a3e589e571e505e5a3e4;
    decBuf[759] = 256'h49e4f8e3aee3bce397e31ee36ce296e15ae033df26de78dd58ddaedd65de6bdf;
    decBuf[760] = 256'ha4e020e285e326e51fe773e81aeb49ee22f2d4f72a00260a3a16d9249c32b242;
    decBuf[761] = 256'hd451975ff364d3694d6b46672c6168595450c9470540f6388a32b52ce325a21d;
    decBuf[762] = 256'ha613910732fcf4eb25e162d372ca93c525c17cc226c6b2cbc6d450dd4ce7b2f0;
    decBuf[763] = 256'h3cf900010c06770ca210f015c21a241f2023c0261a29622a8d2b9c2c932d092f;
    decBuf[764] = 256'h6d31ad33e336e1399a3ca93da03ec03df43c3b3c923bc53bad3c7c3ea8404943;
    decBuf[765] = 256'h0d45a946f346af46ff440643923f473c9337f131a32c6f269a204c1b1815980d;
    decBuf[766] = 256'h880647fe83f674ef33e7a7e1a0deb5dde0dca2ddb3dfd4e2ade53be795e993ec;
    decBuf[767] = 256'h4cefe4f386f9d4fe0805dd0aaf1145161b1ce51f57233725ed266826ff24b623;
    decBuf[768] = 256'hfe20cf1dd11a511707140811890d2f0b0b091a070a065d06d207360a640e6012;
    decBuf[769] = 256'h11185f1dd120f323a8252c26c324a022ae20801da6190716bc12080ea6098604;
    decBuf[770] = 256'hb3ff11fac3f490eebae86ce39ade38da83d8f5d66dd791d910dd4ce16ce63eeb;
    decBuf[771] = 256'he0f02ef662fce203f60c81157d1f3326be2e4a345539403a153b533ae136c033;
    decBuf[772] = 256'hc42f1b2bba269a21c71c65184613730ed108830311006ffaa5f633f352f1c0f0;
    decBuf[773] = 256'h4ef289f6ccfc4d04610dec15b01dbf245529d52b972c482de82d332cae2b5429;
    decBuf[774] = 256'h5626d6229b1e7b19a91447106e0dcf097507510527041703c502100364041406;
    decBuf[775] = 256'h5e09990d95113e16a01a9c1e3b2295249427be28ce29202ad529f927d724fd20;
    decBuf[776] = 256'h551cb2166411920c70099806f8029e007bfec2fb49f9aef7a2f5d6f414f5bcf5;
    decBuf[777] = 256'h87f7b3f954fccdfe5602a1059f08580bd10d1110f11035117c10630f640ec30c;
    decBuf[778] = 256'h3a0b6f09bf07c60562037e00c5fd97fabdf627f4bdf29af036f091f0e3f0c3f1;
    decBuf[779] = 256'h8ff2c4f3ddf442f6e3f76cf937fbe7fc70fe3b00700118024b02c001ee0047ff;
    decBuf[780] = 256'hdefcfaf97af63ff243eea3ea68e68fe302e2a8df84dd93dbced933d853d70fd7;
    decBuf[781] = 256'h4cd746d9aadb32df7de231e753ea4feeeef12af626fabdfc07002b0255036504;
    decBuf[782] = 256'h1204c803740248003dfe51fbd1f787f4adf00eedc3e9c4e6d3e40ee3bce271e2;
    decBuf[783] = 256'hb5e2eae373e5d8e679e8e3ea23edc3ef3df27df41df7e2f8d9f923fadff9a2f9;
    decBuf[784] = 256'hf9f860f8d5f7abf738f789f62ef52ff3cbf0e7edf6eb7ce9e1e76be69fe5e6e4;
    decBuf[785] = 256'haee415e443e4c2e4cee54ee719e945eb50ed3cf0f4f26ef5aef7b9f995fbcafc;
    decBuf[786] = 256'h72fd3ffd57fcdcfa11f961f7d8f5d9f4f1f3caf2bdf184f0b4ee88ec7deaa1e8;
    decBuf[787] = 256'hf1e6d8e53fe56ee5ece5ace615e773e790e7aae7c2e703e865e806e99de927ea;
    decBuf[788] = 256'h5cea8dea43eab0e9d8e8d6e756e68be45fe2bedf90dc6cdab4d7efd554d409d4;
    decBuf[789] = 256'h4dd407d5afd514d759d828dad8dbd1dd35e075e216e544e843eb50f084f6afff;
    decBuf[790] = 256'haa0af4170a282c37de48c254915f66699c67fc658e6129582e4dd842213c9733;
    decBuf[791] = 256'h0b2e00293f266a201c1b27129c0968fd09f2bfe4d0dbb0d34eccf7ca2fccbbd1;
    decBuf[792] = 256'hcbd8e1e246ecd1f495fca0010b088c0a560e671088136116f718511b9a1cc41d;
    decBuf[793] = 256'h891f24212f231b26d428022cdc2f7b33d535d338fe39583aab3aca3976384237;
    decBuf[794] = 256'h99366636f1366d38d239733b8c3c253d3d3c6d3ac637e3333a2fd82adc263422;
    decBuf[795] = 256'hd21dd61936160a11370c9506c3ff58f9d7f1c8ea32e607e23dde2cdc8cdbfada;
    decBuf[796] = 256'h75daeeda36dc61dd25df0ae289e5c4e9c1ed60f19cf598f937fd820080037205;
    decBuf[797] = 256'h8106d4068906bd050405cc04330461043704c4031503b90118001ffe43fc0efb;
    decBuf[798] = 256'h66fafffafdfce9ff6803a4077d0a1c0e850fce106a105b0f1b0de509e606a002;
    decBuf[799] = 256'ha3fefbf999f579f008eda6e8aae40ae1cfdcf6d956d6fdd3d9d13dd24cd330d6;
    decBuf[800] = 256'hb0d9ebdde7e190e6f2eaeeee96f3f8f718fdeb018d07db0cad110f16e818751a;
    decBuf[801] = 256'hee1aa5197b1801161d139e0f440d450a5408da053f043402e000abff92fe2dfd;
    decBuf[802] = 256'he9fb16fb56fa33fad1fa0efc31fed2004c0330062108e609380a830a3f0a010a;
    decBuf[803] = 256'h5909c00891081308a00737075a061e05f703ea02b001de006a004800a6007001;
    decBuf[804] = 256'hc3026504ce060e09af0b280e6810de113213eb132314f013c213ef122f123b11;
    decBuf[805] = 256'ha00f170e800b06092206a30258ff35fd7cfa4ef72af572f2adf06deef8eca4eb;
    decBuf[806] = 256'heaeab2eae5ea70ebefeb62eccaec69edf8ed4cef91f060f210f499f5fef689f7;
    decBuf[807] = 256'h08f8e1f7bef720f757f6a0f5caf4c8f3d3f2f6f1f3f0ffefe3ee23eebaed1ced;
    decBuf[808] = 256'hffec19ed31ed47ed82ed70ed5fed6eed61ed6deda4edaeeda5ed7ced0bed79ec;
    decBuf[809] = 256'ha1eb9eeaaae98de834e793e50ae4d9e1cedff2ddc6dbbbd9dfd7aad691d55ed5;
    decBuf[810] = 256'h30d55ad51ad6c8d6e5d73ed926daa1db06dda8de30e0fbe1ace3a5e581e731e9;
    decBuf[811] = 256'h2aeb7eecb3ed5beef4ee7fef55ef7cef59effaeeddee8fee48ee07eecceddeed;
    decBuf[812] = 256'h0eee1dee45ee6aee49ee17eec5ed4cedb9ec7eec25ecf4eb03ec2bec50ec9dec;
    decBuf[813] = 256'hbbecd6ecefecf6ec19ed5ded9dedf8ed4dee84ee7aee5eee04eeafed78ed5aed;
    decBuf[814] = 256'h51ed7aed81ed5fed1aed91ecbaebf0ea39eac3e904eadbea18ec93ed5eef93f0;
    decBuf[815] = 256'h1bf21af302f4d5f448f5f6f5d4f62af744f72cf76af6b3f5ddf4a1f3cef2c2f1;
    decBuf[816] = 256'hcef0b1efa4ee6aed98ecd8eb6feb50eba6ebf4eb6becd7ec12ed24ed14ed22ed;
    decBuf[817] = 256'h15ed6aedf9edaaeeafefa3f041f15ef10ff13af08aee56ed3dec3eebb3ea89ea;
    decBuf[818] = 256'h16ea67e90be80de6a9e36ae1f4df18de5fdd97ddcaddb2de84df44e038e1d6e1;
    decBuf[819] = 256'hd9e213e437e66de921ee45f64100550cf41aa52c4b3d6e4c315a206300687a69;
    decBuf[820] = 256'h7365595f5d55f84b6d43a93b9e363330082c3e286b23881c48144c0a37fed8f2;
    decBuf[821] = 256'h76eb10e267de4bdd4edee3e264ea78f303fcff05640f7e150a1b111ed120a621;
    decBuf[822] = 256'he4209521f4206320de1f661fd31f701fca1f1c2092216e239a253b28b42af42c;
    decBuf[823] = 256'h6a2ebe2f77309031f53296348f367b39fb3c45404443c3461d49414ba44b4a4b;
    decBuf[824] = 256'h0a49d445fa41523df038d033fd2e5b290d243b1f98194a14170e41086f01dafc;
    decBuf[825] = 256'h04f73af3c8efa7ec15ec88ea00eb92eaf6ea05eca1edacef20f36bf644faedfe;
    decBuf[826] = 256'h0e02e7047d07f5073e09da083509e3080208be078107b907ec0777084a09090a;
    decBuf[827] = 256'h430b160c890c7d0ddc0df90db00eb50f3511661306168018641b1d1ee11fd820;
    decBuf[828] = 256'h8d20c11f951d5f1a8616e612ab0eae0a0606a401cbfe2cfbe1f7e3f42af266f0;
    decBuf[829] = 256'hcbee55ed89ec42ed5bee26f0cdf2fbf5d5f974fdb00189042808820a800d3910;
    decBuf[830] = 256'h671366161e19981b331da91eed1eaf1e261d5b1bb4183b16fb13851231117810;
    decBuf[831] = 256'hb010af11f4121a14c115d916d8176318e2185519491a231c0f1f56237628482d;
    decBuf[832] = 256'hea32b436c6386639b1371134e52eb228dc228e1d5b173013ea10780d970bbe08;
    decBuf[833] = 256'h3107c8057f045503fa024c032d048105ac074d0a310ed9127b18c91d3b219d25;
    decBuf[834] = 256'h5227e02867281f276624ed21091fc21ac6162613fa0d2809c604ca002afdc1fb;
    decBuf[835] = 256'h79fadcfaa1fce0fe8101fb033a06db08a00a3b0c1b0d6f0ead0ee50eb20e270e;
    decBuf[836] = 256'h540d480c820a56084b06d7028dffd8fa76f67af2d2edb0ead8e74ae6e1e473e4;
    decBuf[837] = 256'hd7e431e528e673e6c7e7fce885ea50ec7bee1cf196f3d5f5e1f7bdf96dfb15fc;
    decBuf[838] = 256'h48fc1afc9bfb8ffa55f92ef888f66ff50af469f250f1ebefa7ee80ed73ecc5eb;
    decBuf[839] = 256'he7eae5e936e959e8c9e77be7c2e72ee8dfe8b5e97eea35ebdbeb1cec2fec65ec;
    decBuf[840] = 256'h75eca2ece4ecf1ece6ecdcec9cec62ec5aec46ec72ecbbecedec1aed44ed1eed;
    decBuf[841] = 256'hfcece9ecb6eccbec10ed50edcbed48ee9aeee3ee41ef65ef86efcceffaef34f0;
    decBuf[842] = 256'h77f093f0abf0d1f0caf0c4f0d5f0c5f0caf0f9f018f156f1b1f1edf124f242f2;
    decBuf[843] = 256'h15f2a9f107f119f0fdeea3ed02ec79ea14e9cfe7a8e6e9e53ae59ce446e42ce4;
    decBuf[844] = 256'h14e455e490e4e9e45be5c2e53ae6cde608e761e7d3e7ffe75de8b1e8d2e8f0e8;
    decBuf[845] = 256'h1ee905e9e0e8bde860e802e8dee77be738e744e74fe7bde77de868e945ea81eb;
    decBuf[846] = 256'ha8ec68ed5ceebbeed8eef2eeabee13ee8aede9ec27ec3beb1feac5e881e7b1e5;
    decBuf[847] = 256'h86e37ae19edf73ddfddba9daf0d947d9aed8ddd807d9e0d803d962d97fd9cdd9;
    decBuf[848] = 256'h44dab0da88db8bdcc5dd40df0be1bbe295e514e940ee74f4f4fb080504104e1d;
    decBuf[849] = 256'hd0296f384342334b5253cc547553cb4f3f4a3043ef3a2b33202e8a29b423ea1f;
    decBuf[850] = 256'h781c1718d311fe0ba803e4fbd0f2b6ec2ae727e612e792e964f0d0f6fbff8508;
    decBuf[851] = 256'h49105917191a991cd71b271b06182d1597124c0f030ed90cc90b770b570c9b0c;
    decBuf[852] = 256'hd00d590f24115013f1156a184e1b071e802009245427522ad22d0d32e6348538;
    decBuf[853] = 256'hd03bf33d1e3fc33ecd3dc13b4d3812341630642a16254420e21bc216f0118e0d;
    decBuf[854] = 256'h6e089b03f9fd2ffa5df5fbf0ffec68ea0ee8c6e662e608e65ae63ae706e83be9;
    decBuf[855] = 256'h54ea53ebdeeb05edc4edb9ee96ef26f074f0bbf04ff0c6efddee00ee37edb4ec;
    decBuf[856] = 256'h6dec57ec92ecc8ec5aede3ed84ee47ef32f04ff1f5f27ef4aff64ff9c9fb52ff;
    decBuf[857] = 256'h9c0276060c09570c7a0ea50f4a0f540ede0cf209720628034effaffb64f841f6;
    decBuf[858] = 256'h88f30ff1cfeec4ece8eab3e99ae867e896e8bde9afeb13eef8f077f4b3f8affc;
    decBuf[859] = 256'h4e00a802a7059807a808fa08af08f3083a08020869073a07bc0649069b053c05;
    decBuf[860] = 256'hac045e041604010414046e040005ff053907b408190aba0b430d420e2a0ffd0f;
    decBuf[861] = 256'hbd106b110912991250139713ad137213ad128e113410930e0a0da50bbd0aeb09;
    decBuf[862] = 256'h780955097409cb09810a570b5a0c940dbb0e1410591180128c13c614ed154617;
    decBuf[863] = 256'h2e185519c819eb190e19d11702165b13e110fd0d7e0a240825056d02f3ff58fe;
    decBuf[864] = 256'h4dfc71fac0f838f739f6f4f421f4aef346f3e7f2caf218f360f3ccf355f4d2f4;
    decBuf[865] = 256'h23f550f578f56cf561f543f53af521f50af5daf4a2f45ef41ff4d4f3b6f39bf3;
    decBuf[866] = 256'h93f3a9f3bef3d1f3edf3fcf3f7f3d1f399f346f3e3f286f249f212f2f4f1ebf1;
    decBuf[867] = 256'h04f20bf212f2fff1e3f1bff196f185f175f17af176f162f13cf104f1c0f06ef0;
    decBuf[868] = 256'h21f0efefafef65ef1fefbaee27ee4fed86ec9bebbeeaf4e972e9fbe8bae87fe8;
    decBuf[869] = 256'h91e8a1e809e981e934ea0aeb0cec00eddeede1eed5efb2f0b5f1a9f205f4a6f5;
    decBuf[870] = 256'hbff624f868f93bfaaefa17fb76fb92fbe1fb28fc69fccbfcddfcedfcdefc81fc;
    decBuf[871] = 256'h2cfcc9fb36fbacfa2ffa7df9d6f83ff8b6f738f7e7f680f63df631f610f62ef6;
    decBuf[872] = 256'h6ef6d9f65ef722f8d9f880f96dfa0cfb9bfb1efc95fc7ffc6bfc12fc5ffb8afa;
    decBuf[873] = 256'hc0f9a1f894f7a0f684f52af4e6f2bff165f021ef4eeedbedb8edd8ed67ee1eef;
    decBuf[874] = 256'hc5efb2f090f120f2d6f21ef35ff372f319f3e8f29ef25bf237f258f28af2eef2;
    decBuf[875] = 256'h82f30bf464f475f42bf462f35ff2e0f07befd9ed31ed98ecc6ec45ed05eef9ee;
    decBuf[876] = 256'h97ef27f0d8ef32ef19ee73eceaea1fe96fe7e6e5e7e4ffe381e35ae337e357e3;
    decBuf[877] = 256'h3ae320e3d9e26de20be2b1e1a1e1cde146e239e3b9e4eae68be96eed17f2f9f8;
    decBuf[878] = 256'h65ff90088b13e11df6295535b73c1c46364c8a4f884ec84bf245203fdf365331;
    decBuf[879] = 256'h442aae252e23641f531d311a5917b0124e0e2f095c04faff21fd94fbfdfcfcff;
    decBuf[880] = 256'h09053c0bbd12cd1938206324a926f82518241b206a1a1c154910e70b0f098107;
    decBuf[881] = 256'h090751080a0b380e1212b115ed19e91d8821d324ad284c2ca62e7f321f366a39;
    decBuf[882] = 256'h683ce83f414265448f45ea454f44ae417f3ea63afd355b300d2b9b273a233d1f;
    decBuf[883] = 256'ha71c4d1a2918381628158d1317123b10100e040ca0090508fa05a604ed034403;
    decBuf[884] = 256'hab02da020403dd020003e1025102ce01f90083ff1efe20fc44fa18f80df631f4;
    decBuf[885] = 256'h77f35ff22cf25af22df339f4b9f584f7b9f842faa7fbebfc12fe1fff59008001;
    decBuf[886] = 256'hd9027a0473064f087b0a1c0d950f7a126b147b15cd15ed141113ee0fef0c7009;
    decBuf[887] = 256'h250627036e005fff68feb3fef7feb0ffe8ff810053007d00570034005300e300;
    decBuf[888] = 256'h0202a903a2050608450a510c2d0e610f9a0fcd0f410f1b0e5b0d210c4e0b420a;
    decBuf[889] = 256'h9309b608ed0736078f062306e805fa056c062c0717087309b70a330c980ddc0e;
    decBuf[890] = 256'haf0f6f10d710b810d41086109e10b310ee106b11dd1144126d124812cf11fc10;
    decBuf[891] = 256'hf90fbf0e980dd90c700c900c1f0d0a0e660f08119112f613dd1404167716e016;
    decBuf[892] = 256'h001756177017b717cd17b9178417121752163315d91338123f10630e370c9609;
    decBuf[893] = 256'h1d07dd04d202f600cafe54fd88fc54fbabfa78fa4afa20fa93fab6fad5faf2fa;
    decBuf[894] = 256'hd8fa91fa25fa9bf9d7f820f84af781f6caf524f58cf403f462f39ff2e9f142f1;
    decBuf[895] = 256'h54f0b6efedee6aee53ee68eea3ee20efd3ef79f067f145f20ef3c5f33bf4a8f4;
    decBuf[896] = 256'he2f4adf47cf432f4d5f398f38df383f38cf3a5f39df389f36af32cf3f2f2bdf2;
    decBuf[897] = 256'h64f20ff296f1e3f00ef044ef59ee7cedb3ecfceb26eb5dea72e9d4e80ae888e7;
    decBuf[898] = 256'h40e72be73ee774e7e6e712e855e8aae80de985e938eaafea46ebcfeb05ec36ec;
    decBuf[899] = 256'h62ec55ec49ec6aec4cec42ec5bec63ec77ecc9ec16ed84ed26ee92eef4ee71ef;
    decBuf[900] = 256'he3ef68f0e5f016f142f185f160f16bf19df1b9f103f285f202f394f31ef4bff4;
    decBuf[901] = 256'h2bf5b4f50df63ef64df625f6d0f56df5f5f4a3f495f487f4acf4e3f401f5f7f4;
    decBuf[902] = 256'hdff48cf413f460f35bf267f14af0f1ee09ee8bed18ed3bed99edf0ed3eee26ee;
    decBuf[903] = 256'h8feddeec09ec06eb57ea38ea1bea9eeaa3eb97ecf3ed94efadf012f2faf278f3;
    decBuf[904] = 256'hebf30ef4aff359f3d6f260f2c8f18df110f1bff075f0fdef8bef06ef66eeceed;
    decBuf[905] = 256'h1eeda7ec0fecd5eb7beb4aeb1eebf6eaeaeac9ea97ea69ea1feac5e970e9f7e8;
    decBuf[906] = 256'h85e81ee8a6e755e728e71be73fe78ce7d2e724e887e8e5e83ae9c9e952eaf3ea;
    decBuf[907] = 256'h0cec19ed99ee64f00bf339f613fabbfe5e04300b9b111b192b209626c12a8b2e;
    decBuf[908] = 256'h9c303c31872ff12ca629cd252421031e2a1b94182a17e215b714f312b310120e;
    decBuf[909] = 256'he40ae5072d05b302180163013f03e605ca09720ed412ad154c19c51957192d18;
    decBuf[910] = 256'hb31586118a0dea099f067c045103f70292049d06110a4d0e4912e9153319571b;
    decBuf[911] = 256'h0f1e1f1fba209a2166221f23382437257c264e275b28c428a428db275326e923;
    decBuf[912] = 256'haa21731e9a1a0318b91495126b11a60f540f090f4d0f100f480f150f8a0e630d;
    decBuf[913] = 256'h090cc50af50845072c06c704e003b902ac01b800dbffd8fe29fe8bfd35fde7fc;
    decBuf[914] = 256'h9ffcb5fc7afc21fcd0fb2dfb96fa0dfa8ff93ef96af9c8f94dfa12fb95fbdcfb;
    decBuf[915] = 256'hf2fbb7fb81fb30fb04fbf6fa02fb39fb93fb31fcf4fc13fe6cff0e0107035b04;
    decBuf[916] = 256'h0b06b3064c07c106ef059504f4026b01a0ff6bfe53fdbafce8fc12fdd2fd80fe;
    decBuf[917] = 256'h1fffaeffc8ffb1ff9bff87ff99ff0b00e80005025e03000518067d07c2089509;
    decBuf[918] = 256'hbb099809fa08f707bd064205dd039902c6015301ea00cb00e700cd00b5007500;
    decBuf[919] = 256'h610073008300af000d017a01e101240279029a02900287025e02290215022702;
    decBuf[920] = 256'h4f029c0215038603ee0330043d0432040004ad0360031a03ed02d402eb022803;
    decBuf[921] = 256'ha40345040805f305d00699071c08c2085a09e309840a1b0bcc0b430caf0cea0c;
    decBuf[922] = 256'hb40c630cde0bf60a180aa3083e079c05a303c70117001efecafc19fb01fa02f9;
    decBuf[923] = 256'h1af847f7d4f6b1f692f675f65bf614f6a7f51ef5a1f4eef348f3b1f24ef2f5f1;
    decBuf[924] = 256'ha4f178f14ff143f122f1dcf09cf031f0caef87ef63ef6eefa0ef16f0c9f06ff1;
    decBuf[925] = 256'h32f21df3faf3fdf4f1f5cff65ef715f88cf8cdf8e1f8f2f803f92ff957f994f9;
    decBuf[926] = 256'hf7f91ffa43fa38fab6f915f927f80bf7b1f56df446f339f28bf1aef01ef0cfef;
    decBuf[927] = 256'h29efbdee5bee02ee90ed46ed03eddfecbeecb4ecbdecd6ecfbec47edb5ed1cee;
    decBuf[928] = 256'hafee39ef6eef9fefaeefa0efacefe3ef29f0b2f063f139f23bf330f40df5d6f5;
    decBuf[929] = 256'h8df604f770f7f9f72ff8a1f808f99bf924fac5fa31fb94fbc9fbd9fbe8fbf6fb;
    decBuf[930] = 256'he9fbf4fb12fcf7fbbdfb7afbf1fa68fac7f9d9f83bf871f7eff678f637f64bf6;
    decBuf[931] = 256'h80f6f2f63cf7b4f747f8a9f802f953f9bbf9fdf96bfa97faa4fa98fa77fa45fa;
    decBuf[932] = 256'h05fabbf975f923f9c0f862f80df8c0f78ef773f75af735f705f7b3f650f60df6;
    decBuf[933] = 256'hd1f5c6f50cf670f603f7b4f72bf897f8aaf8bcf88cf842f8fff7c2f78bf759f7;
    decBuf[934] = 256'h2cf702f7b0f663f61df6b9f576f551f530f526f52ff5f6f4b2f43cf489f384f2;
    decBuf[935] = 256'h8ff134f0efee1cee10ededeccdec23ed0feeeceeefefe3f081f111f25ff277f2;
    decBuf[936] = 256'h61f226f214f245f2acf225f3f8f3fbf4eff5ccf6cff77df89af9a7fae1fbb0fd;
    decBuf[937] = 256'h60ffca01ae0466074a0be90e34123215b2180c1b541cb81c5d1c0b1c951ab918;
    decBuf[938] = 256'h09178015b51389111410c00e0f0df70b920aaa092c0905092809c6098f0ae30b;
    decBuf[939] = 256'h840dee0f2e12ce1448178819281ced1d881f68203421f7204e204f1f0b1ee41c;
    decBuf[940] = 256'h241c751b561bac1bfa1b711c091d431d551d251ddb1c981c741c691cc31c301d;
    decBuf[941] = 256'hd21d951e4b1f2120ea20a12148220a23592341235623f4225322bc21e4201b20;
    decBuf[942] = 256'h641f8e1e8c1d971cba1b441a7918c916601420127f0f060d6a0bf50929096f08;
    decBuf[943] = 256'ha808db08c209950aa20b960cb20dbf0eb30f91102011d7117d12be12f912e712;
    decBuf[944] = 256'h7612d311ba10140f8b0dc00b94098907ad05fd03e402e501fd00d300fa001d01;
    decBuf[945] = 256'hbb0184026f03cb0410063607dd08f509f40adc0b060c2d0c0a0c2c0b2a0a3509;
    decBuf[946] = 256'hda0738062005bb037602a301e3007b005b007800c6003d01d401ac0276039504;
    decBuf[947] = 256'hee0590071909e40a940c1d0e1c0f04108210a810cb10ac101c10990fc30ec10d;
    decBuf[948] = 256'hcd0cef0bec0af8095a09ca084808d1073a07ff06c90698068a067c0670067b06;
    decBuf[949] = 256'h8506a106eb0631077107cb07f00711080708d9078f074907d2064006b7053a05;
    decBuf[950] = 256'ha7041e04c5039403a303cb0307048004f2047705f4056606ea068b074e083909;
    decBuf[951] = 256'h560a620b9c0c6f0d2f0edd0efd0ea60e240e4e0dd80b730a750899066d04f802;
    decBuf[952] = 256'h1c01e7ffcefe35feaafd2cfd6cfcbefb1ffb1dfa29f98af8c1f773f72cf716f7;
    decBuf[953] = 256'h02f7cdf67bf6f7f57af5c7f421f489f300f383f211f26ff103f1a0f023f0f3ef;
    decBuf[954] = 256'hc6efd4ef10f073f006f1def1e1f21bf496f595f6daf701f9c0f929fac7fa57fb;
    decBuf[955] = 256'hdafb50fc91fca5fc6ffc1efc5efba7faa2f9aef891f738f650f529f4d0f2e8f1;
    decBuf[956] = 256'h15f109f0a0ef02ef72eef0ed79ed0ded83ec2aecd9ebcaebf2eb5fec01edefed;
    decBuf[957] = 256'h0cefccefc0f05ef1b4f103f2bbf14ff1edf04cf0e0efa5ef93efe5ef69f00af1;
    decBuf[958] = 256'hcdf184f22af396f3d1f3e3f3d3f3e1f30af446f4d5f45ff523f6daf6b0f779f8;
    decBuf[959] = 256'h30f9a7f9e8f9fbf97ef9ecf814f811f763f685f52ff5adf465f424f49bf31ef3;
    decBuf[960] = 256'h6bf2c5f102f180f0d9ef99ef36ef25ef35ef61efbfef5cf01ff10af227f333f4;
    decBuf[961] = 256'he2f4fef5bef66df70bf89af81df994f900fa14fa02fad1f987f92af9bcf838f8;
    decBuf[962] = 256'hdef74cf7c3f669f6d7f54ef5f4f483f41bf4f3f3b7f396f38cf35ef314f3cef2;
    decBuf[963] = 256'h45f2bbf11bf158f0a1effbee63eeb3ed3cedd0ec47ecedeb5bebd2ea78eae6e9;
    decBuf[964] = 256'h35e9bfe852e8f0e7bbe7aae77ee7a6e79ae7bbe7ede752e8cae89de966ea1deb;
    decBuf[965] = 256'hc4eb5bec96ecefecffec0eed36ed42ed63ed95edc3edeced12ee0beef8edd1ed;
    decBuf[966] = 256'h84ed21eda9ec37ecd0eb8deb81ebb8eb3aecfeece9ed45ef8af005f26af3aff4;
    decBuf[967] = 256'h81f58ef6f6f655f772f758f740f72bf717f770f7c2f70bf869f88df898f8a2f8;
    decBuf[968] = 256'h99f8b2f813f9a7f97efa81fbbbfce2fd3bff8000a70100034504c0058b07c008;
    decBuf[969] = 256'h490aae0b950cbc0d7c0ee50e830f13106110d81019117b11b011e111f011fd11;
    decBuf[970] = 256'hd911a2115c111c11c110b510c01006118f116712301350145c1550162e173018;
    decBuf[971] = 256'hdf187d19d319561a9d1a091b1d1b521b631b541b2c1bbf1aff191419f7179e16;
    decBuf[972] = 256'h5915321426137712d9114911fb10b4109e10d9103211a41164121b13c1135814;
    decBuf[973] = 256'hbb14f0142115f514971412144d132e12d410330faa0d790b6e0992075d064405;
    decBuf[974] = 256'h45041704ed03c703e903ca03ad03c703af03c50300045904ab04f4040205f604;
    decBuf[975] = 256'hbf0465041004ad033403e3027c021e02c9017c013601e4008100090077ffedfe;
    decBuf[976] = 256'h70fefefdd2fdfafd4ffec8fe5affe4ff3d008e00bb00c800bc009b007d002b00;
    decBuf[977] = 256'hdeff70ff08ffabfe56fe1ffe15fe0cfef3fdddfdacfd68fd16fdc9fc97fca0fc;
    decBuf[978] = 256'heafc58fdfafd92fe42ffe8ff55008f00a100910065003d00180023005500a700;
    decBuf[979] = 256'h0a018301b401e001d201ae0177016d018801e30181021803c9039f04f5047705;
    decBuf[980] = 256'h8f057a051705be046d040604dd03b903c403e203100439047c04aa04b204ab04;
    decBuf[981] = 256'h5104cc0307031c020001f3ff45ffa7fe17fec8fd52fde6fc35fc8ffbf7fa6efa;
    decBuf[982] = 256'h15fac3f9b5f9ddf919fa66fad4fa3cfb99fb06fc6efc96fcd2fcf3fcfdfcd0fc;
    decBuf[983] = 256'ha6fc45fccdfb5bfbb9fa4cfac3f98df97df98cf9cff924fab3fa15fbb6fb22fc;
    decBuf[984] = 256'habfc05fd76fda3fde5fd22fe2dfe37fe2efe15fef0fddbfdaffdaafda5fda9fd;
    decBuf[985] = 256'hb6fdc2fdbefdb5fd95fd55fd03fda0fc28fcb6fb4ffbf1fab5fa94fa8afaa5fa;
    decBuf[986] = 256'hcefa12fb52fb8bfb93fb8cfb6dfb2ffbe5fab3fa60fa29faf7f9b8f96df927f9;
    decBuf[987] = 256'hc3f865f841f820f83ef86cf8b6f8fcf83cf975f9c8f915fa6ffadcfa43fb86fb;
    decBuf[988] = 256'hc3fbcefbb0fb94fb6bfb46fb08fbcefa6dfa0ffaa2f93bf9ddf888f867f849f8;
    decBuf[989] = 256'h2ef815f80df8f9f7e6f7ecf7f1f7fff703f816f828f83ef869f8baf81df995f9;
    decBuf[990] = 256'h07fa8cfa2dfb99fbd4fb2dfc3dfc2ffc21fce5fb82fb3ffbd2fa6afaf2f980f9;
    decBuf[991] = 256'hdef847f86ff76cf6bef5e0f417f460f319f3d8f213f349f3baf33ff498f40af5;
    decBuf[992] = 256'h54f561f586f591f5aff5dcf537f68cf6d9f61ff74df755f72ff7e4f68af61df6;
    decBuf[993] = 256'hb5f558f51bf5e4f49ef44cf4fff3a5f338f3d1f28ef239f218f20ef217f261f2;
    decBuf[994] = 256'he3f284f347f432f50ff6d8f65bf7d2f713f875f8cef81ff9a4f945fadcfa66fb;
    decBuf[995] = 256'h2afcadfc53fdebfd74fecdfe1fff68ff91ff9dffbeff04006800fb00ac018202;
    decBuf[996] = 256'h840378045605e605d1063007f907b0085609190a040be10baa0cca0d8a0ec30f;
    decBuf[997] = 256'hea10aa11e412b713771425158415da15f415dc159c1561154f15fe140c153415;
    decBuf[998] = 256'ha21561164c172a182d19211afe1ac71b7e1c241de71dd21e701f73202121ff21;
    decBuf[999] = 256'h8f2245238d23f9233424fe23cd238423f0228e223522c321b4218c2168218921;
    decBuf[1000] = 256'ha721b021ea210022f9210022d8218b2112218020f71f9d1f6d1f401f691fa51f;
    decBuf[1001] = 256'hb01fe21fb51f491fc51e001e151d371c351b411aa219d918ee17111747162815;
    decBuf[1002] = 256'h6814ba13dc12c01271122a121412da118011ee103d10970fd40e1e0e480d7f0c;
    decBuf[1003] = 256'hc80b210b8a0ad9093309c7083e08e40793072c0799063706b90548051b05f304;
    decBuf[1004] = 256'hcf04f004fa04f1040a05110518052b051a05ec04b3044304b1034f03d1026002;
    decBuf[1005] = 256'h5102440250028702a502ae02a6028f0251021702b6013e01cc004700caff58ff;
    decBuf[1006] = 256'h0effe6fef2fe13ff6dfff3ff700002016401be01ce01dd01cf0193015c012a01;
    decBuf[1007] = 256'hfc00d300ad009900860080007b0077006a005e003f001800e0ff9dff4afffdfe;
    decBuf[1008] = 256'h8ffe28fee5fdc1fdccfd12fe76fe09ffbaff31009d00ff003501450154017c01;
    decBuf[1009] = 256'hb80105027302f8027503e70331047404980477045904f5037c03ca02f4012b01;
    decBuf[1010] = 256'h3f0062ff5ffeb1fdd4fc44fcc1fb4afb0afba7fa72fa41fa15fad2f97df904f9;
    decBuf[1011] = 256'h72f8c1f71bf758f6d6f52ff5eff4b4f4a2f4d3f41cf5aff512f68ff600f70ff7;
    decBuf[1012] = 256'h02f7c5f64cf6daf556f5d9f487f45bf44ef442f44df443f427f41ff4eaf3c8f3;
    decBuf[1013] = 256'hc2f3c7f300f461f4daf44bf5b3f5f6f5e9f5c8f546f5c9f417f470f3d9f250f2;
    decBuf[1014] = 256'hf6f1c5f1b7f1c4f1d0f1f1f1d3f181f11ef18bf002f0ccefbcef05f099f070f1;
    decBuf[1015] = 256'h3af259f3ccf37bf49af47df4fbf384f3c1f2d6f138f1a8f05af072f087f0eaf0;
    decBuf[1016] = 256'h43f194f185f178f10bf186f0e5ef4eefc5ee6bee1aee0bee19ee3dee74eef6ee;
    decBuf[1017] = 256'h73ef05f08ff030f19cf14cf294f200f362f3bbf3ecf318f4f0f3b3f37cf30ef3;
    decBuf[1018] = 256'hc5f2b7f2abf2ccf226f37bf3b2f3f8f3eff3d6f3a2f33bf3d3f290f254f233f2;
    decBuf[1019] = 256'h65f292f2fef2a0f30cf495f413f523f514f5ecf47ff4faf3a1f34ff323f34bf3;
    decBuf[1020] = 256'ha0f32ff4e0f486f5c7f502f685f5f2f41bf4def20cf2fff051f031f04ef068f0;
    decBuf[1021] = 256'hdff076f1fff159f2aaf2d6f2c9f2bdf2b2f294f29df284f27df284f24bf208f2;
    decBuf[1022] = 256'hb6f127f176f0d0ef0def56eee0ed48edbfec42ecf0eb89eb61eb0cebebeae1ea;
    decBuf[1023] = 256'hd8ea01eb27eb65ebbfeb45ece6eca8ed93ee71ef3af0f1f068f1a9f1bcf1aaf1;
    decBuf[1024] = 256'h9af1a9f1b6f10bf284f2f6f298f32ff492f4ebf41cf50df500f5f3f4fef444f5;
    decBuf[1025] = 256'hcdf5ccf606f82df987facbfb46fd45fe2dff00000c01bb0198029b038f042d05;
    decBuf[1026] = 256'h3006240701080409f809d60a9f0b560ccd0c0d0d210d0f0dff0cd30cc50cd10c;
    decBuf[1027] = 256'h080d3a0d8d0df00d4d0ed30e730f361021117d12c2133d15a2164318cc19cb1a;
    decBuf[1028] = 256'h561bd51bfb1bd81bb81b9c1b4d1b651b7b1b671b791b481bc31a231a6019a918;
    decBuf[1029] = 256'hd3177d172f174617de17b618b819f21a191cd91ccd1d2c1e821e681e211eb51d;
    decBuf[1030] = 256'h041d5e1cc71b161b701a041a7a192119af180d181f1742163f150514de121e12;
    decBuf[1031] = 256'h2a11cb103b10b90f420fd60e250eaf0dec0c350cbe0b520bf00aba0a8a0a5d0a;
    decBuf[1032] = 256'h350af909960938099a08d80755077f06f0056d05c7042f04cd035003be025c02;
    decBuf[1033] = 256'hbb014f01ed0070003f00130005002a0061009300c000c8008500fcff24ff21fe;
    decBuf[1034] = 256'he8fc15fc55fbecfacdfa23fba6fb4cfce3fc1efd0cfdbbfc19fc56fb9ffa29fa;
    decBuf[1035] = 256'he8f9fbf955fae7fa98fb3efcd5fc37fd25fdd4fc14fcf5fa9cf957f830f724f6;
    decBuf[1036] = 256'h75f516f5faf4dff427f568f5a2f5d8f54af6b1f60ff77cf7c6f7eef7c9f766f7;
    decBuf[1037] = 256'heef65cf6faf5e8f518f6bbf67df79df85df90bfaebf922f99af7a1f5b5f2fdef;
    decBuf[1038] = 256'hceecabeab9e85fe855e9f6eb25efd9f33bf837fcd7ff30029e027301fafe16fc;
    decBuf[1039] = 256'h96f84cf503f4d9f233f32af435f699f8d9fa4ffc1bfdddfc54fb23f982f609f4;
    decBuf[1040] = 256'h6df2f8f0b4f0e8f152f436f7b6fa00feff00f0024b0354024900d5fc8af9b1f5;
    decBuf[1041] = 256'h1af3c0f053f0b6f0c6f1aaf49bf6caf9edfb18fd27fed5fdf5fc29fc79faf0f8;
    decBuf[1042] = 256'h8bf746f6c8f5a1f5c4f523f6b3f66af7b1f7f2f706f8f4f7e3f7f2f750f806f9;
    decBuf[1043] = 256'hf1f90dfb67fcabfd7efe8bfff3ff1300bdff3aff64fe62fd28fc01fbf4f900f9;
    decBuf[1044] = 256'h62f80cf8f2f7daf7eff703f8f1f7e1f7d2f7c5f7d1f7f2f738f878f8d3f80ff9;
    decBuf[1045] = 256'h1af924f9e4f879f812f864f78ef6c5f50ef538f4a9f3f2f2aaf26af256f244f2;
    decBuf[1046] = 256'h54f263f270f295f2b6f2fcf260f3d9f38bf432f5f4f5abf651f714f897f80df9;
    decBuf[1047] = 256'h4ef989f9bff9aef982f975f950f945f963f991f9ecf959fac0fa39fbaafb12fc;
    decBuf[1048] = 256'h6ffcacfce3fc29fd44fd5dfd64fd5efd57fd52fd57fd6efdaefd00fe4dfebbfe;
    decBuf[1049] = 256'h05ff47ff54ff5fff2dff11ffe8fee0fef5fe21ff6affc4ff31007b00be00e200;
    decBuf[1050] = 256'hed00e300b5009d0095009c00c80011017f010402a5026703ea039004fc045e05;
    decBuf[1051] = 256'h9405a40595056d051805cb045d04d9035c03c902190272010601a4006f007f00;
    decBuf[1052] = 256'hab0009018e01e7015902a302cb02ef0210031a0336034f0356037803b103e503;
    decBuf[1053] = 256'h31049f042405c4055c060c078307ef072a086008500841084e087308aa081809;
    decBuf[1054] = 256'hba09510a020bd80b670c520df10dba0e3c0f1210a2102511cb116212ec126913;
    decBuf[1055] = 256'hda1342148514a914e014ea14e114fa1410151715361552155715651561154615;
    decBuf[1056] = 256'h5015601574159c15f015a61691176e18fe18e919871a171b651bad1b971b831b;
    decBuf[1057] = 256'h721b611b531b7b1b871bea1b621cd41c761d0e1e701ec91efa1ece1ea51e511e;
    decBuf[1058] = 256'hd81da71d7b1d6d1dda1d5f1e241f0f20ec207c21ff21462230221d229f21ed20;
    decBuf[1059] = 256'h7620b31ffc1e861eee1d3e1df61c8a1c281cf31bc21b781b351be01a511aef19;
    decBuf[1060] = 256'h4e198c1809189217fb1699163f16ee15c2157f155b15661548152c152415f014;
    decBuf[1061] = 256'h96144114b21302135b12c41113119d100510a30f6e0f3d0ff30ecb0e5e0ed90d;
    decBuf[1062] = 256'h5c0da90cd30b440b8d0ae709a60944093209420951099409d009db09d109a409;
    decBuf[1063] = 256'h2809630878075b064f051504ee02e101ed00100047ff90fe19fed8fd9dfd8bfd;
    decBuf[1064] = 256'h7bfd4ffd0cfdb7fc28fc9ffbdafa58fa82f9f2f8a4f82df8c1f786f72df7fcf6;
    decBuf[1065] = 256'hd0f6a7f69bf690f69af6c8f6f1f626f764f77cf784f78bf778f75cf757f740f7;
    decBuf[1066] = 256'h33f71ff7ebf689f611f67ff5f5f478f407f4bdf395f370f339f31bf3dbf281f2;
    decBuf[1067] = 256'h44f2e1f183f147f1e4f086f019f0b2ef39efe8ee81ee74ee80eeb7ee25efc7ef;
    decBuf[1068] = 256'h8af075f152f21bf306f4a5f434f5b7f5fef514f627f616f6a4f55af5fcf4a8f4;
    decBuf[1069] = 256'h71f467f482f4ccf426f57bf5c8f50ef617f630f637f631f643f66bf6a3f6f6f6;
    decBuf[1070] = 256'h6ff7e0f765f8e2f854f980f98ef951f9d8f846f86ef7def627f6b0f570f55cf5;
    decBuf[1071] = 256'h4af55af569f541f51df5e6f478f4f3f376f304f39df28ff283f2baf228f38ff3;
    decBuf[1072] = 256'h23f4acf405f577f5def521f676f6eff640f7c5f742f873f8bdf8e5f8c0f889f8;
    decBuf[1073] = 256'h2ff8aaf72df7bbf636f6b9f568f501f5a3f44ef4d5f384f33af312f306f33df3;
    decBuf[1074] = 256'h83f3d5f338f460f43cf4d9f310f30ef2d4f0adef53ee6ced99ecd9eb70eb51eb;
    decBuf[1075] = 256'h34eb82eb6beb80eb94eb5eebedea68eaa3e9ece876e835e821e89ee830e908ea;
    decBuf[1076] = 256'h0bebffebddec6cedefed36ee77ee8bee9deeadeebceec9ee06ef27ef59efbdef;
    decBuf[1077] = 256'he5ef09f040f04af066f07ff095f0aaf0e2f0daf0e1f0e8f0b5f093f080f064f0;
    decBuf[1078] = 256'h69f089f096f0a9f0bbf0a5f091f07ef05bf022f0fdefbfef85ef60ef14eff6ee;
    decBuf[1079] = 256'hedeec4eecbeed2eecceeddee01ef21ef61efd7ef49f0cef06ff106f2b7f25df3;
    decBuf[1080] = 256'hf4f3a5f41cf5b3f53df6baf62bf793f70bf85cf8a6f804f940f98df9d3f913fa;
    decBuf[1081] = 256'h5dfaa3fabffae8fafffa05fb18fb29fb4dfb92fbecfb59fcfcfc93fd1cfebdfe;
    decBuf[1082] = 256'h55ffdeff7f00eb007401ce0140028902e7023c037303a503d203fc033f047f04;
    decBuf[1083] = 256'hea046f051006d30689075f08ef08a6091d0ab40a3d0b970b290cb20c530deb0d;
    decBuf[1084] = 256'hc20e8c0f431048113c125913b2149a156c16e016021722179216db1535154714;
    decBuf[1085] = 256'ha9131913cb1284129912ad12bf1210131f132c1351135c137a13a71302146f14;
    decBuf[1086] = 256'hf414951501168a169c168c166016e7153515be1426149d134413f212a9126612;
    decBuf[1087] = 256'h2912c61183114711fa10b41074103a10421056108e10ff1091111b12bb122813;
    decBuf[1088] = 256'h3b134d13fc1295121c12aa112611a9105710f00fad0f580f0b0fb10e2c0e8b0d;
    decBuf[1089] = 256'hc80cdd0b000bfd094f09b1085a080c08c507af074d07d0063e06b4055b052a05;
    decBuf[1090] = 256'hfe040b0530053b051d05ef0484041d04a4031203b00256022602170224023002;
    decBuf[1091] = 256'h51026f0266023d02fa018301f1006700eaff78ff11ffb4fe8ffe6efe64fe6dfe;
    decBuf[1092] = 256'h97febcfedefe17ff2dff34ff2eff06ffcefe9afe40fed3fd6cfdf3fc61fcd8fb;
    decBuf[1093] = 256'h37fb74fabdf9e8f8e5f737f759f6c9f57bf563f579f58df5c2f5f3f51ff62df6;
    decBuf[1094] = 256'h39f65af68cf6ccf616f75cf777f76ff749f7fef6a4f64ff602f6d0f5b5f5bdf5;
    decBuf[1095] = 256'hd3f503f648f688f6c2f6e7f6fcf6f6f6daf6a1f66df63df604f6dff5caf5b7f5;
    decBuf[1096] = 256'ha7f5a1f59df599f5a4f59af58af57cf554f52df513f505f512f535f55ff586f5;
    decBuf[1097] = 256'haaf5a5f5a1f59df5a1f5c3f508f64ef68ef6c8f6b2f681f630f6cdf58af566f5;
    decBuf[1098] = 256'h87f5f5f597f65af745f822f9ecf9a2fa49fb8afbecfbfefbedfbdffbd1fbc5fb;
    decBuf[1099] = 256'he6fb18fc6afccdfc2bfd80fd8bfd81fd1cfda4fcf1fb1bfb8cfad5f92ff997f8;
    decBuf[1100] = 256'h35f8fff7eff7fef726f87bf8c8f822f977f9c4f9f6f911fa2afa31fa38fa32fa;
    decBuf[1101] = 256'h2cfa3cfa65faaffa1dfbbffbadfc8afd53fe0affb0fff1ffdeffa8ff57fff0fe;
    decBuf[1102] = 256'h92fe55fe1efe14fe0bfe24fe49fe7afeb2fed7fefafe19ff35ff44ff5cff68ff;
    decBuf[1103] = 256'h83ffaaffd8ff10006300b0001e016801aa01b701ac015201e400420080ffc9fe;
    decBuf[1104] = 256'h22fe60fd11fd9bfc5afc46fc58fc48fc57fc64fc40fc09fcd7fb84fb37fbf1fa;
    decBuf[1105] = 256'hc4faabfab3fab9fad9fa00fb2efb66fbaafbeafb34fc7afca8fcf2fc24fd64fd;
    decBuf[1106] = 256'haefd08fe5dfeaafef0fe0bff03ffedfebcfe9dfe81fe86fea7fed5fe0eff42ff;
    decBuf[1107] = 256'h72ff78ff68ff2fffddfe64fed1fd48fdcbfc39fcd7fba1fb70fb44fb1cfbdffa;
    decBuf[1108] = 256'h92fa4cfafaf9c3f991f976f97ef985f9b6f907fa54fad6fa53fbe5fb47fca1fc;
    decBuf[1109] = 256'hd1fce0fcd3fc96fc75fc6bfc62fc8bfcc0fcd4fcf4fc05fd14fd34fd74fdfdfd;
    decBuf[1110] = 256'haefeb3ffa70084014e0204037b03e70322045804a904f3045005be0507068006;
    decBuf[1111] = 256'hf10676071708da089109960a440be20b720cf50c3c0d520d650d770d870db40d;
    decBuf[1112] = 256'hc10dfe0d4b0e7d0ecf0e320f750fe20f4910c1103311b8111112831208136113;
    decBuf[1113] = 256'hf3137d141e150b16e916b217d118de198c1a2b1bba1bd41bbd1ba71b451bec1a;
    decBuf[1114] = 256'h7a1af519bf196e195f196d19a919ca19241a611a6c1a621a471afc19b6196419;
    decBuf[1115] = 256'h0119be1882184b18551870188918bd18e018da18bd187118e21731175b165815;
    decBuf[1116] = 256'haa14cd13031381123a12f9110c121e122e125b124d1229121e12d811aa119211;
    decBuf[1117] = 256'h9911a011cc11fe11211259127e129312a612951267122f12cd115511e3105e10;
    decBuf[1118] = 256'he10f6f0f080f750ec40def0cec0bf80a1a0a1809af081108bb076c07f5065e06;
    decBuf[1119] = 256'hd50510055904b3034703bd0264021302ac0169011401c70081002f00ccff6eff;
    decBuf[1120] = 256'h01ff9afe21feb0fd48fdebfc96fc49fc03fcd5fbbcfba6fb9ffb8cfb65fb37fb;
    decBuf[1121] = 256'hfffacafaa8faaefae1fa3afb8ffbdcfbfafbdefb73fbd1fa3afa62f9d2f84ff8;
    decBuf[1122] = 256'hd9f7c3f788f752f701f79af622f68ff5dff438f4a1f33ff3c2f271f244f237f2;
    decBuf[1123] = 256'h5bf292f2d8f22af3a3f3f5f33ef49cf4a8f4c9f4bff4b6f4aef4b5f4a1f49af4;
    decBuf[1124] = 256'h8af447f4f5f392f319f3a8f27bf253f247f27ef2b0f2def2f7f2eff2cdf294f2;
    decBuf[1125] = 256'h51f211f209f2f2f122f274f2d7f26af3f3f394f400f58af5bff5cff5a3f560f5;
    decBuf[1126] = 256'h0bf5bef464f428f407f4e9f3e0f3e8f3c2f3a0f374f32bf3e5f2b8f27ef267f2;
    decBuf[1127] = 256'h6ef274f27af294f28ff29cf2bff2dff21ff395f307f4a9f46cf523f6c9f635f7;
    decBuf[1128] = 256'h97f786f775f72cf7cef691f62ef6ebf5dff5bef5c8f5f6f50ff616f61df6e5f5;
    decBuf[1129] = 256'h92f52ff59cf4ecf345f3aef2fdf1b6f175f13af105f1d4f0a8f080f05bf03af0;
    decBuf[1130] = 256'h58f061f08bf0bff0c6f0b3f097f04af0fdefb7ef77ef3eef36ef14eff4eefaee;
    decBuf[1131] = 256'he0eed3eee8eee4eee0eef0eed0eea2ee76ee2deefbed16ee3feeb0ee83ef4cf0;
    decBuf[1132] = 256'h38f115f2def22df374f389f34ff3f5f2a4f278f26af246f23bf245f22af2f0f1;
    decBuf[1133] = 256'hbbf154f1edf0aaf055f0f2efafef2aefadee3beed4ed76ed52ed47ed79edefed;
    decBuf[1134] = 256'h61ee03efc6ef49f0bff02cf166f19cf1acf19ef190f16cf14bf141f15cf1a6f1;
    decBuf[1135] = 256'h14f2b7f24ef3fff3a5f43cf59ef5d4f5c4f5d3f5c5f5d1f5f2f54cf6b9f63ef7;
    decBuf[1136] = 256'hbbf74ef8d7f854f9a5f90dfa6afaa7fa0afb4dfba2fb05fc62fce8fc88fd20fe;
    decBuf[1137] = 256'hf8fe87ff3e008600c60001011301230132017501e2014902c20213033f034d03;
    decBuf[1138] = 256'h2803f102bf0292029a02ce023603ba035b041e05a0051706af06e9061f075007;
    decBuf[1139] = 256'h7c07bf07fc074908a308100977090a0abb0a610b240c0f0dad0d760ef90e6f0f;
    decBuf[1140] = 256'hb00feb0ffd0f2e105a108210bf100c115211b6112f1280120513821314149d14;
    decBuf[1141] = 256'h1a156c15b515de15b915981552150015c914ab147d1475148c14ae14f3145715;
    decBuf[1142] = 256'hb5152216a716dc164e177a176d1761174017fa16ba165f160a16a7154a15f514;
    decBuf[1143] = 256'ha814621422140914f313c313a313711333130a13e412c212e11214135113bd13;
    decBuf[1144] = 256'h24144c14701465141f14cd136a13f212c1129512a212c712e812de12c2127812;
    decBuf[1145] = 256'he2114b119a10f40f5c0fd30e320ec60d3d0d9c0c300c7f0b080b710a0f0a9209;
    decBuf[1146] = 256'h40091409ec08f8082f097509fe09870a280bc00b490c7f0cd00cc10c990c5c0c;
    decBuf[1147] = 256'h0f0cc90b9c0b620b3d0b360bfd0aba0a680ad9092809b108ef076c07f506b506;
    decBuf[1148] = 256'h7a0668067806870679066d064c06060690051e0599044004ef03e00308045d04;
    decBuf[1149] = 256'hc0041d0542054d0507057e04cd03c802d401f700f4ff45ff68fe9ffd1cfda5fc;
    decBuf[1150] = 256'h39fcd7fba2fb71fb62fb55fb49fb28fb0afbcafa90fa4cfa1ffa06fafff9f8f9;
    decBuf[1151] = 256'h0afa05fae1f9b7f963f90ef9c1f87bf84df856f85df880f8abf8bcf8b7f8a9f8;
    decBuf[1152] = 256'h7af84ff833f80ff801f805f8f9f7eff7ecf7c6f7a3f779f746f716f7eaf6adf6;
    decBuf[1153] = 256'h62f608f69bf516f599f428f4a3f36df33cf310f338f344f37bf3adf3c9f3e2f3;
    decBuf[1154] = 256'he9f3d4f3c2f3b1f3a1f3a6f3d5f30df460f4d9f44af594f5d7f5e3f5c2f590f5;
    decBuf[1155] = 256'h2cf5cef491f45af43cf446f46ff4a3f4fdf452f5cbf53cf686f6e4f639f75af7;
    decBuf[1156] = 256'h78f781f768f751f758f75ff786f7d3f720f87af8e7f813f93bf960f955f937f9;
    decBuf[1157] = 256'h2ef925f92df94ff955f945f92bf9e6f850f8b8f708f761f6f5f593f581f591f5;
    decBuf[1158] = 256'hbef5e6f53bf65cf68ef6a9f6b1f6b9f6cdf6e0f6f1f61ff74bf77ef7d7f714f8;
    decBuf[1159] = 256'h61f8a7f8d4f8edf8f4f8e0f8b4f898f86af857f873f897f8d3f82ef96bf9a2f9;
    decBuf[1160] = 256'hc0f992f958f906f98df81bf8d1f774f737f700f7cef68ef654f602f6b5f55bf5;
    decBuf[1161] = 256'heef486f444f4eff3cef3ecf3f5f31ef453f467f461f445f4f8f3abf379f339f3;
    decBuf[1162] = 256'h41f376f3c1f32ff4b4f40ef57ff58ef581f544f5f7f49df448f411f407f435f4;
    decBuf[1163] = 256'ha0f425f5c6f532f6bbf615f766f775f782f78ef76df777f792f79bf7c0f7f0f7;
    decBuf[1164] = 256'h29f86cf8acf8d5f80af92cf932f943f934f926f933f937f956f996f9faf958fa;
    decBuf[1165] = 256'hf5fa62fbebfb68fcb9fc03fd61fd85fdbcfd02fe30fe69febcfef3fe61ffe6ff;
    decBuf[1166] = 256'h6300f500cd019602b603c204b60594065d07e00756089708ab08e00832097b09;
    decBuf[1167] = 256'hf409a70a4d0b0f0cfb0c990d9b0e4a0fe80feb109911761240132b140815d115;
    decBuf[1168] = 256'h8816ff16961720187918eb1835195d199919a4199a199119891964196a197119;
    decBuf[1169] = 256'h7619c319261a841a091baa1b161ca01cf91c4a1d941df21d161e791ef11e431f;
    decBuf[1170] = 256'he51f5120b3203021612170217d2171213a2130211521eb20f320fa20e7200e21;
    decBuf[1171] = 256'h28213621652177217221772156211721c5206220ce1f6c1f131fa11e3a1edc1d;
    decBuf[1172] = 256'h571dfe1c6b1ce21b411baa1ad219091952184c179e168115c214cd132f136612;
    decBuf[1173] = 256'he3116d110111c6106c10fb0fb10f530fce0e510ebe0d350db80c460c1a0c0d0c;
    decBuf[1174] = 256'h190c3a0c800c9b0cb40cac0c7c0c1e0c8b0bdb0a050a3c095108b207e9066706;
    decBuf[1175] = 256'hc0055405f2045104e50334035f02cf01180172000600a4ff4aff19ffedfee0fe;
    decBuf[1176] = 256'hbbfe9afe7cfe4ffef4fd87fd20fd72fcccfb34fb84faddf946f995f81ff887f7;
    decBuf[1177] = 256'h25f7a8f636f6cff571f535f5fef4ccf4c3f4baf4d1f4f3f406f52df551f57bf5;
    decBuf[1178] = 256'hb9f5f2f545f6a8f6ebf640f777f781f753f72af7b9f627f69ef5fdf465f403f4;
    decBuf[1179] = 256'haaf359f32cf31ff3e2f2c1f253f2cff152f19ff0f9ef8cef03efcdeedeeeecee;
    decBuf[1180] = 256'hfaee36ef2bef21ef06efabee56ee09eeafed5bed24ed06edeaece2ecdaece1ec;
    decBuf[1181] = 256'hf4eceeece9eceeecd9eccdeccaecbaecb1ecc9ecd9ecfeec4bed82eddced31ee;
    decBuf[1182] = 256'h7eeeb0ee02ef23ef55efa7efdeef38f0a5f0eff032f156f14bf105f1c5f05af0;
    decBuf[1183] = 256'h10f0e8efc4efcfef01f01cf035f04bf01bf0e3ef9fef29efd8eeabee83ee8fee;
    decBuf[1184] = 256'hdcee22ef87ef1af07cf0d5f027f153f17bf19ff1c0f1def10cf235f25bf2a6f2;
    decBuf[1185] = 256'hd8f218f362f394f3e7f334f466f4a5f4dff405f519f539f533f52ef53cf526f5;
    decBuf[1186] = 256'h1bf525f51cf530f557f58af5d6f544f68df6ebf658f767f78ff783f74cf706f7;
    decBuf[1187] = 256'hc6f67cf64af62ef626f63df66df699f6b5f6cef6aef677f633f6bdf54bf501f5;
    decBuf[1188] = 256'ha3f47ff474f47ef487f4b0f4a9f4a2f476f422f4b5f34ef3d5f263f237f20ff2;
    decBuf[1189] = 256'h1bf252f25cf278f290f27af265f246f21ff205f21cf231f264f2aff2e1f20ff3;
    decBuf[1190] = 256'h38f331f30ef3eff2a6f274f246f20df2f6f1e1f1c2f1b1f1a2f178f146f116f1;
    decBuf[1191] = 256'hd1f091f057f014f0e6efbdef97ef90ef97ef91ef96efa4efa0ef9cef91ef82ef;
    decBuf[1192] = 256'h7fef97efbfef14f099f016f1c9f16ff2dbf23df373f383f392f385f391f3def3;
    decBuf[1193] = 256'h38f4bdf45ef521f6a3f649f7e1f743f89cf8eef81af95df9b2f915fa8dfafffa;
    decBuf[1194] = 256'h83fb24fc90fc1afdbbfd52fe03ffa9ff970074013d02f402ca0393044a05f005;
    decBuf[1195] = 256'hb3066a0740080909c009660afd0a870b280cbf0c480dc60d580eba0e370f880f;
    decBuf[1196] = 256'hd20ffa0f371058109e100211951146121c13e513d014ad1577162e17d4176b18;
    decBuf[1197] = 256'hf518b919701a461b491cf71c141ed31e821f2020e9203821ae211a227d22d622;
    decBuf[1198] = 256'h27235323b123ee23f9233f247f24b8240b256e25962503266a269226cf260627;
    decBuf[1199] = 256'h10272b2734270e270727dc2687264b26fe257c25fe248d24ea235323ca222922;
    decBuf[1200] = 256'h912108214320c11f1b1f581ea11d2a1d681ce51b3f1ba71a1e1a7d19bb186c18;
    decBuf[1201] = 256'hf5175e174a171517e416f316cb1676163f16bd151c158514fb133713b4123d12;
    decBuf[1202] = 256'hd1116f111611a4103d10a90ff90e530e900da50c070c3d0b870ae00949099808;
    decBuf[1203] = 256'h2208b5072c07af063d06b8053b05a90420047f03e70237029101ce004b00a5ff;
    decBuf[1204] = 256'h0effacfe76fe25fef8fd06fee1fdd6fdccfd9ffd76fd5ffd2ffd03fdfefce4fc;
    decBuf[1205] = 256'hdffcecfcf0fc01fd24fd3bfd50fd64fd59fd3dfd12fdbefc69fc06fc8efb1cfb;
    decBuf[1206] = 256'hd2fa75fa38fa17fa0dfa16fa2ffa45fa68fa87fa8dfaa6faabfa9efa9afa97fa;
    decBuf[1207] = 256'h8dfa90fa93fa9afaa9fab7fabcfac7fac6fab7faa1fa7bfa43fa00fac0f975f9;
    decBuf[1208] = 256'h43f904f9ebf8e3f8eaf809f93cf97af9b4f9f7f925fa3efa54fa4dfa3afa2afa;
    decBuf[1209] = 256'h10fa02fa06fa1afa32fa61fa91fab0fae3faf8fafefa04fbf4fad4faaefa7ffa;
    decBuf[1210] = 256'h47fa22fafff9f9f90afa19fa30fa46fa3afa14fad1f95af9e9f864f8e7f795f7;
    decBuf[1211] = 256'h69f741f74df758f762f76bf763f73ef71bf7fcf6d5f6bbf6c0f6bbf6c7f6dff6;
    decBuf[1212] = 256'hfcf626f759f77bf79af7cdf7eff71bf84ef870f883f89ff890f882f875f862f8;
    decBuf[1213] = 256'h50f853f85cf86ef892f8acf8c3f8d8f8dcf8d1f8cef8aff888f864f832f801f8;
    decBuf[1214] = 256'he2f7c6f7b7f7c5f7d1f7ddf7fcf7f8f7edf7dbf7acf77cf750f71ef7fbf6f5f6;
    decBuf[1215] = 256'hfbf6f6f616f71af716f71af710f7fcf609f71af736f770f7cbf707f854f886f8;
    decBuf[1216] = 256'hb4f8cdf8d4f8cdf8ecf809f937f994f9f2f95ffae4fa3dfb8ffbf6fb03fc0ffc;
    decBuf[1217] = 256'h1afce8fbbbfba2fb6dfb4bfb51fb40fb27fb35fb1ffbf5fad9fa96fa44faf7f9;
    decBuf[1218] = 256'h9df930f904f9a6f869f85ef82cf811f8f8f7b5f787f75ef71af7fff6f7f6eff6;
    decBuf[1219] = 256'hf6f615f71bf716f708f7c8f688f63ef6d0f5a4f57cf557f578f5d2f50ff672f6;
    decBuf[1220] = 256'hd0f6f4f615f71ff7dff6b6f672f60ef6e6f5c1f5b6f5c0f500f62af67cf6c9f6;
    decBuf[1221] = 256'h0ff761f782f7a0f797f77ef74af735f716f710f753f7b7f74af822f9ecf9d7fa;
    decBuf[1222] = 256'hb4fb44fcc6fc0efd4ffd89fd9bfdedfd54feccfe7fff55001e01d501da028803;
    decBuf[1223] = 256'h2704f0047205e9058106e3063c07ce075808b10864090a0acd0ab80b950c5e0d;
    decBuf[1224] = 256'h4a0e270fb70f6e10e4102511af1108125912c0123913ab134d140f1592156816;
    decBuf[1225] = 256'h3117b4175a18f1185319ad19fe192a1a6d1a921ac91a231b771bda1b6e1cf71c;
    decBuf[1226] = 256'h501de31d1d1e531e631e721e4a1e561e4b1e411e811e9a1ece1e1a1f381f531f;
    decBuf[1227] = 256'h6c1f551f331f141fcb1e851e571e0d1edb1dad1d631d1d1ddd1c721ced1b941b;
    decBuf[1228] = 256'h011b781a1f1a8c192a19ad183b18b7173a176616d71520151a146c138f12c511;
    decBuf[1229] = 256'hda103c10ac0ff60e7f0ebc0d3a0d930ca50b070b3e0a53097608e6072f078906;
    decBuf[1230] = 256'h1d066c05c6042e047e03d70240028f01e90052007affeafe68fec1fd2afdc8fc;
    decBuf[1231] = 256'h27fcbbfb59fbb8fa4cfac2f921f98af801f860f7c8f666f6e9f598f54ef5d6f4;
    decBuf[1232] = 256'h85f43bf4c2f351f307f3a9f285f264f246f261f26af262f25bf23cf2fef1c4f1;
    decBuf[1233] = 256'h81f12ff10ef1f0f0d4f0ccf0d4f0cdf0d3f0c2f0b3f0aef099f07ef06cf050f0;
    decBuf[1234] = 256'h3df032f01cf019f02cf038f04ff07ef0a0f0ccf0f3f0f9f0f4f0f8f0edf0e9f0;
    decBuf[1235] = 256'h05f120f155f1a7f1def124f276f2adf2b7f2d3f2dbf2e3f2f7f20af331f35ff3;
    decBuf[1236] = 256'h7ff3b1f3d4f3cdf3b1f398f352f30cf3dff2a5f27ff286f28df29df2b7f2bcf2;
    decBuf[1237] = 256'ha6f2a3f26ef23af217f2dff1b9f1b3f193f182f192f17bf165f15af133f105f1;
    decBuf[1238] = 256'hf2f0b5f07bf055f017f0cdef87ef35efe8eea2ee62ee28ee03eed3edb4eda3ed;
    decBuf[1239] = 256'h75ed3ced17edcbec85ec58ec1eecf8ebffebf9ebffeb2dec3fec50ec74ec70ec;
    decBuf[1240] = 256'h74ec78ec6dec64ec67ec5aec57ec6aec6dec8cecccecf9ec43ed9deddaed11ee;
    decBuf[1241] = 256'h43ee4cee54ee5cee47ee4eee6aee83eebfee1aef6fefd2ef30f06cf0b9f0ebf0;
    decBuf[1242] = 256'hf4f01ef143f166f19ef1f0f13df297f2ecf239f37ff3d1f31ef464f4c9f40cf5;
    decBuf[1243] = 256'h60f5adf5b7f5d3f5cbf5a5f590f597f59cf5caf51cf669f6aff613f73bf760f7;
    decBuf[1244] = 256'h81f777f780f777f77ff794f7bff7f2f730f87af8acf8ecf826f94bf96ef999f9;
    decBuf[1245] = 256'hb5f9e4f90ffa37fa65fa91fac3faf3fa38fb66fb8ffbc3fbe6fb12fc2efc29fc;
    decBuf[1246] = 256'h24fc20fc05fcecfbd0fbadfb8dfb80fb74fb71fb80fb95fbacfbc8fbd4fbd7fb;
    decBuf[1247] = 256'hd4fbc0fbaefb98fb84fb82fb8efba5fbcefbf5fb0ffc1cfc18fcf5fbccfb8efb;
    decBuf[1248] = 256'h44fb12fbd2fab9faa2fa8efa88fa82fa73fa6efa7bfa86fa98fac7faf7fa2ffb;
    decBuf[1249] = 256'h82fbcffb29fc96fcfdfc75fd08fe6afe0bff77ff00005900cb0032019001fd01;
    decBuf[1250] = 256'h8202ff02b2032904c0047105e70528068a06e40635079c07fa077f084409c609;
    decBuf[1251] = 256'h9c0a2c0be30b5a0cc60c280da50d170e7e0e110fc20f3810fb10b2112912eb12;
    decBuf[1252] = 256'ha213481436151416dd16c817a5183519ec19631afa1a841b241ce71c9e1da31e;
    decBuf[1253] = 256'h521f2f20f8207b2121228d22c8224523d7233a24da247225d4257526b626f126;
    decBuf[1254] = 256'h4a279b27c7274028b228fb288e29f129262a572a662a232a2f2a0e2af0291e2a;
    decBuf[1255] = 256'h572a7d2ac82afa2adf2ae72aa42a2d2adc297529fc28ab2861280428df279227;
    decBuf[1256] = 256'h1027b7264526a3253725ad240d247523ec2227227021ca200720511faa1ee81d;
    decBuf[1257] = 256'h651dbf1c271c9e1bd91a231a7c198e18b117e81631162c157d14a013d7122012;
    decBuf[1258] = 256'h1b1126100a0ffd0d090dec0be00a310a540951085d0780067d0589046c036002;
    decBuf[1259] = 256'h6c018e00c5ff0eff38fe6ffdb8fce2fb19fb62faecf929f9a6f830f8c3f73af7;
    decBuf[1260] = 256'he1f62ef6b7f520f56ff4c9f35df3fbf2c5f2b5f289f27bf26ff24ef208f2b6f1;
    decBuf[1261] = 256'h53f110f1a3f077f069f05df07ef0c4f004f13ef181f19df194f18df16bf14bf1;
    decBuf[1262] = 256'h2ff10bf1fdf002f1fef00ff132f149f167f191f1adf1c7f1f1f101f225f23cf2;
    decBuf[1263] = 256'h49f25df275f278f292f2c0f2dff228f382f3d7f324f492f4dcf41ef55bf57cf5;
    decBuf[1264] = 256'haef500f637f691f6fef648f7c0f732f87cf8f4f866f9b0f9f3f948fa69fa87fa;
    decBuf[1265] = 256'ha2fa89fa73fa5efa32fa21fa27fa2bfa49fa7bfa90faaffaaafa86fa53fa07fa;
    decBuf[1266] = 256'hadf958f90bf9d9f8acf8a3f89cf895f88ff867f839f801f8bef76bf734f7daf6;
    decBuf[1267] = 256'h9ef667f621f6cff598f552f524f5fbf4e4f4ddf4f0f401f510f515f5f7f4c5f4;
    decBuf[1268] = 256'h87f42cf4d7f3a0f36ef365f39ff3d4f311f44bf462f45bf42ff4dbf36ef324f3;
    decBuf[1269] = 256'habf25af22ef206f2e1f1d6f1b8f19df184f15ff13cf136f11af100f1f3f0c4f0;
    decBuf[1270] = 256'h8cf057f0feefc1efa0ef96ef9fefd9effeef3cf076f07ef077f064f031f01df0;
    decBuf[1271] = 256'h16f01cf040f07cf0b6f0eaf01af12df13ef158f15cf17af1b4f1ddf112f250f2;
    decBuf[1272] = 256'h69f27ff294f281f287f2aaf2c2f201f366f3c3f318f47bf4bef4e2f4edf4f7f4;
    decBuf[1273] = 256'h01f519f530f552f58af5b0f5d2f5f2f5f7f5f2f500f604f618f63ef658f66ff6;
    decBuf[1274] = 256'h8df689f68cf696f698f6b5f6eff64af7b7f73cf895f8e7f830f93ef94af929f9;
    decBuf[1275] = 256'hf7f8dcf8d3f8dbf8fdf835f96af9a8f9e2f907fa1cfa2efa29fa24fa28fa24fa;
    decBuf[1276] = 256'h28fa40fa5dfa8ffabffaf7fa3bfb7bfbb4fbf8fb26fc3efc46fc3ffc2cfc10fc;
    decBuf[1277] = 256'he2fbb6fb78fb4ffb2afb15fb1bfb37fb65fb9efbe1fb21fc4afc70fc84fc8bfc;
    decBuf[1278] = 256'h9cfcbffce9fc3dfddbfd9efe55ff5a000801e601af02fd027403e0031b049804;
    decBuf[1279] = 256'h0a058f0553060a07e007a9089409720a3b0bf20b980c2f0db90d5a0ef10e7a0f;
    decBuf[1280] = 256'h1b10b3108a111a120513a3136d14ef1496152d168f1630177117fa177718e918;
    decBuf[1281] = 256'h6e19eb195d1ac41a221b5e1bab1b191c631cdb1c6e1dd01d4d1e9e1eca1ef21e;
    decBuf[1282] = 256'hff1ef41efe1e2b1f541fc51f5720e120812119227b22d422e522f3220123f522;
    decBuf[1283] = 256'h00231e234b23642398239f2374234c23ff22862215229021ef208320d21f2c1f;
    decBuf[1284] = 256'h951ee41d3e1da61cf61b4f1bb81a071a321968187d176116541560148313b912;
    decBuf[1285] = 256'h02125c11f0103f10990fd70eeb0d0e0d450c250b190a6a098d08fd074607d006;
    decBuf[1286] = 256'h3806af050e054b049503bf02f6010a012d002aff36fe59fd90fcd9fb32fb70fa;
    decBuf[1287] = 256'hedf947f984f8cdf7f8f62ef678f572f4c4f3e7f21df29bf124f1b8f056f0fcef;
    decBuf[1288] = 256'habef44efe6ee91ee44eeeaed95ed48ed02ed9eec5beceeeba4eb61eb0debd6ea;
    decBuf[1289] = 256'hb8ea9ceaa4eabbeac2eae1eafdea0deb11eb0debeaeacaeaacea89ea84eaabea;
    decBuf[1290] = 256'hd9ea2aeba3eb15ec7cecdaec16ed63ed81ed9dedb5edf9ed39eeb5ee55efedef;
    decBuf[1291] = 256'h9df044f1dbf18cf232f39ef300f47df4cff418f576f59af5d1f517f633f65cf6;
    decBuf[1292] = 256'haef6e5f653f7d8f732f8a3f80bf94df95af97bf95df966f96ef984f9b5f906fa;
    decBuf[1293] = 256'h53fa99fad9fa02fb18fb1ffb0dfb07fb0cfbfefa0bfb1efb1bfb24fb2dfb20fb;
    decBuf[1294] = 256'h14fb12fbfcfae8fadafab7fa7efa59fa1bfae1f9bcf97ef955f93ef90ef9d6f8;
    decBuf[1295] = 256'ha1f848f8dbf774f7e0f67ef601f6b0f584f55cf537f516f5f8f4b8f45ef4f0f3;
    decBuf[1296] = 256'h89f311f3c0f258f215f2d9f1a2f15cf11cf1d2f078f03bf004f0e6efefefe7ef;
    decBuf[1297] = 256'hdfefe6efc7efa0ef7cef49ef19ef1fef30ef68efcaef42f0b4f01bf15ef19bf1;
    decBuf[1298] = 256'ha6f1b0f1a7f19ef197f1abf1cbf1f2f135f287f2d4f21af35af383f3a8f3cbf3;
    decBuf[1299] = 256'hc5f3caf3daf3e7f316f467f4b4f40ef57cf5c5f508f62df64ef658f661f669f6;
    decBuf[1300] = 256'h9df6e9f657f7dcf77df8e9f872f9ccf91dfa49fa71fa7dfab4fafafa4cfbaffb;
    decBuf[1301] = 256'h0dfc62fcc5fc08fd2cfd4dfd6bfd87fd9ffdb6fdcafdeafd06fe15fe23fe30fe;
    decBuf[1302] = 256'h43fe6afe98fec4fe0dff3fff7fff97ffaeffb5ffaeffa9ff99ff95ff99ffa5ff;
    decBuf[1303] = 256'hb6ffc6ffd4ffe7fff7ff060020003900550068007a0076006e00560040002c00;
    decBuf[1304] = 256'h1f00260039005600790090009d008a006a003300feffc0ff97ff90ff97ffb6ff;
    decBuf[1305] = 256'hddff01002100480061007800a700df0023017501d80136028b02d8021e037003;
    decBuf[1306] = 256'hbd0317049c043d05a9055a06d0063d079f07d407050831087408c9084209d409;
    decBuf[1307] = 256'h850a2b0bc30b250ca20cf30c3d0d9a0d200e790eeb0e700fc90f1a109f10d510;
    decBuf[1308] = 256'h6711f0116d122013f61386143d15e3154f168a16e316f3165b17b8173e180219;
    decBuf[1309] = 256'hed198c1a8e1b821ce11cab1df91d401eac1ee71e1d1f8f1f13206d201f219621;
    decBuf[1310] = 256'h0222b3222a239623f82375248524b224a42480245f2441240124092411241824;
    decBuf[1311] = 256'h5c248a24822489244b24e0237923e6223522be212721c5206b203b20d31fab1f;
    decBuf[1312] = 256'h561ff31eb11e431ea11d351dac1ce71b641b8f1aff194819a2183618d4175617;
    decBuf[1313] = 256'he5167d16ea15121549145e1341123511fb0fd40e140e660dc80cfe0b480b720a;
    decBuf[1314] = 256'ha90989083007eb05c404b8037e02ab01eb003d0060ffd0fe19fe43fd7afc8ffb;
    decBuf[1315] = 256'hb1fa22fa6bf995f805f84ef7a8f611f687f5e7f47af418f49bf329f3c2f24af2;
    decBuf[1316] = 256'hb8f12ef1b1f01ff095ef18efc7ee60ee02eec6ed79ed33ed05edcbec97ec67ec;
    decBuf[1317] = 256'h22ecd0eb83eb15ebadea50ea13eadce9e6e9efe908ea4cea79eab3ead8eadfea;
    decBuf[1318] = 256'hd9eadfeacfead4ea03eb2eeb83eb08ec85ecf7ec99ed05ee68eec1ee12ef3eef;
    decBuf[1319] = 256'h81efa6eff3ef39f079f0c3f031f198f110f282f2e9f262f3d4f300f443f47ff4;
    decBuf[1320] = 256'h8af4bcf4eaf403f546f586f5d0f516f668f69ff6e5f625f74ff774f7a4f7c3f7;
    decBuf[1321] = 256'hf6f726f852f890f8daf80cf95ef9c1f904fa59fabcfafffa3bfb72fb90fb9afb;
    decBuf[1322] = 256'hb2fbabfbb2fbc4fbbffbc4fbd2fbcefbd1fbd5fbccfbc3fbc0fbabfb97fb8afb;
    decBuf[1323] = 256'h66fb2efbf9faaefa54fa17facaf998f97df974f97cf990f997f986f962f91df9;
    decBuf[1324] = 256'h9bf81df8acf744f71cf710f71bf761f78ff7c9f7dff7d8f7b9f786f748f70ff7;
    decBuf[1325] = 256'he9f6c7f6c1f6ddf6ecf6faf618f71cf71ff722f71af712f70bf7f3f6ddf6c3f6;
    decBuf[1326] = 256'h9df66ff650f628f619f60bf607f60bf615f612f60ff607f6fbf5f1f5eff5e9f5;
    decBuf[1327] = 256'hf5f508f615f62bf64af657f67af69af6c1f6f9f62ef76bf795f7baf7cff7d5f7;
    decBuf[1328] = 256'hdbf7d6f7e3f701f834f87ff8c5f805f93ff946f932f9f9f8c5f887f85ef874f8;
    decBuf[1329] = 256'h97f8f4f852f9a7f9f4f926fa1dfa04fad0f99ff98df9a9f9ebf950fac8fa5afb;
    decBuf[1330] = 256'hbdfb16fc47fc73fc66fc59fc4efc58fc86fcc0fc12fd75fdeefd5ffea9feecfe;
    decBuf[1331] = 256'h29ff60ff7eff99ffb2ffd7ff15004f00a100ee00340162018b01a201a901af01;
    decBuf[1332] = 256'h9e01a301a801bd01e8010f023302530269026c02700273028d02c10214037703;
    decBuf[1333] = 256'hef036104e6043f0570059c05aa05ce0505067306da0688072e08c60828098109;
    decBuf[1334] = 256'hb209c109b309bf09e009120a770aef0a610bc80b0b0c2f0c240c1a0cff0be60b;
    decBuf[1335] = 256'hee0b1e0c560cb80c150d520d890da70d9e0da60d9f0d980db70df50d3f0ead0e;
    decBuf[1336] = 256'h320f8b0f1d108010d9102a117411b7110c128512f61299133014e11487151e16;
    decBuf[1337] = 256'h8016fe162e1720172d17391744177617c81715188318cd18f5180119ca185c18;
    decBuf[1338] = 256'hf5177d170b17fc1609172e177b17ad17b6179d174b17a616ff1568150615d014;
    decBuf[1339] = 256'hc014cf141215361541150f15ab1418146713c1125512f211e111d011fd11ef11;
    decBuf[1340] = 256'he311ac112a118910c70fdb0e3d0eae0d2b0de40ca30c410c0b0c990bf70a340a;
    decBuf[1341] = 256'h7e0978088407e6061d066605ef048304fa03a0030e035d02b701c900ecff5cff;
    decBuf[1342] = 256'ha5fe2ffec2fd88fd52fd01fd7cfcfffb6dfbbcfa16fa7ef9f5f8bff86ef842f8;
    decBuf[1343] = 256'h34f8f8f7abf729f788f6c5f50ef568f4d1f36ff339f329f31af30df3b8f255f2;
    decBuf[1344] = 256'hc2f111f16bf0a8ef26efdeeec9eeb5eeebee1bef2aef1defe0ee7dee05ee93ed;
    decBuf[1345] = 256'h0eedd9ecc8ecd7ec35ed8aededed4aee6fee64ee32eee0ed7ded3aed15ed20ed;
    decBuf[1346] = 256'h8eedf6ed89ee39efb0eff1ef05f0cfef9eef54ef2cef08ef29ef6fefc1ef24f0;
    decBuf[1347] = 256'h67f08bf080f04ef0fcefc5ef7fef64ef7defa2efe0ef3bf077f098f0b6f0adf0;
    decBuf[1348] = 256'ha5f0acf0c1f0f9f06af1fcf185f226f3bef320f49df4cef4faf422f546f593f5;
    decBuf[1349] = 256'hedf542f6bbf62df794f7d7f72cf84df87ff888f880f878f872f85ff84ef853f8;
    decBuf[1350] = 256'h4ef85bf87ef88cf8a1f8b5f8aaf894f886f85ef842f83df82ff83cf85ff876f8;
    decBuf[1351] = 256'h94f8aff8c0f8d0f8e4f8f7f811f945f96bf9a9f9e2f917fa2bfa4bfa3afa2afa;
    decBuf[1352] = 256'h1dfafff9ebf9e8f9e5f9e8f9f0f9e4f9d1f9b4f981f951f919f9d5f896f85cf8;
    decBuf[1353] = 256'hfaf79df730f7c8f66bf616f6dff5c1f5caf5c2f5baf598f553f501f59ef426f4;
    decBuf[1354] = 256'hb4f36af35df381f3cef328f495f41af573f5a4f5b3f5a5f599f58ef584f58df5;
    decBuf[1355] = 256'hc7f50bf65df6d6f627f78ef7d1f70ef819f837f81bf813f81bf814f81af836f8;
    decBuf[1356] = 256'h50f879f8a1f8baf8dbf8f0f803f915f931f94cf973f9a1f9c0f9f3f907fa1afa;
    decBuf[1357] = 256'h20fa1bfa16fa2bfa46fa7bfacdfa30fb8efbfbfb62fca5fccafcd5fcdffce8fc;
    decBuf[1358] = 256'hf0fc15fd53fdaefd1bfe82fefbfe4cffb3ffdbffe8ff0900130040007a00ae00;
    decBuf[1359] = 256'h08015d01aa01f0011d0247025d028d02ac02f6025003a40307048004d1041b05;
    decBuf[1360] = 256'h430567058805ce050e06690607079e074f08f508b7093a0ab10af20a540b890b;
    decBuf[1361] = 256'h9a0be30b410cae0c330dd40d400ec90e460f980fa60fb40f8f0f840f660f4b0f;
    decBuf[1362] = 256'h640f980fc80f26109f10cf1037115f11531148112a11fc10f4100a111f117011;
    decBuf[1363] = 256'hd3114b12bd1242139b13ed13191441147e149f14d11423158615c9154e16a716;
    decBuf[1364] = 256'hf9166017a317c717fe1730184b188518ba18c118ec18f218ce18c01891184018;
    decBuf[1365] = 256'h0918d71797177f176817381725170917c61699165f160d16d615a41576158f15;
    decBuf[1366] = 256'ha515ba15ff153e166816ab16d916e116f816f116d116cc16bc16a516bb16d616;
    decBuf[1367] = 256'he716161738173f1744171617b8165b16d5155815e71462140814d813ab136913;
    decBuf[1368] = 256'h44130d139f1238128a11b4102510390f5c0ecc0d150d9f0c5e0c230ced0bbd0b;
    decBuf[1369] = 256'h900b330bc60a410aa00909097f08de079d073b070607160707072f0754074907;
    decBuf[1370] = 256'h3f073607eb06910624069f052205b1042c04d20381033703f502d00299025302;
    decBuf[1371] = 256'hef015c01ab00d5ff0cff21fe44fdb4fcfdfb86fb45fb0afbf9fac8fa7efa3bfa;
    decBuf[1372] = 256'hcef967f9eef85cf8faf77df72cf7e2f69ff67bf670f666f65df665f66cf673f6;
    decBuf[1373] = 256'h86f675f647f61bf6d2f58cf54cf502f5e4f4dbf4e3f409f539f558f55ef56df5;
    decBuf[1374] = 256'h56f527f508f5caf490f46bf448f429f40df4f3f3dcf3d8f3ccf3d0f3ecf3fff3;
    decBuf[1375] = 256'h18f43af448f444f438f412f4e4f3d1f3c0f3c5f30af450f4c7f439f5a0f5fef5;
    decBuf[1376] = 256'h53f674f67ef699f680f688f68ff688f6a4f6bef6def6fcf627f743f767f790f7;
    decBuf[1377] = 256'h96f79bf797f779f746f716f7c5f68ef670f667f680f6b4f600f75af7aff7e6f7;
    decBuf[1378] = 256'h18f821f819f811f818f812f823f851f889f8dbf828f96ef9aef9f9f917fa44fa;
    decBuf[1379] = 256'h6dfa93faa8fac7fac1fabcfab7fa9afa77fa69fa5cfa58fa6afa6dfa70fa6dfa;
    decBuf[1380] = 256'h4afa07fac7f95cf9f5f897f82af8e0f7b8f794f75df73ff711f7d7f6a3f665f6;
    decBuf[1381] = 256'h2bf615f600f6faf50bf605f60af617f613f616f626f629f636f650f654f65df6;
    decBuf[1382] = 256'h66f659f651f654f64ef656f66ff680f696f6b0f6acf697f66bf627f6e7f59df5;
    decBuf[1383] = 256'h6bf54ff557f56ef59ef5d6f5edf501f6eff5bcf57ef534f5daf49df47cf472f4;
    decBuf[1384] = 256'h8ef4c7f40bf56ff5cdf522f685f6c8f6ecf623f741f74af763f788f7b9f70af8;
    decBuf[1385] = 256'h83f8f5f879f91afa86fa10fb69fb9afba9fbb6fbaafbb5fbbffbc8fbe1fb15fc;
    decBuf[1386] = 256'h45fc7efcb2fce2fc0efd35fd59fd83fdaafdcefde5fdfafdfefd02fefffd07fe;
    decBuf[1387] = 256'h29fe5cfea8fe16ff7dfff6ff6700cf002c0169018a01a801c301ec0112025e02;
    decBuf[1388] = 256'hb80225038c03ea035704a004e30438056f05a105e1051b06400670069c06b806;
    decBuf[1389] = 256'hd206e906070731076407a207ec0746089b08e8082e095c0974096d0958092d09;
    decBuf[1390] = 256'hfa08ca08ab08a508b408f0083b098109e509280a340a3f0a0d0abb096e091409;
    decBuf[1391] = 256'hbf089e08a808d60830098509e8092b0a500a450a270ae7098c094f090209d008;
    decBuf[1392] = 256'hb508ad08a5089e08a508940899088b087e088a0886087d0886087e0868085a08;
    decBuf[1393] = 256'h3d081a08160811081d084a088308c608060950096e099c0994098c0978096509;
    decBuf[1394] = 256'h3d0938092a0926093a094b095b0975098d09900993098609670949091709d908;
    decBuf[1395] = 256'hb0086c083f080508df07af0784075c0738070f07e706b9068d065b062b06ff05;
    decBuf[1396] = 256'hcc058e0555051105bf04880456042804100408040f042204270422041e04f703;
    decBuf[1397] = 256'hc90385034503fa02b40275023b0224020202fc01eb01d101b10182013d01eb00;
    decBuf[1398] = 256'h720000007cffdbfe43febafd61fdeffc88fc45fcf0fbcffb89fb49fbeefa99fa;
    decBuf[1399] = 256'h0afaa8f907f99bf839f8e0f78ff762f755f761f76cf776f77ff777f760f723f7;
    decBuf[1400] = 256'he9f696f633f6d6f581f534f516f5faf4f2f4faf40ef515f51af50bf5e1f4baf4;
    decBuf[1401] = 256'h6df420f4eef39cf365f347f32bf323f33af333f346f356f351f356f363f34ff3;
    decBuf[1402] = 256'h3ef32ef303f3d7f2bbf297f280f27cf278f28af2b2f2cef2e8f212f32ef33df3;
    decBuf[1403] = 256'h5df362f36df37ff375f378f385f37ef389f3a3f3b4f3ddf31bf455f498f4eaf4;
    decBuf[1404] = 256'h21f53ff56df565f55df549f529f524f529f537f55df595f5caf508f652f684f6;
    decBuf[1405] = 256'hc4f6edf604f718f71ef702f7e9f6d2f6abf69cf6aaf6b7f6e1f62af770f7c2f7;
    decBuf[1406] = 256'h0ff841f86ff888f871f85df83df816f811f81ff83df877f8c1f807f959f9a6f9;
    decBuf[1407] = 256'hd8f906fa2ffa45fa4cfa46fa35fa1cfa04fadef9d9f9e7f9fcf936fa91fae6fa;
    decBuf[1408] = 256'h33fb8dfbcafbebfbe1fbc5fbacfb78fb56fb36fb3cfb4bfb75fbbefbf0fb30fc;
    decBuf[1409] = 256'h6afc80fc87fc81fc59fc2bfc00fccdfb9dfb7efb56fb47fb4bfb47fb5bfb6cfb;
    decBuf[1410] = 256'h6ffb6cfb64fb41fb1dfbfdfad6fabdfaaffaa2faa6faa2fa99fa90fa83fa73fa;
    decBuf[1411] = 256'h68fa72fa89fab1faeffa3afb80fbbffbe9fbf0fbf7fbe4fbdffbdafbf1fb28fc;
    decBuf[1412] = 256'h7afcddfc56fde8fd4afea4fed4fe01ff29ff35ff2aff20ff29ff31ff48ff5cff;
    decBuf[1413] = 256'h95ffc9ff15005b009b00c400f8000d010701eb00d1009e007c00690063007d00;
    decBuf[1414] = 256'hb000ee004801b601ff015d02b202e902070334033d03440359036c039e03dc03;
    decBuf[1415] = 256'h26049404fc04740506066806c20613073f0732073e07490753078107ba070d08;
    decBuf[1416] = 256'h7008cd0822099b09ed09360a790ace0a050b4b0b8b0bb40bda0b0a0c1d0c440c;
    decBuf[1417] = 256'h5e0c750c9b0cde0c0b0d660dbb0d080e760ec00ee80e0c0f2d0f230f1a0f220f;
    decBuf[1418] = 256'h0c0f200f4c0f730fc00f3910ab103011ad11de1145126d12611256123812f811;
    decBuf[1419] = 256'hf011e811e1111a126c12cf124813b91303144614831478146e144014f613d813;
    decBuf[1420] = 256'haa1381139713ba13d9132d149a14e4145d15ae15bd15ca158d152a15cd146014;
    decBuf[1421] = 256'hf813b513a9139e13f81335148214dc140015f514d71497142c14e21385133013;
    decBuf[1422] = 256'hf912db12c012e912ff1206133e1355135c13621351130f13cf1284121612cd11;
    decBuf[1423] = 256'h8a114d114211381154116c1183117c1169112b11d11094103110ee0fb10fa60f;
    decBuf[1424] = 256'h880f7f0f770f520f2f0fea0e980e350ed80d830d4c0d1a0dec0cd30c9f0c610c;
    decBuf[1425] = 256'h270cd50b720b140ba70a220ac9095709f008ad08700839081b0812080a081208;
    decBuf[1426] = 256'hef07b70773070f0797062506a0052305f204c604d304f8041905370552053905;
    decBuf[1427] = 256'h1405d6046b04e6036903f70272021902e801bc01af01a3019801a20186015d01;
    decBuf[1428] = 256'h1901a300110087ffc3fe0cfe65fdcefc6cfc36fc06fcd9fbccfba8fb71fb2bfb;
    decBuf[1429] = 256'hb4fa22fa98f9f7f88bf802f8a9f757f72bf71ef712f707f7fdf6f3f6ebf6e4f6;
    decBuf[1430] = 256'hcff6b0f688f665f628f6eff5baf58af552f52cf518f505f50bf505f513f520f5;
    decBuf[1431] = 256'h24f512f5f6f4bcf461f40df4aaf34cf3f7f2c0f2a2f2bdf2e7f20cf358f376f3;
    decBuf[1432] = 256'h7ff387f353f315f3dbf289f252f234f218f220f255f277f2a3f2e1f20af330f3;
    decBuf[1433] = 256'h60f366f377f391f38cf390f394f38af38df3acf3c2f3fcf356f4abf4f8f466f5;
    decBuf[1434] = 256'hb0f5d8f5fdf5f2f5d4f5a6f56cf556f54ff555f571f5b4f5e1f52cf672f69ff6;
    decBuf[1435] = 256'hc9f6dff6caf6b8f69cf66df64ef649f639f65af699f6d9f623f77df7a2f7c3f7;
    decBuf[1436] = 256'hcdf7b1f788f754f708f7d6f6cdf6c5f6dbf60bf72bf747f760f75cf757f74cf7;
    decBuf[1437] = 256'h2cf720f714f702f7f3f6f0f6def6d2f6d4f6cef6d7f6eff607f72af74af757f7;
    decBuf[1438] = 256'h4bf73af70bf7dbf6a3f67df668f67bf697f6daf61af754f779f78ef76ef73cf7;
    decBuf[1439] = 256'h0cf7c7f699f691f699f6bbf6f3f637f777f7a0f7b6f7aff790f75ef720f7e6f6;
    decBuf[1440] = 256'hb1f68ff695f6a6f6caf606f72ff764f779f772f761f73ef701f7c8f6a2f68ef6;
    decBuf[1441] = 256'h94f6b0f6e8f62cf790f7d3f728f85ff87df886f88ef878f871f884f895f8b8f8;
    decBuf[1442] = 256'hfef858f9c5f92cfa8afadffa16fb48fb51fb49fb41fb3afb40fb51fb7ffbc4fb;
    decBuf[1443] = 256'h04fc5ffcb4fcebfc1dfd26fd2efd27fd20fd0dfd07fd17fd2efd54fd97fdd7fd;
    decBuf[1444] = 256'h21fe67fea7fee0fe06ff28ff54ff65ff7fffa8ffdbff19007300e1004801a501;
    decBuf[1445] = 256'hfa01470279029502ad02c402d902f8022a037603bc030e044504770493049b04;
    decBuf[1446] = 256'h840470045d04570467047e04a404c804df04f404f804ee04e404dc04cf04cc04;
    decBuf[1447] = 256'hd304d504e104ec04ee04f704fb0405051a05340553058205a105bd05cd05db05;
    decBuf[1448] = 256'hce05d205ce05d105f105170645067e06b206c706e606e006c706b00689065b06;
    decBuf[1449] = 256'h3c06200606060206fd05010605060e060506fe05e305b6057e053a05e8049b04;
    decBuf[1450] = 256'h69043b0444044b047b04b404d904ee04f404c10476041c04af0347030403e002;
    decBuf[1451] = 256'hd502070322035c038203890369033703eb0291023c02d9019601720167015d01;
    decBuf[1452] = 256'h66015e0165016c01590149011a01e2009f005f001500e3ffa3ff8aff73ff6dff;
    decBuf[1453] = 256'h66ff6cff67ff50ff32ff07ffd5fe97fe5dfe38fe15fe02fefdfdf8fdeafdddfd;
    decBuf[1454] = 256'hc2fd9bfd6dfd42fd0ffddffcb3fc97fc73fc65fc50fc35fc1cfcfafbc7fb97fb;
    decBuf[1455] = 256'h5ffb1bfbdbfa91fa4bfa1dfaf4f9def9e5f9f7f9fdf90cfa08faeaf9bff976f9;
    decBuf[1456] = 256'h1cf9e0f893f861f845f84df864f886f8b2f8cef8e8f8daf8b4f890f84af8f0f7;
    decBuf[1457] = 256'hb4f767f735f707f7fff606f71bf73af762f790f796f790f76df727f7cdf678f6;
    decBuf[1458] = 256'hfff5aef582f55af566f587f5a5f5d2f50cf605f6f0f5d1f588f542f502f5b8f4;
    decBuf[1459] = 256'h86f47cf464f47af49df4c8f4f0f428f54ef562f581f571f557f52df5fbf4cbf4;
    decBuf[1460] = 256'habf49af4a0f4c0f4def408f530f53ff531f51cf5e2f4a8f483f452f44cf45df4;
    decBuf[1461] = 256'h62f479f497f493f482f46cf441f421f41cf421f438f478f4a5f4dff405f519f5;
    decBuf[1462] = 256'h13f502f5def4d0f4d5f4e0f40ef546f58af5c9f503f629f64bf66af67bf69ff6;
    decBuf[1463] = 256'hc9f6e5f609f729f736f749f762f771f791f7c8f70cf84cf8a6f8e3f81af938f9;
    decBuf[1464] = 256'h41f928f912f9eff8e9f8faf814f947f992f9c4f904fa3efa72fa95fab4fabafa;
    decBuf[1465] = 256'hd3faeafaf7fa0afb23fb39fb5efb97fbdafb2cfc8ffcedfc42fd8ffdadfdb6fd;
    decBuf[1466] = 256'h9dfd69fd46fd40fd46fd7efdd0fd33feacfefdfe29ff51ff45ff24fff2fee9fe;
    decBuf[1467] = 256'he1fe06ff44ff8fffe9ff3d008a00bc00ea00030119012e014d0175019801c201;
    decBuf[1468] = 256'hf501250251028302b302f802380361038703a903af03aa03a503a003b503e003;
    decBuf[1469] = 256'h1e046804c2041705640582058b0572056b0556055c058405bc050f068806d906;
    decBuf[1470] = 256'h40078307c007e107ff070808310856087908be08fd0837098a09d7091d0a6f0a;
    decBuf[1471] = 256'hd20a150b6a0bb70be90b280c410c490c5d0c700c810caf0cf40c340d8e0de30d;
    decBuf[1472] = 256'h1a0e4c0e680e5f0e670e6e0e4f0e540e4f0e410e4e0e5a0e5d0e860ead0edb0e;
    decBuf[1473] = 256'h130f480f6a0f8a0f8f0f760f710f5c0f410f4b0f670f920fe60f3b107210b810;
    decBuf[1474] = 256'he610ee10f510ef10cf10ca10c510b710d410e010e410f310f610e910f510ff10;
    decBuf[1475] = 256'hfd1018111c1111110811e810b1108b105b103c1036103b1037105d1062105410;
    decBuf[1476] = 256'h50102d10fa0fd80fac0f850f800f7b0f6e0f7a0f6f0f4d0f3f0f2a0f070f0c0f;
    decBuf[1477] = 256'h180f1c0f3c0f490f450f410f2b0f000fe10ed00ec10ed80ee50ee80e010ff80e;
    decBuf[1478] = 256'hd20eae0e7b0e3e0e250e0e0efa0d000e060eec0dd50da60d550d1e0dd80caa0c;
    decBuf[1479] = 256'h910c8a0c830c890c8f0c800c720c540c220cff0bec0bd00bd50bd10bcd0be00b;
    decBuf[1480] = 256'hdc0bcd0bd00bd20bd50bf50b1e0c3a0c680c6f0c530c390cfd0bc30b9e0b890b;
    decBuf[1481] = 256'h8f0bb70bef0b140c370c3d0c0a0cda0b890b260bfe0ac10ab60aac0ac80abf0a;
    decBuf[1482] = 256'hc70aa50a790a460a080acf09b809b1099e09a40995096b093809fb08b0087e08;
    decBuf[1483] = 256'h510838083f0846084d08520843082208fc07c407800740070707d206b0067806;
    decBuf[1484] = 256'h43060506cb0588055a052105fb04d904a0046c042e04c3035c03e30271020a02;
    decBuf[1485] = 256'hc7018b016a014c0143013a012401f400c8008a0040000e00ceff84ff3efffefe;
    decBuf[1486] = 256'hb4fe5afe1dfed0fd9efd83fd6afd71fd5dfd3dfd00fda5fc1ffc7ffbe7fa37fa;
    decBuf[1487] = 256'hc0f954f919f907f917f908f9fbf8bef871f817f892f715f783f6f9f57cf52bf5;
    decBuf[1488] = 256'he1f49ef47af459f43bf444f43cf425f41ef4fff3d8f3b4f381f343f31af303f3;
    decBuf[1489] = 256'heff202f31ef342f37ef3a7f3dbf3fef304f4fef3f9f3e2f3bcf3a2f379f351f3;
    decBuf[1490] = 256'h2df30df3eff2ebf2e8f2ebf20bf317f31bf31ff3f6f2c4f293f242f20bf2edf1;
    decBuf[1491] = 256'hc0f1b7f1cef1e2f102f229f22ef23cf251f246f242f24cf249f251f26bf267f2;
    decBuf[1492] = 256'h71f27ff272f279f290f29af2bff2edf20cf334f358f35cf361f35df344f33bf3;
    decBuf[1493] = 256'h38f326f323f32ef324f322f324f313f30df317f319f327f345f352f365f370f3;
    decBuf[1494] = 256'h66f352f340f321f314f320f338f367f3cef336f4aef420f587f5caf507f63ef6;
    decBuf[1495] = 256'h5cf689f6b2f6e7f633f779f7cbf744f895f81af973f9c4f92cfa54fa60fa55fa;
    decBuf[1496] = 256'h37faf7f9cef9b7f995f99bf9b7f9d1f9faf917fa26fa18faf2f9aff96ff925f9;
    decBuf[1497] = 256'hdff8b1f8a9f8a2f8c4f8e3f80bf91af928f91bf908f9eff8d3f8c8f8c4f8c7f8;
    decBuf[1498] = 256'hdbf803f92af958f984f9b7f9e7f906fa22fa31fa36fa29fa1efa1afa1dfa37fa;
    decBuf[1499] = 256'h6cfaaffaeffa4afb86fba7fbb1fb96fb5cfb0afbbdfa8bfa82fa8afacdfa32fb;
    decBuf[1500] = 256'h8ffbfdfb64fca7fccbfcecfce2fcd9fce1fce9fc0bfd50fda2fd05fe7dfeeffe;
    decBuf[1501] = 256'h74ffcdff3f008900e6000b0116010c01f000c700b1008e0088009900b200e500;
    decBuf[1502] = 256'h23014c017201790166013301f6009b004600f9ffc7ffacffb4ffbbffdefffdff;
    decBuf[1503] = 256'h2400480072008e009d00ab00af00ac00a800a500a800bf00e2001e016801ae01;
    decBuf[1504] = 256'h00026302a602e3021a03380365037e0386039a03ad03a703a20394037f036403;
    decBuf[1505] = 256'h530349034c035e0374038e039f03960376033f03ec0289022c02d701a0018201;
    decBuf[1506] = 256'h8b01a401d80116023f02650287028e02880279026102440229020902f401e801;
    decBuf[1507] = 256'hec01fb0121024f027b02ad02d002d602c5028d023a02d70179010c01a5006200;
    decBuf[1508] = 256'h3e00490053005c0075008b00840072004a001200ceff8eff44ff12ffe5feccfe;
    decBuf[1509] = 256'hc4fee7fe12ff50ff8affceff0d0037003e004500320021001c00210036005900;
    decBuf[1510] = 256'h9500cf00210158018a01a601bf01d501ce01c801c201a9019201740149010b01;
    decBuf[1511] = 256'hd2008e003c000500bfff91ff58ff32fff4feaafe64fe12fec5fd7ffd2dfdf6fc;
    decBuf[1512] = 256'hb0fc82fc59fc24fc02fceffbeafbf9fb19fc40fc6efca6fccbfce0fce6fccafc;
    decBuf[1513] = 256'hb1fc90fc72fc67fc71fc9afcd8fc33fd87fdd4fd1afe36fe4ffe47fe32fe07fe;
    decBuf[1514] = 256'hdffdbbfd9bfd8efd92fda4fdc6fdf9fd29fe61fe87fe9bfe95fe6efe2bfed9fd;
    decBuf[1515] = 256'h8cfd46fd18fd10fd27fd57fd8ffdd3fd12fe2bfe33fe1efef2fdcbfda7fd87fd;
    decBuf[1516] = 256'h7afd7efd88fd98fdacfdaffdacfda2fd84fd66fd43fd10fde0fcb4fc76fc3dfc;
    decBuf[1517] = 256'h08fccafb91fb5cfb3afb0efbf2fac4fa98fa65fa35fafdf9d7f9c3f9bdf9c2f9;
    decBuf[1518] = 256'hdcf9fcf922fa32fa40fa44fa31fa2dfa2afa33fa4ffa7afab8fa02fb5cfbb1fb;
    decBuf[1519] = 256'hfefb44fc84fcbefcf2fc15fd34fd39fd3ffd3afd3efd42fd5bfd83fdc1fd0bfe;
    decBuf[1520] = 256'h65febafef1fefbfee0fea6fe36fec4fd5dfdfffcc2fccdfcebfc2bfd86fddbfd;
    decBuf[1521] = 256'h12fe44fe3bfe22fedefd8cfd3ffde5fcc1fca0fcbefcecfc36fd90fdfdfd47fe;
    decBuf[1522] = 256'ha4fee1feecfef6fedbfeb1fe8cfe5cfe49fe4ffe5efe7efeb6feeafe28ff51ff;
    decBuf[1523] = 256'h86ffa8ffc7ffcdffd2ffcdffc1ff9eff7dff4fff23ff12ff0dff24ff5bffaeff;
    decBuf[1524] = 256'h11006e00c300fa002c012301fa00d400a40085008b00af00f4006201e7016402;
    decBuf[1525] = 256'hd6023d039a03d703f80316041f0427042f0436043c044d0467048704a504d704;
    decBuf[1526] = 256'h0705330566058805a705ad059305730544050c05c8049b0461044a0444044a04;
    decBuf[1527] = 256'h7c04ba0405055f05b305000632064e06560640061d06fe05f805080631068606;
    decBuf[1528] = 256'h0b07ac074308f4086b09020a3d0a4f0a3f0a300aed09c909a8099e09b909030a;
    decBuf[1529] = 256'h710ad80a6c0bce0b270c370c290ce60b790bd60a6a0ae1098709570948097009;
    decBuf[1530] = 256'had09fa09180a330a2b0af609ab095109e4089a0857083308540872089f08d908;
    decBuf[1531] = 256'h1c093809510967096009730979097e099509aa09b609c009bd09a90997097809;
    decBuf[1532] = 256'h510942093409270933094c095b0975098709770963093b09f208ac086c082208;
    decBuf[1533] = 256'h0408e907f107170847087f08c208f008190921091a09ee08d2089a0865085108;
    decBuf[1534] = 256'h4a08450869089b08d90824096a09a909e309eb09e409c50987092c09d7087408;
    decBuf[1535] = 256'h1608f207d107c707e207eb0701080808e907ab075007cb064e06bb055905dc04;
    decBuf[1536] = 256'hab047f048d049904ba04c404df04e704d104ca04ab04830474045d0450046304;
    decBuf[1537] = 256'h75048504aa04c404d104e704f20404051a0528053a0550055805510549052e05;
    decBuf[1538] = 256'hfb04cb04870447040d04e703c503bf03c403ca03d703d303b8038b034603f402;
    decBuf[1539] = 256'h91023302de01a70175015a01520159017b019b01b701c601dd01d901d501bd01;
    decBuf[1540] = 256'ha1017e015d014001240121012401380160019201c201fb01110226021302ec01;
    decBuf[1541] = 256'h9f015201e4007c003a00e5ffc4ffbaffc3ffdcfff2ff07000000f0ffadff5bff;
    decBuf[1542] = 256'hf8fe9afe2dfee3fda0fd7cfd87fda5fdc0fdfafd2ffe51fe57fe52fe38fe0efe;
    decBuf[1543] = 256'hdcfdacfd80fd64fd54fd59fd66fd79fd8bfda1fda9fda7fd9bfd7ffd54fd22fd;
    decBuf[1544] = 256'hf2fcc6fc88fc5ffc39fc17fcf8fbdcfbb8fb97fb71fb43fb17fbe5fab4faa2fa;
    decBuf[1545] = 256'h86fa6cfa5efa51fa3efa25fa09fae6f9cff9baf9aef9b2f9cef9f1f92dfa77fa;
    decBuf[1546] = 256'hbdfafdfa37fb5cfb71fb84fb7efb6ffb6afb66fb6afb82fbb1fbeffb39fc7ffc;
    decBuf[1547] = 256'hbffcf9fc1efd33fd20fd04fdd6fc9efc69fc47fc34fc3afc53fc7dfcbbfcf5fc;
    decBuf[1548] = 256'h38fd54fd6cfd65fd42fd17fdcefc88fc48fc0efce8fbeffb02fc35fc80fcc6fc;
    decBuf[1549] = 256'h06fd2ffd37fd15fde9fc94fc40fcddfb9afb5dfb52fb5cfb8afbd4fb06fc46fc;
    decBuf[1550] = 256'h6ffc77fc54fc1cfcd8fb74fb31fbdcfabbfa9dfaa6fad0fa04fb50fb96fbd6fb;
    decBuf[1551] = 256'hfffb06fc0dfcfbfbdefbc5fbaefbb2fbc5fbe5fb1cfc60fc9ffcd9fc0efd30fd;
    decBuf[1552] = 256'h43fd54fd4ffd4afd46fd42fd3efd48fd45fd47fd4afd3ffd35fd33fd2bfd27fd;
    decBuf[1553] = 256'h30fd34fd3afd41fd35fd24fd09fdd5fca0fc70fc2cfcecfbc2fb9dfb96fb9cfb;
    decBuf[1554] = 256'ha2fbb1fbc8fbc4fbb9fb99fb62fb1efbdefa84fa47fa26fa08fa11fa2afa5efa;
    decBuf[1555] = 256'h81faadfac9facefac9faabfa81fa59fa36fa15fa08fa05fa16fa38fa62fa89fa;
    decBuf[1556] = 256'hc2faf6fa19fb44fb55fb65fb69fb5dfb49fb3ffb2ffb32fb44fb63fb9afbedfb;
    decBuf[1557] = 256'h3afc80fcd2fcf3fc11fd1afd01fddcfcbafc9afc89fc84fc92fcb8fcf1fc25fd;
    decBuf[1558] = 256'h55fd9afdb6fdcefdd6fdcffdbcfda0fd86fd66fd59fd4efd58fd68fd82fdaffd;
    decBuf[1559] = 256'hdbfd0efe4bfe75fe9afebdfec3fec8feb9fe99fe7bfe58fe41fe34fe38fe5ffe;
    decBuf[1560] = 256'h97fedafe3fff82ffbefff5ffebffd0ff86ff2cffd7fea0fe6efe77fea0fef3fe;
    decBuf[1561] = 256'h6cffddff4500a200df00ea00cc008c0052000000c9ffabffa2ffcbffffff5900;
    decBuf[1562] = 256'hc6002d018b01e001170221021802ee01ba0160012401ed00cf00c600ef003201;
    decBuf[1563] = 256'h8501e8012a026702720254021402b9014c01c8004a00f9ffafff87ff93ffb4ff;
    decBuf[1564] = 256'he6ff14003d0063005c003d00ffffb5ff5bffedfea4fe7cfe57fe62fe94fed4fe;
    decBuf[1565] = 256'h1eff78ffcdff0400360052005a0052003e001e00f7ffddffd0ffd4ffe7ff1500;
    decBuf[1566] = 256'h5900ac000f016c01c101f8010202e701ad015a01f700b5007800570061008f00;
    decBuf[1567] = 256'hc8000c01390163015b012b01e60082002400cfff98ff66ff5dff66ff7cff91ff;
    decBuf[1568] = 256'ha3ffb4ffafffabff95ff7aff69ff5fff57ff59ff5cff55ff4bff38ff1bfff1fe;
    decBuf[1569] = 256'hc9fe9bfe7cfe76fe7bfe92feb0fedbfef7fe11ff03ffe5feabfe61fe1bfedbfd;
    decBuf[1570] = 256'hb1fdaafdbffdeafd33fe79feccfe03ff35ff3eff35ff1fff0afff8fee7feecfe;
    decBuf[1571] = 256'hfafe0fff32ff5bff8effccff16005c009c00e600180134013c012501f500bd00;
    decBuf[1572] = 256'h7a003a00210019002e005a00a300e90017012f012801f8009a003c00b7ff3aff;
    decBuf[1573] = 256'he9fe81fe59fe4dfe58fe76fea4feddfe03ff18ff1eff0dffdffea7fe63fe23fe;
    decBuf[1574] = 256'he9fdb5fda0fda7fdcefdfcfd41fe93fee0fe12ff40ff58ff60ff4bff1fffedfe;
    decBuf[1575] = 256'haffe75fe50fe3bfe4efe75feb8fe0aff6dffcbff07003e0048002d00f3ffb0ff;
    decBuf[1576] = 256'h70ff36ff10ff0aff1cff4fff9bfff5ff49009600c800f600fe000601e300c400;
    decBuf[1577] = 256'h9200610036000e00f5fff9ff170049009500ef0044019101af01b8018f014b01;
    decBuf[1578] = 256'he7006f00fdff96ff53ff2eff39ff57ff97ffd1ff05001a001400ecffb4ff62ff;
    decBuf[1579] = 256'hfffea1fe4cfe15fe0bfe02fe1bfe4ffe7ffed1fe08ff4eff8dffa6ffbdffd1ff;
    decBuf[1580] = 256'hcbffbaffabff94ff87ff8bff8effa4ffcfff14006600c90027019401de012102;
    decBuf[1581] = 256'h450250023202e00193014d011f0106011d015b01c6012d02c00223037c038c03;
    decBuf[1582] = 256'h60031d0398021b028801ff00a60075008400ac0001014e01bc01050248025402;
    decBuf[1583] = 256'h3302ed01890111019f003800f5ffd0ffdbff21008600fe007001d7011a023e02;
    decBuf[1584] = 256'h1d02eb0199013601d9006b003f00170023005a00b4002101a60123027402be02;
    decBuf[1585] = 256'he602f202bb0275021102b3017701560160018d01e8016e02eb025c03c403ec03;
    decBuf[1586] = 256'hf803d70391032d03cf027a024302390242026b02af0201036403c20317044e04;
    decBuf[1587] = 256'h6c0475045c042704ea039f0359032c030203fb021d0349039203d80318044104;
    decBuf[1588] = 256'h49043404fc03b80354031103bc02850267025e0277029c02da0225036b039803;
    decBuf[1589] = 256'hb103c703b303940361032303e902c402af02a902c502f3021f03520374039303;
    decBuf[1590] = 256'ha403a9039b039703930390038d038f0388038a03880386039203a403be03ec03;
    decBuf[1591] = 256'h17043f046d0480048504760455042704fb03c80398038503800370037e038303;
    decBuf[1592] = 256'h8e039903a803b103b903c003be03b803a80388035f0337031303f302e602ea02;
    decBuf[1593] = 256'h0a03380364039703c703da03ea03d103a70369031f03d902990270024a024402;
    decBuf[1594] = 256'h4a0266029402cc02f2022203350324030a03ce0284023e02fe01c401ae01b501;
    decBuf[1595] = 256'hd40112024b028f02bd02e602ed02e602c702a00267022402e401bb0195018e01;
    decBuf[1596] = 256'h9501b101e9012d027f02b602fc020503fd02d7028c023202dd0190015e015501;
    decBuf[1597] = 256'h5d018201b201de0106020b02fd01d7019e015b011b01d1009f005f0046002000;
    decBuf[1598] = 256'h0c00f9ffffff180039005f009700cc00ee000d011301f900d900b30085005900;
    decBuf[1599] = 256'h48004d006e00a500e80028017201b801e601ee01d801b5017d012b01de009800;
    decBuf[1600] = 256'h6a00620069008c00c400f8002901480142011e01e20098003e00e9ff86ff5eff;
    decBuf[1601] = 256'h21ff00fff6feedfee5feddfed7fed0fed6fed1fed5fed1febefe97fe69fe24fe;
    decBuf[1602] = 256'he5fdabfd94fd8dfda0fdd3fd1efe78feb5feecfe0aff01ffc7fe93fe47fe01fe;
    decBuf[1603] = 256'hd3fdbbfdc2fde5fd1dfe60fea0fec9fefefe13ff19ff13fffafee2fecdfebafe;
    decBuf[1604] = 256'haffeacfebbfed2fef5fe1eff46ff69ff8affa8ffbbffbeffc2ffbfffb7ffabff;
    decBuf[1605] = 256'h98ff85ff75ff66ff60ff5eff6aff80ffa9ffd0fff4ff0b000f00fcffd5ff9dff;
    decBuf[1606] = 256'h5aff1affe0fec9feb5fec8fee4fe08ff1fff2bff28ff0fffe6feb4fe91fe72fe;
    decBuf[1607] = 256'h61fe5cfe6afe7ffe9afeacfebcfecafecdfed4fed6fed8fedafedbfeddfedefe;
    decBuf[1608] = 256'hdffee3fee4fee5fee9fef1fef4fef7fefafefbfefcfefefe01ff0eff24ff38ff;
    decBuf[1609] = 256'h55ff70ff7bff84ff81ff74ff68ff59ff4bff49ff4bff56ff62ff71ff77ff78ff;
    decBuf[1610] = 256'h7aff6fff66ff62ff5cff59ff59ff54ff53ff4fff47ff41ff42ff47ff50ff65ff;
    decBuf[1611] = 256'h79ff8cff97ff9eff94ff81ff64ff41ff17fff0feccfeacfe8efe7afe70fe60fe;
    decBuf[1612] = 256'h5dfe5bfe54fe52fe4cfe3ffe2afe0bfee4fdb6fd8afd63fd54fd58fd6efd90fd;
    decBuf[1613] = 256'hc3fde6fd05fe0bfe05fee5fdb6fd7efd59fd36fd23fd29fd38fd59fd7ffda3fd;
    decBuf[1614] = 256'hbafdc7fdd2fdcffdccfdcffdd7fddefdedfdfffd0ffe22fe35fe45fe58fe66fe;
    decBuf[1615] = 256'h71fe80fe8afe90fe98fe99fe98fe94fe8afe78fe63fe43fe1dfef9fdd9fdc3fd;
    decBuf[1616] = 256'hb8fdbbfdc5fddefdf7fd07fe15fe08fef2fdcdfd9ffd73fd57fd3dfd42fd57fd;
    decBuf[1617] = 256'h7afda4fdcbfde5fdf3fdf7fddcfdbcfd96fd72fd52fd45fd39fd44fd54fd68fd;
    decBuf[1618] = 256'h85fda0fdb8fdd4fdeffd01fe11fe19fe1cfe19fe1cfe1afe1bfe27fe34fe47fe;
    decBuf[1619] = 256'h5ffe6ffe77fe7ffe73fe5cfe46fe21fef3fdd3fda1fd7efd6cfd4ffd4afd46fd;
    decBuf[1620] = 256'h41fd4dfd58fd5bfd5efd5bfd4ffd3cfd2afd0ffdfefcf5fcf2fcfffc14fd28fd;
    decBuf[1621] = 256'h3bfd47fd3cfd26fd01fdd2fca7fc8bfc67fc62fc6ffc7afc9afcb8fccbfcddfc;
    decBuf[1622] = 256'he0fcddfcd0fcc9fcbefcc4fcd0fcdffcf9fc18fd2efd41fd52fd4ffd47fd34fd;
    decBuf[1623] = 256'h1afdfbfce5fccafcb2fca8fc94fc8cfc8afc84fc7afc7bfc77fc6ffc73fc77fc;
    decBuf[1624] = 256'h81fc93fca4fcb7fcc4fccbfcc5fcbffcabfc99fc8dfc82fc84fc94fca3fcb1fc;
    decBuf[1625] = 256'hc1fcbffcb5fc9afc68fc38fc0cfce5fbcbfbd0fbe5fb10fc42fc72fcabfcd0fc;
    decBuf[1626] = 256'he5fcdffccefcaafc89fc6cfc58fc55fc6bfc85fcabfcd9fc05fd21fd30fd35fd;
    decBuf[1627] = 256'h28fd15fdeefccbfcb3fc9efc9afcacfcc8fcebfc1efd40fd6cfd93fda3fda7fd;
    decBuf[1628] = 256'ha3fd9ffd95fd91fd89fd8bfd97fda2fdb4fdcefde0fdeffd03fe10fe1cfe27fe;
    decBuf[1629] = 256'h31fe3afe45fe4dfe53fe5cfe64fe73fe86fe99feb3fed2fef0fe13ff33ff51ff;
    decBuf[1630] = 256'h74ff82ff8eff9aff9eff8eff85ff7dff76ff70ff6eff70ff7bff89ff95ffa3ff;
    decBuf[1631] = 256'hadffb3ffaeffa3ff8fff75ff5cff40ff25ff1bff1eff2cff3eff5dff7bff96ff;
    decBuf[1632] = 256'hafffbeffc7ffc4ffb8ffaaffa0ff97ff98ffa3ffb5ffd4fffaff280047006f00;
    decBuf[1633] = 256'h9300a000ad00b100ae00a400a700aa00b100c800de0003012701480165018101;
    decBuf[1634] = 256'h8b018e018b017e01720163015d015c016101650171017d0184018b018f018e01;
    decBuf[1635] = 256'h8b0185017f017c017d017e018b019901a201b301bf01c601d001d101d001d401;
    decBuf[1636] = 256'hd301d401dc01e901f90110022602340247024e024802420235022a0228022f02;
    decBuf[1637] = 256'h3b02510273029402ba02d402e202e602e202d002c102ad02a0029d029f02ad02;
    decBuf[1638] = 256'hc102d802e802fc0209030b030903ff02ec02df02d302c802c602d302de02f502;
    decBuf[1639] = 256'h110324033d034c034f0357035503460340033a033203340338033c0344034703;
    decBuf[1640] = 256'h46034803470341034b035703660380039803ae03c203d503d703d503cf03c303;
    decBuf[1641] = 256'hbe03bf03c103d403eb0301042104360442044c04430429040904ec03c903b203;
    decBuf[1642] = 256'ha503a103b903d603f8032b044e046d047e0483046c04570434040a04f903e003;
    decBuf[1643] = 256'hdb03e803fb030d042f043d04410435042b040904e803c2039e03900383037803;
    decBuf[1644] = 256'h82039203a603c303e603fd031b04360439043c043a042c041c040d04ff03fa03;
    decBuf[1645] = 256'hfb0303041504250434043e04430438042e041e040804fa03ed03e103df03e903;
    decBuf[1646] = 256'hee03fa0304040804110419041604170416041104110411040a040404f903e503;
    decBuf[1647] = 256'hd803c303a3038e037b0362035f0368036a0380039403a103a803a60394038303;
    decBuf[1648] = 256'h68034d0342033f0342035f038203a203c003d303d703cd03b3038d0369034903;
    decBuf[1649] = 256'h2b031f031c032503330341033e033c032e031e030b03f902e802e602e802f102;
    decBuf[1650] = 256'hff0211031d032c032e032c0324031a030b03090307030c0319032d033f035003;
    decBuf[1651] = 256'h5a035403480330030903e502c502a70294029702ad02cd02f302210340035103;
    decBuf[1652] = 256'h4c033e032003f602ce02ab028a0286029202aa02c602e902090316031a030203;
    decBuf[1653] = 256'he502b30275023b021602e601e001e501f501150244026f028c029b02a0029302;
    decBuf[1654] = 256'h780251022d02160209020d0218022e024d0263026e0279026f0261024f023402;
    decBuf[1655] = 256'h1c020002ec01db01cb01c301b601b301b101b701b901c101cb01dd01e901f401;
    decBuf[1656] = 256'hf601f101df01c901af0197017b0167015d015a0157015a01650168016a016401;
    decBuf[1657] = 256'h590142012001f600da00b6009f009b009700a200ab00bf00cc00d300d100c700;
    decBuf[1658] = 256'hb4009700740054003f00240012000200f4ffecffe5ffd6ffccffc7ffbfffb4ff;
    decBuf[1659] = 256'hadffa5ff98ff86ff76ff63ff50ff44ff3eff40ff45ff54ff66ff77ff81ff87ff;
    decBuf[1660] = 256'h85ff81ff76ff67ff59ff4dff45ff40ff3fff3dff3fff40ff3fff3cff38ff32ff;
    decBuf[1661] = 256'h31ff2cff28ff25ff21ff17ff0eff00fff4fee8fedbfecffecdfecbfecafecbfe;
    decBuf[1662] = 256'hcffecefecbfec3feb7fea8fe96fe7cfe64fe54fe40fe38fe3afe3cfe42fe4ffe;
    decBuf[1663] = 256'h54fe58fe51fe41fe2efe16fe00feecfddffdddfde3fdedfdf2fdfafdfcfdf5fd;
    decBuf[1664] = 256'hecfddbfdc6fdb8fdb0fda9fdaffdb5fdbefdccfdcefdcdfdc5fdbafda8fd98fd;
    decBuf[1665] = 256'h89fd83fd88fd90fda1fdb4fdc1fdcdfdd7fdd1fdc2fdaefd97fd81fd73fd60fd;
    decBuf[1666] = 256'h59fd64fd6efd7dfd91fd9efda0fd9afd84fd6afd4afd24fd0afdf3fce7fce3fc;
    decBuf[1667] = 256'hedfcf7fc05fd12fd10fd05fdf7fcddfcc2fca2fc84fc71fc6efc64fc67fc6ffc;
    decBuf[1668] = 256'h71fc6ffc75fc70fc6bfc67fc5dfc54fc51fc4efc4bfc4cfc4dfc4efc50fc4afc;
    decBuf[1669] = 256'h46fc43fc3bfc34fc2ffc27fc21fc1efc1afc15fc18fc14fc0dfc0dfc03fcf9fb;
    decBuf[1670] = 256'hf3fbe9fbe2fbe6fbe7fbecfbf6fbfcfb03fc0bfc0afc03fc01fcf4fbeafbddfb;
    decBuf[1671] = 256'hcffbc5fbc3fbb8fbb0fbacfba6fba2fba5fba3fba2fba5fb9efb98fb92fb85fb;
    decBuf[1672] = 256'h77fb75fb6dfb69fb6afb70fb7dfb8ffb9afba5fbb3fbb1fbb0fba8fb99fb8bfb;
    decBuf[1673] = 256'h7ffb73fb6ffb70fb6ffb75fb80fb87fb94fba2fba4fba9fbb2fbb0fbaffbb0fb;
    decBuf[1674] = 256'hadfbaefbb2fbb5fbc0fbd2fbdefbf1fb03fc0ffc1afc1cfc1afc18fc14fc0afc;
    decBuf[1675] = 256'h01fcfefbf9fbf8fbfefb03fc0bfc1bfc27fc36fc48fc59fc63fc71fc7afc82fc;
    decBuf[1676] = 256'h8afc8bfc87fc8dfc90fc96fca3fcb1fcc1fcd8fceefcfdfc05fd02fd00fdf6fc;
    decBuf[1677] = 256'he3fccbfcbcfcadfca0fc9efca0fcaafcbdfcd5fcebfcfffc0cfd18fd1afd14fd;
    decBuf[1678] = 256'h04fdf5fce7fcdbfcddfce7fcf9fc1dfd40fd61fd87fda1fdaffdaafd9ffd8dfd;
    decBuf[1679] = 256'h77fd63fd5bfd59fd5ffd75fd95fdbbfddffd09fe25fe3efe56fe5afe56fe52fe;
    decBuf[1680] = 256'h49fe4cfe4ffe5afe72fe8efeb1fed1feeffe02ff0dff10ff07fffafeeefee4fe;
    decBuf[1681] = 256'hdafed8feddfeeafefafe09ff17ff23ff2fff39ff40ff4bff5cff6fff86ff96ff;
    decBuf[1682] = 256'haaffbdffc4ffc6ffc8ffc3ffbeffbcffbbffc1ffcbffd5ffdeffe5ffe8ffe8ff;
    decBuf[1683] = 256'he0ffd3ffc1ffb6ffabffa5ffa7ffafffc2ffdafff6ff19003000450059006300;
    decBuf[1684] = 256'h60005d005b0058005a006000700083009b00aa00b900c100c300c100b700b200;
    decBuf[1685] = 256'hb000b500c600dc00fb00190134015401690175017801750172017a017c017f01;
    decBuf[1686] = 256'h8d01a001b201c301cd01d301d201c301ad019901810165015a014f0152015b01;
    decBuf[1687] = 256'h72019501b501d301e601f801f501ec01df01ce01bf01bd01c601d501ef010e02;
    decBuf[1688] = 256'h2c023f024a0247023e022c0212020002ea01dc01d901d701d901e301ec01f401;
    decBuf[1689] = 256'hfb01fd01fe01ff01fe01fd01020208020a0216021b021f0221021d0215021202;
    decBuf[1690] = 256'h0802ff0100020602110224023c0252026b027602790270025e0249023a023202;
    decBuf[1691] = 256'h350248026a029402c602f60216033203370329031403f902d202c302b502b102;
    decBuf[1692] = 256'hc402dd02f9021c033c0349034d034903390325030803ed02dc02d202ca02d702;
    decBuf[1693] = 256'hec0206031f033b035603600364035b0353034c033d032f032a03250326032503;
    decBuf[1694] = 256'h21031e0319030f0308030003f802f702f402f002f102ee02e102d302c002a802;
    decBuf[1695] = 256'h98028a0282028e029d02b702d602f402080319031c0314030603ec02c602ac02;
    decBuf[1696] = 256'h950288028c029702b302d602ff0227034b0358035d03510332031403f102d102;
    decBuf[1697] = 256'hc402cf02e10203032d03540378038f039403800361033a030203dd02ac029a02;
    decBuf[1698] = 256'h8902840288029e02a902bb02c402cd02cf02c802b9029f028702710251024502;
    decBuf[1699] = 256'h3902350239024102540264026f02750277026e025e0247022a020f02f001db01;
    decBuf[1700] = 256'hcf01cb01c801d101e301f9010d022402340237023a0229021202f501da01c901;
    decBuf[1701] = 256'hb901b601b901c501d401e601f201f401ee01e501d301be01af01a2019b019d01;
    decBuf[1702] = 256'ha301ac01bb01c101c601ce01d201d101d201d101cc01cd01c901c301bc01b101;
    decBuf[1703] = 256'ha6019e0192018a0188018401850189018a0189018d0192019401970198019901;
    decBuf[1704] = 256'h990192018c0185017a017101670163015d0159015401500148013c012d012301;
    decBuf[1705] = 256'h10010301f700ec00e600dd00dc00d700d600d200cc00c900ca00cf00d100d400;
    decBuf[1706] = 256'hd300d600d500cf00c900c100b400a6009c008f008b0080007c007b007a007f00;
    decBuf[1707] = 256'h860091009d00ac00b600bb00b900af009d008700730061005a00600072008c00;
    decBuf[1708] = 256'hac00c100d400d800c800ae0088005a002200fcffdaffc7ffcdffe6ff07002400;
    decBuf[1709] = 256'h470068006c00600048001f00f8ffcaff9eff82ff7dff81ff96ffb2ffd8fffcff;
    decBuf[1710] = 256'h130017000c00ecffc6ff98ff6cff45ff2bff1dff19ff25ff36ff46ff54ff5cff;
    decBuf[1711] = 256'h63ff61ff5fff5aff52ff4aff40ff35ff2bff21ff16ff0eff0dff13ff22ff34ff;
    decBuf[1712] = 256'h49ff63ff75ff7eff7bff6eff54ff2dff09ffe9fecbfeb0feadfeb6fec4fedcfe;
    decBuf[1713] = 256'hf8fe1bff32ff47ff4bff41ff25fffafed3feaffe98fe8bfe87fe99feb5fed0fe;
    decBuf[1714] = 256'heffe05ff10ff0dfff7fed1fea3fe78fe50fe37fe29fe2dfe39fe51fe6dfe88fe;
    decBuf[1715] = 256'ha1feb7fec5fed2fed9fedbfed9fed4feccfec8febefeb5feb4feb7febafec5fe;
    decBuf[1716] = 256'hd0fedbfee2fee3fee0fed5febefea2fe87fe6efe52fe37fe26fe23fe25fe38fe;
    decBuf[1717] = 256'h52fe71fe8ffeaafec3feccfec9febcfea2fe7cfe62fe42fe35fe31fe3bfe51fe;
    decBuf[1718] = 256'h71fe8ffeaafeb4feb7fea9fe91fe75fe5afe50fe46fe4ffe67fe83fea6fecffe;
    decBuf[1719] = 256'hebfe05ff13ff17ff1bff10ff07fff9fef1feeafee3fee5fee4fee5fee4fee2fe;
    decBuf[1720] = 256'hdcfed6fecbfec4febdfeb7febafebffec5fed2fee4fef0fefbfe01fffffefefe;
    decBuf[1721] = 256'hfcfef5fef6fe01ff0dff1fff2fff3eff44ff46ff3eff30ff1dff0bfffffef4fe;
    decBuf[1722] = 256'heafee9fee7fee5feeafeedfeeefef3fefafefefe06ff0bff0eff13ff15ff13ff;
    decBuf[1723] = 256'h0dff08ff00fffbfef8fef7fefdfe08ff14ff21ff2eff2fff31ff32ff2cff26ff;
    decBuf[1724] = 256'h23ff1aff10ff07fffffe00ff03ff07ff14ff32ff50ff6bff84ff93ff9cff94ff;
    decBuf[1725] = 256'h84ff70ff5eff44ff39ff30ff33ff3bff50ff6aff83ff9fffaaffb5ffb8ffaaff;
    decBuf[1726] = 256'h97ff78ff5bff38ff21ff0bff07ff19ff3bff65ff98ffc8fff3ff10000a00fdff;
    decBuf[1727] = 256'hd6ffa8ff7cff55ff3bff40ff4dff68ff95ffc1ffddffedfffbffeeffdaffbbff;
    decBuf[1728] = 256'h95ff71ff50ff44ff38ff3cff45ff53ff6bff87ff9affacffc2ffcaffc8ffcaff;
    decBuf[1729] = 256'hbbffa5ff91ff7aff64ff55ff53ff55ff5bff6dff83ff9dffb5ffd1ffe5fff6ff;
    decBuf[1730] = 256'hf9fff1ffd9ffb7ff96ff79ff65ff62ff71ff9cffd5ff09004700700087008e00;
    decBuf[1731] = 256'h6e0047001900e1ffacff98ff91ffadffd1ff040034006d0083008a0084006800;
    decBuf[1732] = 256'h44002300fdffe3ffd6ffd1ffddffeeff04001e00370046004f004c0040002900;
    decBuf[1733] = 256'h1300f9ffe8ffdeffd6ffdeffeafff8ff06000f0017001c001d00210027002c00;
    decBuf[1734] = 256'h320038003a003a003200250017000900f9fff3fff1fff9ff08001a002f003e00;
    decBuf[1735] = 256'h40003e0038002a001a000f0009000b00100014001e00240028002f0035003700;
    decBuf[1736] = 256'h3a00390035002d001e0010000400f9fff4fff0fff4fffcff0700110018001e00;
    decBuf[1737] = 256'h240025002200230027002f0037003e00440047003f0030001e000900f5ffe8ff;
    decBuf[1738] = 256'he5ffe8fff6ff02001000160015000d00fcffe5ffcfffbbffaeffa6ffa4ffaaff;
    decBuf[1739] = 256'hb7ffc8ffdefff8ff0900190021001f000e00f7ffdbffb8ffa1ff8bff78ff7cff;
    decBuf[1740] = 256'h7fff93ffa5ffbbffc9ffd1ffcaffb7ff9fff89ff6fff5eff54ff51ff54ff5bff;
    decBuf[1741] = 256'h5dff63ff69ff71ff78ff82ff8dff98ff96ff90ff7fff60ff42ff20fffffeeafe;
    decBuf[1742] = 256'hdefee2fef1fe11ff2fff4aff62ff72ff7bff73ff62ff4bff35ff1bff0aff00ff;
    decBuf[1743] = 256'h03ff0bff25ff3eff60ff8affa6ffbfffcdffc9ffb6ff8fff61ff29ff03ffe1fe;
    decBuf[1744] = 256'hdbfeebfe05ff2fff61ff84ff96ffa7ff98ff8aff6cff49ff29ff14ff00fffdfe;
    decBuf[1745] = 256'h06ff1aff37ff5aff7bff98ffacffb6ffadff99ff77ff56ff30ff16fffffefbfe;
    decBuf[1746] = 256'hfffe09ff2cff43ff61ff6cff70ff6dff64ff57ff50ff4eff50ff5cff6aff78ff;
    decBuf[1747] = 256'h7eff7fff78ff76ff75ff74ff7dff88ff93ffa2ffacffb1ffacff9fff8fff7cff;
    decBuf[1748] = 256'h6aff59ff5bff61ff71ff88ffabffcbfff1ff0b0019002500290026001c001400;
    decBuf[1749] = 256'h0700fbfff9ffffff0e00260042005d006f007e0076006800530033001e001300;
    decBuf[1750] = 256'h0f00180032004b0067007a008c00950092009500970099009f00ac00b400bb00;
    decBuf[1751] = 256'hbf00bc00af00a100930083007d007b0087009500a300b000b800b600b200a700;
    decBuf[1752] = 256'h9900910089008d009400a200b100c000ce00db00e300e700eb00e500dd00d600;
    decBuf[1753] = 256'hcb00bc00b200b000b200ba00c300ce00dc00e100e000de00d700d100d200db00;
    decBuf[1754] = 256'he600fa00110121012a0132012a01240116010601000106011201240139014e01;
    decBuf[1755] = 256'h5b015d015201400126010701fa00ee00f200fb000a011c013101460148014b01;
    decBuf[1756] = 256'h4d0143013d0132012501180113010c010d0116011e012b013b0145014b014a01;
    decBuf[1757] = 256'h41013701280116010f0104010201070113011d01270130013301300126011d01;
    decBuf[1758] = 256'h160115011a012401300135013a013b0135012f012a01260128012b0131013b01;
    decBuf[1759] = 256'h4401480150015301500150014d01470142013b012e0126011f011a011e012201;
    decBuf[1760] = 256'h2d013d0150015d01690167015d014d0136011a010601fc00f900fc0009011e01;
    decBuf[1761] = 256'h380143014c014901410131012601180108010201fc00f700fb0003010a011801;
    decBuf[1762] = 256'h2b01380149014f0151014f014401330120010e01fd00f300f500fa0005011301;
    decBuf[1763] = 256'h1b0124012801210116010e010201f700f200e900e000da00d300cb00c800c500;
    decBuf[1764] = 256'hc400c700cd00d600db00d900d600cd00ba00a30093007f006c006a006c006e00;
    decBuf[1765] = 256'h7a00860093009c00a100a2009e009300860076006700550044003e0038003600;
    decBuf[1766] = 256'h42004f005f0069006f006e00660052003500220009000000fdff050016002d00;
    decBuf[1767] = 256'h3d004b00530050004600380028001d0013000e001300180019001d001e001d00;
    decBuf[1768] = 256'h13000a0003000000fbfffaff0000060012001d002200230022001c0013000800;
    decBuf[1769] = 256'hfafff2fff0ffeefff3fff9ff01000a000b000800fbffe7ffcaffafff97ff87ff;
    decBuf[1770] = 256'h84ff87ff9cffb6ffcfffe5fff3fff0ffe4ffd1ffbaffaaff96ff93ff96ffa5ff;
    decBuf[1771] = 256'hb3ffc6ffd3ffd5ffcfffbdffa8ff99ff82ff72ff6fff72ff79ff83ff8dff9aff;
    decBuf[1772] = 256'h9fffa0ff9fff9bff98ff95ff94ff93ff95ffa1ffa9ffb3ffc0ffc8ffc9ffc8ff;
    decBuf[1773] = 256'hbdffacff99ff91ff8aff84ff8aff96ffa5ffb7ffc3ffc9ffcbffc6ffbaffadff;
    decBuf[1774] = 256'ha1ff9fff9dffa4ffb2ffc5ffd2ffe3ffe9ffe7ffe6ffdaffcaffbbffb1ffa5ff;
    decBuf[1775] = 256'h9dff9bff97ff9bff9cff9dffa1ffa4ff9fff9dff98ff94ff8eff88ff85ff84ff;
    decBuf[1776] = 256'h83ff8aff91ff99ffa0ffa6ffa9ffa6ffa0ff98ff93ff90ff8bff8bff91ff99ff;
    decBuf[1777] = 256'ha0ffa5ffa6ffa2ff9cff96ff8aff7fff77ff79ff7dff84ff8fff9dffa9ffb5ff;
    decBuf[1778] = 256'hb9ffbdffb9ffb4ffadffa3ff9aff93ff94ff97ffa1ffb0ffbeffcaffd6ffdaff;
    decBuf[1779] = 256'hd6ffcdffbdffa7ff99ff8cff85ff87ff91ff9dffafffc4ffd3ffe0ffe2ffdcff;
    decBuf[1780] = 256'hd6ffcdffc2ffbaffb9ffbcffc4ffcdffd6ffdeffe1ffdeffdcffd6ffcfffc9ff;
    decBuf[1781] = 256'hc5ffc1ffc1ffc2ffc3ffc4ffc7ffc6ffc1ffc1ffbaffb8ffbaffc1ffc8ffd7ff;
    decBuf[1782] = 256'he5fff5ff04000e000c000400f6ffe3ffcbffbcffadffa6ffa8ffb3ffc5ffdaff;
    decBuf[1783] = 256'he8fff5fff8fff1ffdfffcaffb6ffa4ff93ff91ff9bffb2ffc7ffe7ff05001800;
    decBuf[1784] = 256'h23002c0023001100fcffe2ffd0ffc1ffb8ffbbffc2ffd1ffe3fff3fffeff0400;
    decBuf[1785] = 256'h0600fefff6ffe7ffd9ffd0ffcbffc7ffceffd9ffe3fff0fffeff000002000100;
    decBuf[1786] = 256'hfcfff0ffe8ffddffd1ffc5ffbeffbaffb6ffb3ffb2ffafffacffabffaeffafff;
    decBuf[1787] = 256'hb0ffadffacffabffa5ff9fff9bff96ff94ff8fff8dff8aff89ff85ff81ff7eff;
    decBuf[1788] = 256'h76ff6cff62ff5aff4fff49ff40ff3cff3bff39ff34ff37ff38ff34ff2fff2dff;
    decBuf[1789] = 256'h2cff2bff2cff2dff31ff32ff36ff3bff3bff39ff36ff30ff28ff20ff17ff11ff;
    decBuf[1790] = 256'h0eff0dff0fff15ff1aff1eff23ff1eff1aff17ff0eff04fffefef8fef5fef6fe;
    decBuf[1791] = 256'hf9fefbfefafefdfefefefbfef5feedfee8fee1fed9fed3fed2fecffec9fec5fe;
    decBuf[1792] = 256'hc2fec0febbfeb9febbfebafebbfebefec2fec3fec2fec1fec1febcfeb3feacfe;
    decBuf[1793] = 256'ha8fea2fe9ffea2fea6feaefeb8febcfec0fec1febcfeb4feadfea4fe9dfe98fe;
    decBuf[1794] = 256'h93fe92fe96fe9bfea2feaafeb3febcfec2febffebefebbfeb7feb1feacfea6fe;
    decBuf[1795] = 256'ha7feaafeabfeb1febafec4fecffed7fedefee4fee7fee4fee0fedafed4fecdfe;
    decBuf[1796] = 256'hc7fec5fecbfed8fee6fef2fe04ff15ff1fff21ff1cff17ff10ff06fffbfef6fe;
    decBuf[1797] = 256'hf5fefbfe08ff13ff1dff2dff33ff34ff33ff28ff1cff10ff06ff02ff03ff0bff;
    decBuf[1798] = 256'h18ff28ff37ff45ff4dff4fff4dff49ff41ff3bff3aff39ff43ff52ff60ff6cff;
    decBuf[1799] = 256'h77ff7cff7dff77ff6dff61ff55ff4eff4fff55ff5fff71ff82ff95ffa2ffa9ff;
    decBuf[1800] = 256'habffa9ffa1ff99ff97ff96ff99ffa4ffb0ffc2ffd7ffe6ffedfff5fff7fff1ff;
    decBuf[1801] = 256'hebffe3ffd9ffd7ffd9ffdaffe1ffecfff8ff02000c00120015001c0021002700;
    decBuf[1802] = 256'h2d003700430048004f0056005500520051004e00480049004d00510059006300;
    decBuf[1803] = 256'h700078007900750072006a005d0054004c004a005400640077009400af00c100;
    decBuf[1804] = 256'hd000d900d600cf00bc00af009e00940092009400a200b400ca00de00f000fc00;
    decBuf[1805] = 256'hfe00f800f300e700d700cc00c600c800d000e100f4000b0121013b0146014f01;
    decBuf[1806] = 256'h52014a01430138012e0122012001220126012f01400150015f0171017d018301;
    decBuf[1807] = 256'h850180017f0177016d016c017001750182019401a401b701ca01d101d701d901;
    decBuf[1808] = 256'hd101c801c101b701b101b001b101bb01c401cf01e001eb01ed01f201ed01e801;
    decBuf[1809] = 256'he401e101db01de01e201e801f60104020c02140219021a02190213020e020c02;
    decBuf[1810] = 256'h09020c02120216021c0228022d022e02320231022b022a022802220224022902;
    decBuf[1811] = 256'h2a023002360238023f0243024002450246024102440245024402460247024602;
    decBuf[1812] = 256'h4b024d024b024f025202510259025c025b026002640260025f025c0252025402;
    decBuf[1813] = 256'h53024d02520255025702610268026b02730274026e026f026c0261025c025802;
    decBuf[1814] = 256'h54025202530254025c026002630269026a02690266025e0254024d0242023802;
    decBuf[1815] = 256'h33022d0228022b02310237023f02440247024c0247023e02340221020f02fe01;
    decBuf[1816] = 256'hf401ea01eb01f001f8010c021b0223022a02280216020502f201da01c401b601;
    decBuf[1817] = 256'hae01b501c001ce01e501f401fd010502f901ea01d801be01a501900187017f01;
    decBuf[1818] = 256'h8b019601a801b801c301c101c301ba01a4018e017a0168015c01550153015901;
    decBuf[1819] = 256'h5d0165016c016d0165015c014c013d012f012301170113011201130116011701;
    decBuf[1820] = 256'h1801190115010d010501fc00f300ed00e600e200df00d900d300cb00bf00b400;
    decBuf[1821] = 256'ha9009a008c0083007b0074006f006c0066005f00570052004b00430036002e00;
    decBuf[1822] = 256'h2a0023001f00190016000f000200f7ffecffddffcbffbfffb0ffa6ffa5ffa3ff;
    decBuf[1823] = 256'h9fff98ff91ff8cff83ff75ff6cff5eff54ff4eff50ff55ff59ff5fff65ff6aff;
    decBuf[1824] = 256'h69ff63ff57ff49ff37ff26ff1bff0dff05ff00ff01ff05ff04ff05ff00fffafe;
    decBuf[1825] = 256'hf0fee4fed5fecbfebffeb7feb3feb4feb3feb6febdfebefebbfebefebbfeb3fe;
    decBuf[1826] = 256'ha9fe9dfe92fe87fe78fe6afe5efe52fe45fe39fe30fe2cfe28fe24fe23fe24fe;
    decBuf[1827] = 256'h20fe1bfe15fe0dfe05fefcfdf1fde7fde0fddefde0fde3fde9fdebfdf0fdf1fd;
    decBuf[1828] = 256'hecfde6fddbfdc9fdbdfdaefda0fd97fd92fd91fd98fd9efda4fdadfdb0fdb2fd;
    decBuf[1829] = 256'hb3fdacfda6fda0fd9afd96fd95fd90fd91fd97fd9afd9dfda3fda0fda3fda5fd;
    decBuf[1830] = 256'ha3fd99fd95fd8cfd82fd7efd73fd6bfd6afd66fd65fd6afd69fd6efd75fd79fd;
    decBuf[1831] = 256'h7afd79fd73fd6dfd67fd5ffd59fd56fd57fd5bfd65fd6cfd75fd7cfd7dfd7bfd;
    decBuf[1832] = 256'h78fd70fd64fd59fd51fd4dfd4efd4dfd50fd5bfd60fd5ffd63fd5ffd57fd4efd;
    decBuf[1833] = 256'h48fd3efd3dfd39fd3efd47fd4bfd53fd5afd57fd55fd50fd47fd3dfd34fd2dfd;
    decBuf[1834] = 256'h2cfd2efd2ffd33fd3afd3afd3bfd3afd33fd2bfd26fd20fd19fd19fd1bfd21fd;
    decBuf[1835] = 256'h2bfd35fd40fd47fd4bfd4ffd4efd4bfd4cfd4dfd48fd49fd4efd4ffd51fd52fd;
    decBuf[1836] = 256'h4ffd52fd55fd52fd51fd54fd4ffd4ffd53fd50fd4ffd50fd4efd4ffd4ffd4ffd;
    decBuf[1837] = 256'h53fd5dfd63fd6cfd76fd7afd81fd82fd7bfd75fd70fd65fd5dfd5bfd57fd5bfd;
    decBuf[1838] = 256'h63fd68fd71fd78fd77fd78fd75fd68fd5efd59fd51fd52fd56fd5dfd69fd78fd;
    decBuf[1839] = 256'h86fd8efd93fd92fd8bfd85fd7afd71fd6dfd6efd73fd7ffd8afd94fd9efda7fd;
    decBuf[1840] = 256'ha8fda7fda1fd97fd93fd8dfd8cfd93fd9cfdabfdbdfdc9fdd4fddafdd8fdd0fd;
    decBuf[1841] = 256'hc9fdbffdb9fdbafdbbfdc1fdcefddcfdecfdfbfd01fe02fe01fef9fdf0fde9fd;
    decBuf[1842] = 256'he4fde3fde9fdf1fd02fe12fe21fe27fe30fe2bfe27fe20fe17fe0ffe10fe11fe;
    decBuf[1843] = 256'h1bfe27fe36fe48fe53fe5afe60fe65fe63fe5ffe5bfe5cfe64fe6dfe78fe89fe;
    decBuf[1844] = 256'h93fe9dfea6fea8fea3fe9afe91fe89fe88fe8bfe8ffe97fea5feaffeb8fec4fe;
    decBuf[1845] = 256'hc8fec4fec0febbfeb6feb3feb4feb8fec5fed7fee8fef7fe05ff07ff05fffdfe;
    decBuf[1846] = 256'heefee0fed8feccfecbfeccfed5fee3fef5fe01ff10ff16ff18ff1aff15ff0eff;
    decBuf[1847] = 256'h0aff09ff10ff1dff2bff42ff58ff66ff79ff85ff87ff85ff80ff7bff70ff6cff;
    decBuf[1848] = 256'h6dff73ff78ff83ff8fff9cffa5ffadffb2ffb3ffafffaeffabffaeffb7ffc1ff;
    decBuf[1849] = 256'hccffdaffe9fff8fffeff040002000000fafff1ffebffe6ffe9ffeafff0fff6ff;
    decBuf[1850] = 256'hfafffdfffefff8fff0ffe8ffe1ffdbffdaffe2ffeefffdff0b001e0030003800;
    decBuf[1851] = 256'h420040003b0033002b00240026002b0034004200520065007200790077006d00;
    decBuf[1852] = 256'h640056004c00430045004c005e0073008d00a600bc00ca00cd00ca00c000b600;
    decBuf[1853] = 256'had00a500a600b000c000d700ed0001010f01160114010a01fa00eb00e100d800;
    decBuf[1854] = 256'hd700e400f40007011f01340143014b014d014701410134013001340138014801;
    decBuf[1855] = 256'h600176019001a101b101b901b701ab01a4019a01920193019b01a701bc01d001;
    decBuf[1856] = 256'he301f301fe0100020202fa01ef01eb01ef01f401010215022c0242025c026702;
    decBuf[1857] = 256'h76027902760274026e02640265026a026f027e0290029c02ab02b502b602bb02;
    decBuf[1858] = 256'hba02b602b702ba02b902c302d202e002f3020603160329033c03480352035c03;
    decBuf[1859] = 256'h62036d037703810391039c03a203ae03bd03c303cc03d403db03e503ee03f303;
    decBuf[1860] = 256'hfe0309040a0415042304280437044904550463047504810494049c04a304ae04;
    decBuf[1861] = 256'hb004ae04b304b504b604bc04c004c304d004d604d404d904dd04dc04dd04e104;
    decBuf[1862] = 256'he004eb04fa0404051a0530053f0556056c0575057d0589058b05910599059b05;
    decBuf[1863] = 256'ha905b805c305d505e605ec05fa05030601060606040603060b0616061d062f06;
    decBuf[1864] = 256'h4506530670068306870696069f069c06a306a606a006a806b406b806c706d106;
    decBuf[1865] = 256'hd706e206e606e006e306de06d106d206d406d006df06ed06f206070715071807;
    decBuf[1866] = 256'h240726072007220723071f07290734073b074d075e0764077207770773077107;
    decBuf[1867] = 256'h6a075a075c075a0758076a077b078a07a007ae07b107b807b1079f0798078e07;
    decBuf[1868] = 256'h7c077907800782079507a207a907b807c207af07a20791077507620751074107;
    decBuf[1869] = 256'h4a07510754076707790777077d0777076107510737071f070f070607fe060a07;
    decBuf[1870] = 256'h19071f0732073a072e072c0722070c07fc06f306e106e306ea06ec06fb060607;
    decBuf[1871] = 256'h0c0711070c07fc06f106df06c506bb06b106a906ab06ae06ac06b206a9069406;
    decBuf[1872] = 256'h85066e0652063e062d061d062006230620062b062906200618060406e205cb05;
    decBuf[1873] = 256'ha505810573056605630566056f056d056f055f0547052b050005d904b5049504;
    decBuf[1874] = 256'h880484048f049804ac04bf04c104bf04ad04890465043c041404fb03e403df03;
    decBuf[1875] = 256'heb03fc030c04150417040204e803c2038903550325030503f402ef02f4020903;
    decBuf[1876] = 256'h1d0327032a031c03fa02d0029d026d02350210020902020208020d021b021f02;
    decBuf[1877] = 256'h1402fb01d901a60176013e010901e700d400ce00d300d800e500e900de00cf00;
    decBuf[1878] = 256'haf0089005b002f001300f9ffe2ffdeffe2ffdeffdbffd8ffcbffb6ff96ff70ff;
    decBuf[1879] = 256'h42ff22fffbfed7fec9feb4fea8fe9efe8efe80fe68fe46fe1cfef5fdd1fdb1fd;
    decBuf[1880] = 256'h93fd78fd5ffd56fd42fd2ffd1ffd03fde0fcc0fc91fc65fc49fc30fc0ffc02fc;
    decBuf[1881] = 256'heffbe5fbd5fbc1fba4fb89fb5bfb30fb08fbe4fabbfaaafa90fa8cfa87fa7cfa;
    decBuf[1882] = 256'h71fa6efa54fa35fa17faecf9c5f9a1f98af975f969f95ff95bf95ef951f941f9;
    decBuf[1883] = 256'h2df906f9dff8b1f885f852f830f811f8f4f7eff7e1f7ccf7c8f7b0f794f780f7;
    decBuf[1884] = 256'h53f727f70bf7e7f6c7f6baf69ff68df684f676f668f65df63df61cf607f6e4f5;
    decBuf[1885] = 256'hbbf59ef57bf55af545f522f50bf5fef4dbf4c4f4b7f4a4f48cf488f474f467f4;
    decBuf[1886] = 256'h65f452f43ff438f41df409f4fff3e3f3cff3d3f3bdf3b4f3b2f3a1f38ef381f3;
    decBuf[1887] = 256'h5df339f322f3f3f2c8f2b7f29df28ff293f288f28bf2a1f293f286f283f263f2;
    decBuf[1888] = 256'h43f236f20cf2f0f1eaf1ddf1d8f1ecf1e8f1ebf1f4f1e2f1c3f1b6f17cf153f1;
    decBuf[1889] = 256'h3cf10cf1f9f0f4f0eef0fcf01af11ef121f137f123f111f105f1e5f0c5f0c0f0;
    decBuf[1890] = 256'ha5f0a2f0bef0c2f0d3f0f6f0f1f0edf0f1f0caf0a6f098f06af04af045f02bf0;
    decBuf[1891] = 256'h30f045f051f062f078f075f06df070f050f02ff02bf010f006f015f012f01ff0;
    decBuf[1892] = 256'h3ef043f04ef060f04af036f02ef00ff0faeff6efe4efe1effbefffef14f034f0;
    decBuf[1893] = 256'h30f034f045f036f027f02ff023f025f03bf044f056f07af089f097f0acf0a9f0;
    decBuf[1894] = 256'ha5f0a8f09af097f0a8f0a6f0b4f0cef0e9f0fbf01df122f126f131f120f11df1;
    decBuf[1895] = 256'h25f11ef129f149f157f16cf197f1a8f1b7f1cef1caf1c6f1d1f1c1f1c4f1dcf1;
    decBuf[1896] = 256'hdff1f9f11ff239f259f27ff285f292f2a8f29cf2a0f2aff2a7f2b4f2cef2e6f2;
    decBuf[1897] = 256'h02f32df349f363f38cf392f3a1f3aff3b4f3b7f3d0f3d9f3f9f31ff443f463f4;
    decBuf[1898] = 256'h92f4b1f4cef4f1f4fff40cf527f52bf534f54ef55ff57cf5a6f5c2f5e6f510f6;
    decBuf[1899] = 256'h2cf646f666f673f686f69ff6a8f6c2f6e1f6f7f619f74cf76ff79af7c2f7e6f7;
    decBuf[1900] = 256'h06f82cf83cf853f871f884f89cf8bff8d6f8fcf82af93df964f993f9b2f9d9f9;
    decBuf[1901] = 256'hfdf914fa3afa5efa75fa9cfac0fae0fa0ffb3afb57fb85fbb0fbcdfbfbfb26fc;
    decBuf[1902] = 256'h43fc66fc90fcacfcd0fcf0fc0efd29fd49fd67fd91fdb9fddcfd06fe2dfe5cfe;
    decBuf[1903] = 256'h87feaffed3fef3fe11ff2cff4bff69ff8cffacffdbff070039006a009500bd00;
    decBuf[1904] = 256'heb000a0126014001570175018801af01dd0108023b026b02a302d80208033403;
    decBuf[1905] = 256'h500374038b03a903c403dc03ff03320454048c04d004fd0437055d058d05ac05;
    decBuf[1906] = 256'hc805d705f8050d06200647067506a106df0629075b078907c207d907fb071a08;
    decBuf[1907] = 256'h15082e083c08520874089e08d1080f0948097d09ad09d909ea09030a110a0d0a;
    decBuf[1908] = 256'h200a400a550a870ac50aee0a320b720b9b0bd00be40bea0bf00bf50bf10b0e0c;
    decBuf[1909] = 256'h290c420c710cbc0cee0c2e0d580d6e0d900da30d9e0dad0dbb0dbf0dea0d110e;
    decBuf[1910] = 256'h3f0e840ec40eed0e220f440f4a0f5b0f560f480f5d0f690f730f9c0fcf0ff10f;
    decBuf[1911] = 256'h29105e1080109f10bc10ac10ba10be10b310cb10e710fb102f1164118611be11;
    decBuf[1912] = 256'he411f8110b121c120d121112161202121b1231123f1266129912ae12d912f512;
    decBuf[1913] = 256'hfb1208130d13f212fc12f912f0120d1328133a1369139913ac13d313ed13df13;
    decBuf[1914] = 256'he313d713b813b413b0139e13c113d813ed1318143f1444145b1457143c143114;
    decBuf[1915] = 256'h1514f213f713fb13f7131e14421450147e1491148014901478144a1437142614;
    decBuf[1916] = 256'h021407141414171437144c145014621465143f143a141a14eb13e513d413c513;
    decBuf[1917] = 256'hd213df13db13fb130814f413f813e813c313b3139c1376137b136d1360137413;
    decBuf[1918] = 256'h7013611369135c133d1331131d13f012e912d912b512b912ad1291129c128c12;
    decBuf[1919] = 256'h6d12681255122f121f121112eb11e611d811ba11b611a51183117e1169113e11;
    decBuf[1920] = 256'h2d111e11f410ef10df10b610b010a110771071104d102d1020100510df0fda0f;
    decBuf[1921] = 256'hcc0fae0faa0f990f700f6a0f460f1d0f0c0ff20ec90ec30eb40e930e8f0e830e;
    decBuf[1922] = 256'h640e570e340e010edf0dc00d820d690d530d300d370d260d160d1b0d060de30c;
    decBuf[1923] = 256'hc20c9c0c640c3e0c0e0cd60bce0bba0ba70bad0bb20ba40b970b7c0b480b130b;
    decBuf[1924] = 256'hd50a8b0a590a2b0af209ea09e309e909fa09f509e709d209a7096a091f09d908;
    decBuf[1925] = 256'h990860083a0826082c08310837084e0841082608f807b40761071407ba067e06;
    decBuf[1926] = 256'h5d063f0636063e0645064c06530636060806d0058d052805e504a90472045404;
    decBuf[1927] = 256'h5d0455046b0472046c045b042d04e803a8035e030403c70290025e0255024d02;
    decBuf[1928] = 256'h54025b026102510237020402c6017c013601e400ad008f006100590060006700;
    decBuf[1929] = 256'h6e0068004e002e00f7ffb3ff61ff14ffcefea0fe77fe61fe68fe6efe73fe79fe;
    decBuf[1930] = 256'h6bfe4dfe1bfeddfd92fd38fdfcfcaffc7dfc61fc59fc61fc68fc7afc75fc65fc;
    decBuf[1931] = 256'h3cfcfefbb4fb6efb1bfbcefa9cfa81fa79fa80fa87fa8dfa9efa85fa64fa2dfa;
    decBuf[1932] = 256'hdbf98ef948f9f5f8bef8a0f897f88ff8a6f8acf8b3f8adf87ff853f815f8cbf7;
    decBuf[1933] = 256'h85f757f71ef7f8f6f1f6ebf6f1f6f6f6f1f6dcf6c1f693f64ff621f6d7f5a5f5;
    decBuf[1934] = 256'h77f54ef537f530f52af519f514f5fdf4d7f4bdf48af45af43bf408f4d8f3d2f3;
    decBuf[1935] = 256'habf39bf397f379f35ef34cf31df3edf2cef29bf279f25af232f20ef201f2e3f1;
    decBuf[1936] = 256'hc8f1b6f18ef166f157f124f102f1eff0bcf0a8f0a1f085f076f071f053f038f0;
    decBuf[1937] = 256'h20f0f1efc1efa2ef6fef3fef2cef10eff6eefbeeddeed2eed5eeb3ee92ee7dee;
    decBuf[1938] = 256'h4bee1beefbedc9eda6edaded90ed96edadeda0ed9ceda0ed7ded5ded3fed05ed;
    decBuf[1939] = 256'hcbecb5ec85ec72ec83ec73ec78ec9eec8fec8aec8eec64ec3cec23ece7ebbdeb;
    decBuf[1940] = 256'hb6eba1eb9bebb7ebb2ebc0ebd5ebcaebb8ebb5eb8aeb6beb5aeb36eb1feb23eb;
    decBuf[1941] = 256'h17eb1beb37eb33eb37eb46eb2ceb1beb1eebfeeaf2eafdeaeceae9ea02ebf1ea;
    decBuf[1942] = 256'heeea02ebeaeadbeae3eac6eabbeacceac3eacceaf3eaf9eafeea1eeb11eb06eb;
    decBuf[1943] = 256'h09ebe7ead9eaddead2eae3ea0ceb1deb36eb69eb70eb76eb87eb63eb43eb3feb;
    decBuf[1944] = 256'h0cebf8ea0aeb10eb34eb79eb97ebd7eb11ec18ec1fec32ec0becf1ebe3ebc5eb;
    decBuf[1945] = 256'hc9ebe9ebfeeb30ec7cecaeecc9ec03edfcecf5eceeecbcec99ec93ec82ec87ec;
    decBuf[1946] = 256'hbaecddec15ed67ed88edbaede8edf0edf8edf1edd2edcceddbedd7edeced1eee;
    decBuf[1947] = 256'h41ee79eeaeeed0eee3eeffeeefeeebeef8eedceed9eeefeef7ee0fef3eef60ef;
    decBuf[1948] = 256'h80efbdefd6effcef2cf032f04ef072f077f094f0b7f0c5f0d2f0f5f0f9f00ff1;
    decBuf[1949] = 256'h32f136f154f17ff19bf1bff1e8f1f9f11df234f238f24cf264f267f27bf2a3f2;
    decBuf[1950] = 256'hcaf203f346f386f3c0f303f41ff448f45ef457f451f462f45df474f49af4bef4;
    decBuf[1951] = 256'hfaf445f577f5a4f5def503f618f62bf630f636f64df662f68df6caf604f748f7;
    decBuf[1952] = 256'h9af7d1f703f830f849f860f874f87bf88bf8a5f8c5f8f4f82cf952f990f9caf9;
    decBuf[1953] = 256'heff911fa31fa42fa65fa7dfaa3fad1fa09fb3efb89fbbbfbfbfb24fc3bfc50fc;
    decBuf[1954] = 256'h62fc73fc83fca3fcd2fcfdfc47fd8dfdccfd17fe49fe64fe6cfe74fe6dfe67fe;
    decBuf[1955] = 256'h78fe91fec4fe10ff6affd7ff3e008100be00df00e900cd00b4008f007a008100;
    decBuf[1956] = 256'ha800f5005801d0016202c5021e032e033d031503d802a10283027a029302e502;
    decBuf[1957] = 256'h5e03f103a10418058405bf05ad057c053305d50480045f04690497040205a405;
    decBuf[1958] = 256'h3c06ec066307a407df07a90758070e07b006740669068706eb067e072f08d508;
    decBuf[1959] = 256'h6d09cf09e109d00987090e09bd08560813081f086c08da087c093f0ac10a380b;
    decBuf[1960] = 256'h790b8d0b7b0b2a0bc20a650a400a1f0a510ab60a2e0be10b870cc80c2a0d3c0d;
    decBuf[1961] = 256'h2c0de20c9f0c320ce80bdb0bcf0b1c0c8a0cf10c840d0d0e430e940ea30e600e;
    decBuf[1962] = 256'h3c0e050ed30db70dc00de50d310e9f0ee90e610f920fbe0fe60fc20f8b0f6d0f;
    decBuf[1963] = 256'h3f0f260f2e0f420f6e0fc30f17104e109410c210ca10d210cb10ac10a610a110;
    decBuf[1964] = 256'h9c10c310e61007113e11641178119711921182117e1171115e116f117f118d11;
    decBuf[1965] = 256'hb511e711ee111a122b121b1220121312f81103120612fd112412411250127012;
    decBuf[1966] = 256'h86128212851276124a12441228120e12261232123e1272129812ad12cc12dd12;
    decBuf[1967] = 256'hcd12c912b312891278125e1247125412601263128c12a812ad12c412c0129d12;
    decBuf[1968] = 256'h98127b12481234122d121c122c12431258128b12ad12c012dc12e112c112b412;
    decBuf[1969] = 256'h91125e123c122912021207121512101233124112451259125512331225120712;
    decBuf[1970] = 256'hd511ce11bb11aa11c411e411f111231246124c125d1258122e121212ee11a911;
    decBuf[1971] = 256'h8b116f1146113f1146113f115b11751170117d11721152113d111a11f010df10;
    decBuf[1972] = 256'hd010b910ce10e210f3101c1138113d11421135110211e0109b105b102210fc0f;
    decBuf[1973] = 256'hcc0fd20fd80fd30ff30f081005100f10ff0fd40fb50f8e0f4b0f300f170f000f;
    decBuf[1974] = 256'h150f280f390f670f7a0f740f6f0f4e0f0f0fcf0e850e2b0e060ecf0d9d0da60d;
    decBuf[1975] = 256'hbf0dc70de90dfc0df60dfb0dd20d940d5a0d160dd70c9d0c860c720c840ca10c;
    decBuf[1976] = 256'hba0cdb0cf00cdc0cc40c950c2e0ce40b870b190bed0ac50aa10ac20ae00afb0a;
    decBuf[1977] = 256'h140b2a0b080be90aa00a460af1098e094b09260905090f093d0966097d099f09;
    decBuf[1978] = 256'h990966092809ce086108f9079c075f073e0734074f0779078f07a407b7079a07;
    decBuf[1979] = 256'h62071007ad064f06fa05ad058f0586058e05a505d505e805e205d305a9056005;
    decBuf[1980] = 256'h1a05b50458041b04fa03dc03e503ee03f5030a041004ff03db03a8035d031703;
    decBuf[1981] = 256'hd7028d025b023f0226021f0218021e0219020902e901c30195015c012801f800;
    decBuf[1982] = 256'hbf009a00780065005f00500039002c000900e9ffbaff8eff5cff1efff4fec0fe;
    decBuf[1983] = 256'h90fe64fe48fe24fe04feeefdd3fdb4fd96fd73fd4afd22fdfefcd5fcb9fc95fc;
    decBuf[1984] = 256'h6bfc4ffc2bfc0bfcedfbc2fb9bfb77fb44fb14fbe8fab6fa86fa5afa32fa04fa;
    decBuf[1985] = 256'he5f9bef99af979f94bf91ff903f9dff8b5f899f880f85ff84af827f807f8e9f7;
    decBuf[1986] = 256'hc6f79cf775f73df708f7e6f6aef679f664f639f611f602f6e2f5c4f5b0f58af5;
    decBuf[1987] = 256'h66f54ff520f5f4f4cdf49ff480f46ff44bf43df439f425f41bf412f4f2f3ccf3;
    decBuf[1988] = 256'hb2f376f33cf317f3d9f29ff289f274f261f267f262f266f273f258f23ff22af2;
    decBuf[1989] = 256'hfef1baf18cf163f12ef127f115f11af134f139f13df150f13ff11cf105f1c5f0;
    decBuf[1990] = 256'h86f04cf017f0f5efefefe9efeeef18f034f043f064f057f03cf02af0fbefb0ef;
    decBuf[1991] = 256'h92ef52ef39ef41ef3aef4def74ef83ef9aefb8efa5ef85ef70ef36ef0defe7ee;
    decBuf[1992] = 256'hc5eea6eeb6eebceedcee0bef1def3aef5def50ef43ef2feffbeec6eeb2ee86ee;
    decBuf[1993] = 256'h75ee85ee80ee95eeb8eec6eedbeef6eee5eed5eecdeea5ee89ee7aee63ee5eee;
    decBuf[1994] = 256'h79ee7dee93eebeeed1eee2eefbeee4eee0eedceebceea7eea3ee8bee88ee96ee;
    decBuf[1995] = 256'h93ee9beeb6eeb2eebdeed3eecaeecdeeddeed7eeddeef4eef7eeffee17ef14ef;
    decBuf[1996] = 256'h1def2fef28ef2eef44ef47ef54ef78ef7def94efa9efa5efa9efb9efa4ef9def;
    decBuf[1997] = 256'h9fef94ef9eefb9efcceff2ef2bf050f073f09ef0a4f0b3f0c1f0acf0a0f0abf0;
    decBuf[1998] = 256'ha2f0b0f0d2f0e9f018f150f176f1a6f1c5f1d6f1d1f1d5f1c0f1adf1b7f1a8f1;
    decBuf[1999] = 256'hb0f1d8f1fff12df27ef2b5f2e7f215f32ef335f34af32bf31af31ff311f31ef3;
    decBuf[2000] = 256'h41f361f398f3dcf31cf455f48af491f4a4f4a9f485f477f46bf457f462f484f4;
    decBuf[2001] = 256'haef4e0f42cf572f5b2f5ecf502f609f60ff6fef5eff5eaf5def5e2f50ff62ef6;
    decBuf[2002] = 256'h6cf6b6f6e8f628f762f779f77ff786f775f765f758f753f75ff77ef7a5f7ddf7;
    decBuf[2003] = 256'h21f84ef888f8cbf8d5f8edf804f9fdf8f7f8fcf8f7f805f92bf94ff982f9c0f9;
    decBuf[2004] = 256'he9f91efa4efa6dfa7efa8dfa7ffa84fa88fa84fa94fab3fad1fafcfa2efb5efb;
    decBuf[2005] = 256'h8afbb2fbd5fbedfb02fc06fc10fc20fc34fc4cfc6efc8efcbdfce9fc05fd29fd;
    decBuf[2006] = 256'h49fd5efd72fd83fd93fda7fdbffdd5fdfafd14fe34fe5afe74fe8bfea0febbfe;
    decBuf[2007] = 256'hcdfee9fe04ff2bff4eff78ff9fffceffedff0900230030003d00490053006900;
    decBuf[2008] = 256'h8900a700d9000901350167018a01a901ba01c901ce01d201d601e101f6011c02;
    decBuf[2009] = 256'h4a028202b702f5021e03430366036c0372036c0371036d0371038903ac03d503;
    decBuf[2010] = 256'h080446047f04b404d604e904fa04ff04f104e404e104dd04ed040c0533056b05;
    decBuf[2011] = 256'h9f05dd0507062c06410647064d063d062f0623061f06300653067306aa06df06;
    decBuf[2012] = 256'h0f0747076d0773077a0774075a07560749073d074f0765077f07ac07e4070a08;
    decBuf[2013] = 256'h2c084c085c08620866085908560852084f085d087a089508bc08ea0809093109;
    decBuf[2014] = 256'h4a094f095c095f095509520955094d095909680976099009ba09cb09ef09060a;
    decBuf[2015] = 256'h130a260a310a2e0a3c0a440a4b0a5a0a700a790a960ab10abb0ad70aeb0aee0a;
    decBuf[2016] = 256'h040b0d0b0f0b200b2b0b310b400b4f0b510b610b6c0b6e0b810b8e0b950bb10b;
    decBuf[2017] = 256'hcc0bdd0bf90b1c0c210c3f0c4a0c470c500c4d0c3b0c420c4d0c4f0c690c8c0c;
    decBuf[2018] = 256'h9a0cc80ce80ced0c070d0c0df60cf20ce80cd20cdb0ce80cef0c0f0d420d640d;
    decBuf[2019] = 256'h9c0dc20dc90dcf0dd50dbb0dad0d980d840d880d910d9a0dc10de90d020e2c0e;
    decBuf[2020] = 256'h480e4d0e5b0e570e430e400e300e220e2a0e3a0e410e5f0e850e940ebe0ecf0e;
    decBuf[2021] = 256'hd40ee20ede0ed20ecf0ec50eb10eb90ebb0eb50ecb0ed90ee10efb0e140f170f;
    decBuf[2022] = 256'h2b0f380f2c0f3b0f390f260f2e0f270f180f1e0f230f1b0f310f3b0f3e0f550f;
    decBuf[2023] = 256'h5f0f560f630f610f490f460f380f200f1d0f1a0f0d0f1e0f2d0f2f0f490f640f;
    decBuf[2024] = 256'h680f770f7a0f680f650f560f380f230f180ff80efc0e000ffd0e190f2c0f300f;
    decBuf[2025] = 256'h460f4e0f410f3f0f2c0f040ff30eda0eb90ebe0ec10ebe0ee00ef70e040f270f;
    decBuf[2026] = 256'h350f280f1d0f040fd50eb30e940e6c0e5d0e580e5c0e780e900ea60ec60ed20e;
    decBuf[2027] = 256'hc70ec30ea70e750e600e340e0d0e080e030eff0d1a0e330e3c0e560e590e4a0e;
    decBuf[2028] = 256'h3b0e190ee60dc40d980d660d510d4b0d450d540d620d670d820d850d6f0d670d;
    decBuf[2029] = 256'h4a0d1f0d030dd50ca90c980c890c720c760c7a0c6f0c730c700c580c4f0c350c;
    decBuf[2030] = 256'h0e0cf50bd40ba60b930b770b5d0b580b4c0b380b350b2b0b170b0f0bff0adf0a;
    decBuf[2031] = 256'hd10aab0a870a670a400a120af309d709b309a50998098509810978095e095409;
    decBuf[2032] = 256'h3e091e090009d608a308810855082e081e080708f207ee07e407ce07bf07a207;
    decBuf[2033] = 256'h78075c072307ef06bf06860661063f061f060e060906fb05ef05eb05d905b705;
    decBuf[2034] = 256'ha005710539051305d5049c047604460427041604fc03ee03ea03d703be03a203;
    decBuf[2035] = 256'h780345030703cd028a025c022202fd01e801e201dc01e201dd01d901c501a601;
    decBuf[2036] = 256'h6f012b01d9008c0046000600ccffa7ff92ff8cff92ff8cff88ff7bff50ff1eff;
    decBuf[2037] = 256'he0fe96fe3cfefffdb2fd80fd65fd5cfd64fd6bfd71fd6bfd5cfd32fd0bfdbefc;
    decBuf[2038] = 256'h5bfc18fcc3fb76fb30fb15fbfcfaf5fafcfaf5fafbfaecfacbfaa5fa62fa10fa;
    decBuf[2039] = 256'hc3f97df92bf9f4f8d6f8bbf8b3f8baf8b3f8c6f8aaf890f867f81df8d7f785f7;
    decBuf[2040] = 256'h22f7dff6a3f66cf64ef657f64ff656f65df64af639f616f6d9f5a0f55cf50af5;
    decBuf[2041] = 256'hd3f4a1f473f45bf462f44ef447f44df433f413f4f5f3bbf371f33ff3fff2c5f2;
    decBuf[2042] = 256'haff27ff26cf266f257f249f245f22af211f2fbf1d0f1a4f188f150f12af116f1;
    decBuf[2043] = 256'heaf0cef0bef095f079f069f040f024f014f0ebefceefbfef9fef81ef75ef4fef;
    decBuf[2044] = 256'h2bef14efe5eec6eeb5ee91ee71ee75ee5aee4fee59ee3fee2dee24eef9edcded;
    decBuf[2045] = 256'hb1ed79ed53ed3eed1fed0eed13ed0fed13ed26ed1ced19ed16edefecc7ecb8ec;
    decBuf[2046] = 256'h85ec63ec50ec34ec2fec46ec41ec45ec65ec58ec54ec58ec2fec08ecf8ebc5eb;
    decBuf[2047] = 256'ha3eb90eb74eb6feb86eb82eb95ebb5eba8ebacebb6eb94eb74eb67eb35eb12eb;
    decBuf[2048] = 256'h0cebf0eae0eaf8eaebeae7ea06eb02ebfeea10ebfaeaeceaf3ead0eab6eabbea;
    decBuf[2049] = 256'h95ea85ea93ea86ea8aeaaaeaa5eab9ead8ead4ead8eae9eacdeabaeab6ea8eea;
    decBuf[2050] = 256'h7dea82ea6bea78ea9beaa8eac6eaf9ea0deb20eb3ceb2deb1feb23ebf8eae8ea;
    decBuf[2051] = 256'hedeadfeaecea1eeb33eb5eeb9cebb5ebdaebefebe9ebd8ebddebb3eba3eba8eb;
    decBuf[2052] = 256'ha3ebb8ebebeb0dec45ec89eca4eccdecf3ececece6ecebecd2ecc4ecd1eccdec;
    decBuf[2053] = 256'hdeec0ded30ed5beda4edc2eddeed07eef1edf7edfeede2eddcedeaede6ed09ee;
    decBuf[2054] = 256'h3cee5eee96eedaeef5ee1fef44ef4bef51ef57ef47ef4cef61ef65ef85efbcef;
    decBuf[2055] = 256'he1ef12f056f072f09bf0cff0d6f0e9f005f115f12cf152f176f19ff1e9f11bf2;
    decBuf[2056] = 256'h48f292f2b0f2def218f32ef343f36ff38bf3aff3ebf314f449f479f4a4f4d7f4;
    decBuf[2057] = 256'h15f52ef562f592f5b2f5e4f514f640f673f6b1f6daf60ef73ef75ef785f7b3f7;
    decBuf[2058] = 256'hc6f7edf71bf847f86ff8a7f8ccf8fdf828f950f969f993f9a4f9bdf9def9fcf9;
    decBuf[2059] = 256'h26fa59fa89fac1faf6fa34fb5dfb91fba6fbc5fbe1fbf1fb11fc2ffc4afc77fc;
    decBuf[2060] = 256'hb0fce4fc14fd4dfd81fdb1fdd0fdedfd06fe27fe3cfe5ffe88febbfeebfe30ff;
    decBuf[2061] = 256'h70ffbaffecff2c0055007b008f00ae00bf00d90003012a016201a601e6011f02;
    decBuf[2062] = 256'h54028402b002cc02e602fd021a03360363038f03c103ff0339046e049e04c904;
    decBuf[2063] = 256'he604f5040c0519052c054c0569059405c705f7052306550678068a06a606ac06;
    decBuf[2064] = 256'hb006bd06c906e1060a07310769079e07ce0706082c0833085208580852086a08;
    decBuf[2065] = 256'h7f088a08b808f008250963099c09d109010a2d0a3e0a570a6e0a7b0a9e0ac80a;
    decBuf[2066] = 256'hef0a320b710bab0bef0b410c620ca80cd50cee0c140d360d550d7d0dab0dd70d;
    decBuf[2067] = 256'h140e4e0e740ebf0ef10e1f0f590f8d0fa20fce0ff50f0f102f10551065108510;
    decBuf[2068] = 256'hab10b010da100111111131114f115a1173118911801193119a118b1195119a11;
    decBuf[2069] = 256'h8b119d11a911a711c111d311d011de11e611d511d711cd11b311af11a5118f11;
    decBuf[2070] = 256'h9711a5119911b411c811c411da11e811db11e211dc11c211cd11c911bb11d311;
    decBuf[2071] = 256'hef11fa11211245125c1282129c129712a412a8129612a012a812a012c412e812;
    decBuf[2072] = 256'hf6122d13621368139413b013ab13b913bd13aa13b413be13bb13e2130a141914;
    decBuf[2073] = 256'h4c146e1468148f1495147414701464143e14391434141f143a144b144f146e14;
    decBuf[2074] = 256'h7b14681472146214371431141514e713ed13e713ce13ee13fb13f71310140c14;
    decBuf[2075] = 256'hf813f613e513c513b713a2138f13a013b013b313da130114071427142b141814;
    decBuf[2076] = 256'h22141f1405141714261435145c149a14c314071534154d1573157a1567156c15;
    decBuf[2077] = 256'h72155a158115a515bc15fb154e166f16b516d016d816e016cb169f168e167516;
    decBuf[2078] = 256'h54166a167d168816b616d916df16f016e116a4167b162916dc15961556151c15;
    decBuf[2079] = 256'h0615f114de14e414ca14a11479143714d21375132013a71255120c12ae11a211;
    decBuf[2080] = 256'h6b11391130110711c31095104b10f10fb50f520ff40ed00e990e670e4b0e320e;
    decBuf[2081] = 256'h1c0e150e020edb0dd60db50d870d740d4d0d1e0d180dfc0ce20ce70ceb0ce00c;
    decBuf[2082] = 256'hf80c020dff0c160d190d110d190d120dfe0cfc0cf00cdd0ce50ce20ce00cf60c;
    decBuf[2083] = 256'h050d0c0d220d250d1d0d1a0d070de50cce0ca80c7a0c670c400c260c180c030c;
    decBuf[2084] = 256'he80bdd0bc70b9c0b7d0b560b130be50a9b0a690a290a000abc09a10978094309;
    decBuf[2085] = 256'h21090209cf08ad08740831080308ca07860758071f07db06c006970671065c06;
    decBuf[2086] = 256'h3d062c061d060606f105dd05c505a2058b056d054b053d052705240527052a05;
    decBuf[2087] = 256'h3305400547054d0553054b053c052e051705fb04e804d604c704be04bb04be04;
    decBuf[2088] = 256'hc004ba04b504ad04990477044d041b04eb03a60366032c03f802c8029c026902;
    decBuf[2089] = 256'h39020102cc0181012701d2006f0011008cff0fffbdfe56fedefd8dfd43fde5fc;
    decBuf[2090] = 256'ha9fc46fce8fb93fb46fbc4fa6bfaf9f974f91bf9a9f85ff802f8c5f78ef75cf7;
    decBuf[2091] = 256'h2ef7f5f6cff691f658f623f6d7f591f564f52af505f5f0f4ddf4d8f4e7f4ecf4;
    decBuf[2092] = 256'hf8f413f517f51af51df50bf5faf4f8f4e6f4dff4f2f4faf414f541f561f588f5;
    decBuf[2093] = 256'hacf5c3f5d0f5dbf5d1f5bbf5b2f59bf58bf588f57bf57df58cf586f588f590f5;
    decBuf[2094] = 256'h7df565f54ff524f5ecf4c6f488f44ff429f4ebf3b2f38cf35cf324f3fef2c0f2;
    decBuf[2095] = 256'h87f261f223f2d9f1a7f167f11df1d7f085f038f006f0c6ef7cef5eef1eeff4ee;
    decBuf[2096] = 256'hedeecbeeabee9aee6cee41ee24eeecedb8eda3ed77ed66ed76ed71ed86eda9ed;
    decBuf[2097] = 256'hc0edd6edf1edededeaedededd0edbdedc0edb1edb9ede1edfded2bee70ee8bee;
    decBuf[2098] = 256'hb4eedaeee1eedaeee0eec6eea6eeaaee87ee83ee98ee94ee9feec1eebceeb0ee;
    decBuf[2099] = 256'hb3ee7fee4aee1aeebded5fed22edd5ec8fec62ec28ecf3ebdfeba7eb72eb42eb;
    decBuf[2100] = 256'he4ea87ea32eab9e947e9fde8a0e832e806e8c3e787e766e734e7f4e6dbe689e6;
    decBuf[2101] = 256'h3ce60ae6b7e56ae538e5f9e4cfe4d7e4b4e4bbe4d7e4d2e4e0e406e50be519e5;
    decBuf[2102] = 256'h37e53ae54ce57be58fe5afe5f8e516e656e6b0e6d5e622e77ce7b8e7efe749e8;
    decBuf[2103] = 256'h86e8bde817e954e98be9d1e9fee938ea8beaaceadeea30eb67ebadebffeb20ec;
    decBuf[2104] = 256'h52ec92ec9aeca1ecb6eca3ec92ec98ec80ec7cec90ec85ec8eecaeecaaeca6ec;
    decBuf[2105] = 256'ha9ec7bec4aec2becd7eb9aeb63eb1debf0eae7eac2eabbeac1eab0eaa1ea9cea;
    decBuf[2106] = 256'h65ea40ea0feacbe98be972e93ee929e93ce941e95be98ee9a2e9cee9f6e905ea;
    decBuf[2107] = 256'h0aea1fea1bea1eea41ea4fea75eac2ea0feb55ebcbeb1dec84ece2ec1eed55ed;
    decBuf[2108] = 256'hafedd4ed0bee51ee90eedbee49ef92ef0bf07df0e4f041f196f1e3f115f255f2;
    decBuf[2109] = 256'h7ef2a4f2d4f2f3f21bf35df38bf3b4f3f8f313f43cf462f469f47bf48cf47df4;
    decBuf[2110] = 256'h8bf498f484f488f497f489f48cf48ef47ff479f47bf469f462f464f452f44bf4;
    decBuf[2111] = 256'h4df43bf434f432f41cf419f41bf419f428f446f464f48ef4ccf4f5f439f579f5;
    decBuf[2112] = 256'ha2f5d7f507f626f659f696f6d0f614f778f7d6f743f8c8f821f993f9faf958fa;
    decBuf[2113] = 256'hacfaf9fa3ffb7ffbdafb2ffc92fc0afd7cfd01fe7efef0fe74ffceffffff4800;
    decBuf[2114] = 256'h8b00b000d100030130016a01ad01ed0138027e029902c202d902d202bf02ae02;
    decBuf[2115] = 256'h8a0273026602530257025a025d025f02580249022f020902db01a2016e013001;
    decBuf[2116] = 256'h0701d200b0009100740065004e0039001e00feffe0ffc5ffa6ff90ff7dff7aff;
    decBuf[2117] = 256'h70ff79ff86ff92ffa9ffbfffd3fff0ff13002a0050008900ae00ec0026016901;
    decBuf[2118] = 256'ha901e30126027902c6020c035e03c1031e047304ec043d05a50502065706ba06;
    decBuf[2119] = 256'hfd0652079f07f9074e089b0809095309b0091d0a670aaa0aff0a200b660b930b;
    decBuf[2120] = 256'hbd0bf10b210c410c7e0cb80cde0c0e0d460d5d0d7f0d9e0da40db30db80db40d;
    decBuf[2121] = 256'hc70dd10dce0de20dfa0d030e1d0e360e390e530e640e610e810e8e0e910eb80e;
    decBuf[2122] = 256'hdc0eea0e210f460f690fa10fd60ff80f301056106a10a310d710f9103e116c11;
    decBuf[2123] = 256'h9511e81135126712b912061338137813c213f41334146d149314df1425155215;
    decBuf[2124] = 256'h8c15c015e3150f162b1626163316381624162816251611161e161b1604160116;
    decBuf[2125] = 256'he715b2158d154115e714ab144814ea13ad1360131a13db12a1124e1201129311;
    decBuf[2126] = 256'h2c11b4102110980ff70e8b0e020e850d130dac0c690c140cb10b530be60a610a;
    decBuf[2127] = 256'h080a7609140996084508fb07d3079707760758073c071307ee06cb0686066b06;
    decBuf[2128] = 256'h42061c0615061c061606440670068c06c406f9061b0754078807aa07ef072f08;
    decBuf[2129] = 256'h5808ba0817095409b709150a510ab40a120b4f0bb20b0f0c640cc70c3f0d910d;
    decBuf[2130] = 256'hf80d560e920ef50e380f750fc20f08104810a210f7102e118811dd1114125a12;
    decBuf[2131] = 256'h88129012b512ca12d012ec12101327135f139313c313081436144e1474147b14;
    decBuf[2132] = 256'h68146e1469145114671482148c14bb140715251565158e15a415b915bf15ae15;
    decBuf[2133] = 256'hb415af159a15bd15dd15fb1535169016b41617173f1763178417a2179917a217;
    decBuf[2134] = 256'ha917a217c117de17ed1720184218481870187f1868186c1849180d18f517c017;
    decBuf[2135] = 256'h7417561729170017da16b8167f165a161c16d21578150b15a3142b1499130f13;
    decBuf[2136] = 256'h921200127711d6103e10b50f380fa60ef50d7e0dbc0c050c5f0b9c0ae5093f09;
    decBuf[2137] = 256'h7c08c5071f075c06da0534059c04ec037503dd022d02b601f3007100cbff33ff;
    decBuf[2138] = 256'haafe2dfebbfd54fdf6fc89fc3ffcfcfbc0fb89fb6bfb3dfb14fbeefaccfaadfa;
    decBuf[2139] = 256'h9cfa8cfa88fa9dfac0faeafa27fb72fbb8fb0afc57fc89fcc9fc02fd37fd67fd;
    decBuf[2140] = 256'hacfdecfd46feccfe49ffbbff5d00f4007e01fb016d02d40231038603d3032d04;
    decBuf[2141] = 256'h8204e5045e05f0057906f6068907eb076808b908e50828094d096e09a009df09;
    decBuf[2142] = 256'h2a0a980ae10a5a0bab0b120c550c7a0c9b0ca50cae0cb60cbd0cd20cf10c190d;
    decBuf[2143] = 256'h510d860dc30dfd0d230e450e580e5d0e6d0e710e650e700e7b0e840ea40ec20e;
    decBuf[2144] = 256'hd50efb0e150f230f380f440f470f510f4e0f3b0f390f260f090ffd0ee50ec90e;
    decBuf[2145] = 256'hbd0eac0e960e8d0e7b0e650e4c0e250ef70dbf0d6c0d1f0dc50c700c0d0cca0b;
    decBuf[2146] = 256'h5d0b140bd10a640a1a0aa1093009ab082e087b07d50612065b05b5041e046d03;
    decBuf[2147] = 256'hf6025f02ae013801a000f0ff1aff8afe9ffdc2fcf8fb0dfb6ffa6cf9bef820f8;
    decBuf[2148] = 256'h57f7a0f6f9f562f5b1f40bf449f392f2bcf12cf175f0cfef0cef8aee13eea7ed;
    decBuf[2149] = 256'h45edebec7aec30ecd2eb7deb30ebeaea98ea61ea2fea02eaf9e9f2e9ebe9fee9;
    decBuf[2150] = 256'h1aea29ea53ea7aea9eead1ea0feb49eb8cebf1eb4eecbbec23ed9bed0deeafee;
    decBuf[2151] = 256'h1befa4ef45f0b1f03bf1dcf148f2f8f29ff30bf494f435f5ccf556f6d3f645f7;
    decBuf[2152] = 256'hc9f747f8b8f83df9baf92cfab1fa2efba0fb07fc64fcb9fc06fd4cfd7afdb4fd;
    decBuf[2153] = 256'he8fd18fe5dfe8bfec4fef9fe29ff3cff58ff72ff76ff72ff76ff6bff68ff71ff;
    decBuf[2154] = 256'h79ff85ff98ffa5ffb1ffbbffadff9eff86ff64ff43ff26ff0bff00ff03ff06ff;
    decBuf[2155] = 256'h18ff33ff3dff40ff43ff2bff0fffecfec3fe90fe6efe5bfe4afe4ffe54fe50fe;
    decBuf[2156] = 256'h5bfe51fe3bfe1bfedcfd9cfd51fd0bfdb9fc82fc3cfcfcfbe4fbaffb71fb48fb;
    decBuf[2157] = 256'hf6fa93fa35fab0f932f9c1f83cf8bff74df7c8f64bf6faf575f5d4f468f4b8f3;
    decBuf[2158] = 256'h11f37af2a2f1d9f056f080eff1ee3aee94edd1ec4eeca8ebe5ea63ea8de9c4e8;
    decBuf[2159] = 256'h41e89be704e77ae6d9e542e5b9e43be4a9e347e3a6e23ae2d8e15be1e9e09fe0;
    decBuf[2160] = 256'h5ce020e0ffdfcddf9fdfa7df91df8adf9ddf97dfa7dfd9dfeedf26e088e0cbe0;
    decBuf[2161] = 256'h38e19fe117e289e22be398e321e4c2e459e5e3e583e61be7cbe772e834e9ebe9;
    decBuf[2162] = 256'hc1ea8aeb41ec17eda7ed5dee33efc3ef46f0ecf083f134f2daf271f322f4c8f4;
    decBuf[2163] = 256'h34f5bef53bf68cf6d6f619f73df774f7a6f7c2f7ebf72ef84af862f888f88ff8;
    decBuf[2164] = 256'h7cf876f834f8f4f7cbf778f741f70ff7e2f6b8f693f670f645f61df6d0f583f5;
    decBuf[2165] = 256'h3df5d9f496f441f4f4f3c2f3a7f38ef387f38ef37bf375f370f359f344f338f3;
    decBuf[2166] = 256'h20f316f325f337f35bf39df3ddf317f469f4a0f4d2f412f53bf561f59ff5c8f5;
    decBuf[2167] = 256'hfdf556f693f6f6f653f7a8f7f5f73bf869f892f8b7f8b1f8b7f8d3f8c4f8c8f8;
    decBuf[2168] = 256'he6f8e2f8edf802f9eef8dcf8c7f89bf83ef8fbf78ef709f7b0f63ef6d7f579f5;
    decBuf[2169] = 256'h0cf5a5f447f4daf355f3d8f246f295f11ef15cf0a5efffee67eedeed3dedd1ec;
    decBuf[2170] = 256'h47eceeeb5cebfaea7dea0beaa4e946e9c1e867e816e8cce789e765e75ae750e7;
    decBuf[2171] = 256'h6be784e7aae7e7e711e845e883e8bde800e952e99fe921ea9fea31ebe1eb88ec;
    decBuf[2172] = 256'h4aed01eea7ee6aef21f0f7f0c0f177f21df3e0f3cbf4a8f571f628f7fef7c7f8;
    decBuf[2173] = 256'hb2f990fa20fbd6fb7dfc14fd9dfd3efeaafe34ffb1ff02008700e00032015e01;
    decBuf[2174] = 256'ha101ad01ce01d801bc01b4019e016e0142011a01d80098005e000c00bfff65ff;
    decBuf[2175] = 256'hf8fe90fe33feadfd30fdbefc57fcdffb6dfb06fb8dfa3cfad5f977f93bf9eef8;
    decBuf[2176] = 256'ha8f868f83ff80af8e8f7c8f7b8f7b2f7caf7e7f712f850f8abf8fff84cf9baf9;
    decBuf[2177] = 256'h22fa9afa0cfb91fb0efca0fc29fdcafd8dfe44ff1900e3009a016f023903ef03;
    decBuf[2178] = 256'h960458050f06b5064d07fd0774083709b909600acc0a550bd20b440cab0cee0c;
    decBuf[2179] = 256'h430d640d960db10dba0db20d9e0d7e0d570d290df10cad0c6d0c230cc90b740b;
    decBuf[2180] = 256'hfb0a890a220a8f0906098808d6075f07c8063e06c1054f05cb047104ff039803;
    decBuf[2181] = 256'h3b03cd02660209029b0134010c01cf00ae00b800c200da00000130015c019a01;
    decBuf[2182] = 256'hd301f90144028a02dd025603c7034c04ed0484053506db069e072008f6088609;
    decBuf[2183] = 256'h3d0ab40a760b2d0cd30c6b0d1b0ec20e840f0710ad101911a311fc116e12b712;
    decBuf[2184] = 256'hfa124f138613b813e613ff1324142b1425141414f013c61388134f13fc12af12;
    decBuf[2185] = 256'h5512e811811123119e102110af0f0d0fa10e170e760ddf0c560cd80b460bbd0a;
    decBuf[2186] = 256'h400ace094909a8086708de0785073307cc06890665062e06fc050506fd05f505;
    decBuf[2187] = 256'h0a0629063a067206b606e4062e079c07e6075e08d0083709e5098b0af70aa80b;
    decBuf[2188] = 256'h4e0c110dc80d6e0e300fe70fbd104d1138121513df1395146b153416eb16c117;
    decBuf[2189] = 256'h51180819ae191a1aa31a211b921b171c701cc21c291d871dc31d101e421e5e1e;
    decBuf[2190] = 256'h871e8e1e6c1e661e3e1e061ed11d941d491d031db11c4e1c0b1cb61b3d1bec1a;
    decBuf[2191] = 256'h671aea195819cf182e18c21711176b16ff157515f81486141f14a7135613ee12;
    decBuf[2192] = 256'h76122512db1163113211e8108a10661045102710301038103110531066106c10;
    decBuf[2193] = 256'h90109d10a210c510dc10f1102b117511bb1120129812e9125113ae13eb132214;
    decBuf[2194] = 256'h54146f1488149e14a514c514ec1406152f15571570157e157a1557152415d814;
    decBuf[2195] = 256'h7e141114aa134c13df1296121d12cc1182110a119810f60f5e0f870ebd0dd20c;
    decBuf[2196] = 256'h340c310b830ae5091c09990822088b0701078406f2056905c804300480030903;
    decBuf[2197] = 256'h7202e801b301610118010a01fe00f300fd0006010f0125013a0133015b017f01;
    decBuf[2198] = 256'h9f01df0131027e0200037d030f0499043a05d10582062807bf077008e7087e09;
    decBuf[2199] = 256'h070aa80a140bc50b6b0c030db30d590ef10ea10f4810b41016116f11a011ea11;
    decBuf[2200] = 256'h2d1251128812ce120e135813b2130714541486148f14971472142614cc137713;
    decBuf[2201] = 256'hfe12ad1246120312c6118f115d113011f61095101c108a0fd90e330e700d850c;
    decBuf[2202] = 256'he70b570ba10a2a0abe095c09020990080c088f07dc0606063d055204b403ea02;
    decBuf[2203] = 256'h3302bd017c011a01e400b3006a002700d2ff43ffb9fe19fe81fdf8fc9efc4dfc;
    decBuf[2204] = 256'h21fc14fc20fc2bfc49fc52fc4afc33fcf5fbabfb65fb01fbbefa81fa4afa40fa;
    decBuf[2205] = 256'h49fa51fa68fa7dfa83fa88fa6ffa3cfafef9b4f95af905f9b8f85ef821f8eaf7;
    decBuf[2206] = 256'hb8f78bf751f7fef6c7f659f6f2f57af5e8f45ef4bdf326f39df21ff2aef146f1;
    decBuf[2207] = 256'he9f07cf014f0b7ef62efe9ee98ee13ee96ed24ed9fec22ecb0eb49eb06ebcaea;
    decBuf[2208] = 256'h93ea89ea80ea88ea8feab2eab8eac9eae2eae7eaf4ea0feb27eb56eba2ebfceb;
    decBuf[2209] = 256'h69eceeec6bedfdedaeee25efbcef45f09ff0f0f057f1b5f13af2b7f24af3d3f3;
    decBuf[2210] = 256'h98f44ef5f5f5b7f63af7b1f71df87ff8d8f809f953f97bf9d0f91dfa77fafcfa;
    decBuf[2211] = 256'h56fba7fb0efc36fc5bfc66fc48fc1afcf1fb9efb67fb35fb08fbeffaf6faeffa;
    decBuf[2212] = 256'he9fafafad6faadfa85fa38fabff94ef9c9f84cf8daf773f715f7d8f6a1f65bf6;
    decBuf[2213] = 256'h1cf6c1f56cf509f591f4fef39cf3fbf264f202f2a8f137f10af1c8f08bf054f0;
    decBuf[2214] = 256'h22f0e2efa8ef47efe9ee94ee31eeb9ed88ed21eddeecbaec83ec65ec5cec32ec;
    decBuf[2215] = 256'h1cec15ecf6ebdaebd4ebabeb83eb74eb4aeb3aeb34eb27eb2beb46eb57eb74eb;
    decBuf[2216] = 256'haeebc6ebddeb1bec23ec2bec31ec2bec1aec1fec08ec04ec1fec2aec4cec88ec;
    decBuf[2217] = 256'ha1ecc6ec04edfcec04ed18edf9ecddecd8ecaeeca8ecb8ecaaecbfece2ece7ec;
    decBuf[2218] = 256'hfcec08edf6ecdaecbfec8aec56ec41ec15ec05ec14ec19ec47ec80eca5ece3ec;
    decBuf[2219] = 256'h0ced23ed45ed64ed5fed6eed8eeda4edd6ed22ee68eeccee44ef96ef1af074f0;
    decBuf[2220] = 256'he6f04df1c5f116f29bf218f38af30ff48cf41ef5cff575f60cf796f737f8cef8;
    decBuf[2221] = 256'h57f9d5f946faaefa26fb77fbdefb57fca8fc0ffd88fdd9fd40fe9efedafe11ff;
    decBuf[2222] = 256'h43ff5fff78ff7fff78ff72ff6cff5dff58ff54ff41ff36ff2dff0dffe7fec3fe;
    decBuf[2223] = 256'h7efe38fee6fd83fd25fdd0fc83fc29fcecfbb5fb83fb56fb2dfbf8fad6faaafa;
    decBuf[2224] = 256'h77fa55fa1dfaf7f9d5f9b6f999f98af985f981f97df981f97ef986f989f98bf9;
    decBuf[2225] = 256'h92f998f9a7f9bbf9cdf9e7f90efa31fa5bfa8efabefaf6fa2bfb4dfb85fbabfb;
    decBuf[2226] = 256'hcdfbecfb08fc18fc26fc3bfc3ffc50fc60fc69fc7bfc90fc99fca6fcb7fcb5fc;
    decBuf[2227] = 256'hb3fcadfc9ffc8dfc81fc72fc64fc5ffc5afc5efc62fc64fc67fc64fc59fc4afc;
    decBuf[2228] = 256'h38fc1efc05fcf6fbe7fbe0fbddfbe4fbeefbfafb08fc1afc26fc35fc43fc53fc;
    decBuf[2229] = 256'h62fc80fc9efcc0fcf3fc23fd5cfd9ffddffd19fe5cfe9cfec5fe09ff49ff83ff;
    decBuf[2230] = 256'hc6ff060040009200df0025018a01cc013a02a102fe025303cc031e048504e204;
    decBuf[2231] = 256'h50059905f70534068106db0617077a07bd0712087508b8080d0944098a09b709;
    decBuf[2232] = 256'he109f709190a390a550a790a990ab70ad20ae30af30aea0add0ac30a960a6a0a;
    decBuf[2233] = 256'h2c0af209af096f0935090109b5086f082f08d40780071d07bf06520608069005;
    decBuf[2234] = 256'h3e05f504970442040b04c50373033c03e2028d0256021002d001a70182015f01;
    decBuf[2235] = 256'h5901530144014901550151016a0180019a01c701f30131027b02d5022a038d03;
    decBuf[2236] = 256'heb033f048c04e6043b058805e2051f066c06c606030750079607d5070f085308;
    decBuf[2237] = 256'h8008aa08de08f30812092e093d095509590955094a093b091b09fd08d308a008;
    decBuf[2238] = 256'h70083808f407b4077b072807db0695064306e00582052e05e10487043204fb03;
    decBuf[2239] = 256'hc9039b0382035d033a0328030c03f202e402d702bc02c002c902cc02e4020603;
    decBuf[2240] = 256'h1d0354038903b903fe033e047704bb040d0544059e05f30540069a0607075107;
    decBuf[2241] = 256'hae071b088308e00835098209c8091a0a510a830ac30aec0a120b340b540b700b;
    decBuf[2242] = 256'h890ba00bb60bba0bbd0bba0bb10b9a0b7e0b5b0b310b0a0bdc0ab00a880a650a;
    decBuf[2243] = 256'h320a020ac90986094609fc08a2084d08ea078c073707ea06a40677063d06f905;
    decBuf[2244] = 256'hcc0592054f050f05c4047e043f04f403c20395036b03550340032e0311030203;
    decBuf[2245] = 256'heb02c502a102770250022c02150208020c021d022d0258028402a002ce02ed02;
    decBuf[2246] = 256'h0a0323033a0347035a0373038303a803d603020440047904ae04ec0426054b05;
    decBuf[2247] = 256'h8905b205d805fa052606420670069c06c306f1062a074f077f07ab07c707eb07;
    decBuf[2248] = 256'hf907f507f107e607d007b607a507890775076b075507470734071a07fb06d406;
    decBuf[2249] = 256'h9c0668062a06f005ca059a0562054c05370524051f0519050205f604da04b404;
    decBuf[2250] = 256'h9a047a0454044404360432043e04560466049104bd04d90407053f0556059405;
    decBuf[2251] = 256'hbd05e20520065a069e06dd0628076e07ae07f8072a0857088108a608bb08da08;
    decBuf[2252] = 256'he008ef08fd080a0915092009230926091e091709ff08dd08b30881084308f907;
    decBuf[2253] = 256'h9f074a07fd06a3063606ec058e053905ec0492043e04db036203f0026c021202;
    decBuf[2254] = 256'h80011e01c50053000900c6ff8aff53ff21fff3fecafeb3fe91fe65fe49fe2ffe;
    decBuf[2255] = 256'h18fe14fe18fe1bfe37fe5afe7bfeb2fee6fe17ff4fff83ffb3ffdfff1d005700;
    decBuf[2256] = 256'h9a00da0014016601b3010d026202af02e10221035b038f03b203c503d503ef03;
    decBuf[2257] = 256'hfd0312041e042f043f0453046004630460045a044b042f040c04e303b0038003;
    decBuf[2258] = 256'h48031303e302b7028502540229020102c901940157011d01d900990060003a00;
    decBuf[2259] = 256'h0a00ebffcfffb5ffa7ff9aff87ff7dff67ff58ff41ff31ff23ff1bff1dff28ff;
    decBuf[2260] = 256'h36ff4dff69ff8cffa3ffc9ffe3fffaff06001a002b0041005b0074009c00c400;
    decBuf[2261] = 256'hf2002a015e019c01d601fc012c024b026702810298029c02a802ab02b502b702;
    decBuf[2262] = 256'hba02bc02c302c102bc02b302a3028c027602500222020302d001a00168013301;
    decBuf[2263] = 256'h0301cb00880048000e00bbff6eff14ffa7fe40fee2fd8efd2bfdcdfc78fc15fc;
    decBuf[2264] = 256'hb7fb63fb00fba2fa4dfaeaf9a7f93af9f0f893f856f809f8c3f795f75cf736f7;
    decBuf[2265] = 256'h22f7f6f6daf6caf6b3f6a6f69bf690f68df68af692f69ef6adf6bff6d9f6f2f6;
    decBuf[2266] = 256'h0ef738f760f798f7cdf70af855f89bf8dbf825f96bf9abf9e4f928fa56fa8ffa;
    decBuf[2267] = 256'hd3fa00fb3afb6ffb91fbbdfbe4fbfefb27fc44fc5dfc74fc92fc96fc99fca9fc;
    decBuf[2268] = 256'ha0fc99fc8dfc6dfc4cfc26fceefbb9fb89fb51fb1cfbecfab4fa80fa4ffa17fa;
    decBuf[2269] = 256'he3f9b3f96ef92ef9f4f8a2f855f823f8d1f79af768f728f7fef6d9f6a9f67df6;
    decBuf[2270] = 256'h6cf648f631f624f619f61cf61ff622f62ff645f64df660f67ff68bf6a7f6cdf6;
    decBuf[2271] = 256'he7f610f743f765f79ef7d2f710f84af87ef8aef8e7f82af958f981f9b5f9d8f9;
    decBuf[2272] = 256'hf7f92afa3efa51fa6dfa72fa80fa8dfa89fa8dfa96fa93fa96fa98fa89fa7bfa;
    decBuf[2273] = 256'h76fa5efa37fa1dfaebf9baf98ff951f907f9d5f895f84af818f8c6f779f747f7;
    decBuf[2274] = 256'h07f7bdf68bf64bf612f6ecf5bcf590f569f530f5fcf4ccf487f459f420f4ebf3;
    decBuf[2275] = 256'hc9f3b6f3a5f3a0f3a5f3b1f3c5f3ddf3edf301f413f416f420f42ef434f442f4;
    decBuf[2276] = 256'h58f46cf48ff4b8f4e0f418f54cf57df5b5f5f8f526f660f6a3f6d1f60bf74ef7;
    decBuf[2277] = 256'h8ef7c8f7fcf72cf858f88bf89ff8cbf8e7f8f7f80ef934f943f964f992f9a5f9;
    decBuf[2278] = 256'hcdf9fbf91afa41fa65fa7cfa89fa9cfa92fa95fa98fa80fa77fa74fa67fa69fa;
    decBuf[2279] = 256'h70fa72fa81fa99faa2fab1fabefabbfab9fab7faa0fa91fa82fa66fa52fa4ffa;
    decBuf[2280] = 256'h3ffa3cfa3ffa3cfa43fa4dfa4bfa50fa5dfa63fa75fa8afa9efabbfadefafefa;
    decBuf[2281] = 256'h1cfb37fb49fb5efb6dfb6ffb77fb79fb7ffb8bfba3fbc3fbf2fb2afc5efcaafc;
    decBuf[2282] = 256'hf0fc30fd6afdadfdc8fdf2fd17fe2cfe3ffe44fe54fe61fe7ffe93feabfed4fe;
    decBuf[2283] = 256'hfbfe1fff49ff70ff8affa1ffb6ffc2ffc5ffbcffb3ffa6ff91ff7cff6aff55ff;
    decBuf[2284] = 256'h41ff33ff1eff0afff8fee7fed8fec6feb5fea7fe99fe8cfe84fe7afe70fe65fe;
    decBuf[2285] = 256'h51fe3ffe2efe13fef8fdd8fdc3fdaffda5fda2fdb0fdcdfdf0fd1afe4cfe8afe;
    decBuf[2286] = 256'hb3fef7fe24ff3dff63ff85ff98ffb4ffceffeeff140042007b00be0010015d01;
    decBuf[2287] = 256'hb7010c025902b302f0023d038303c303fc03220452047e04a504c904e904ff04;
    decBuf[2288] = 256'h1a052b0541055505680582059a05b605d905fa0517063a065106670672066806;
    decBuf[2289] = 256'h58063e061806f405c1059105720555053c0537053b053f0558056e0576058905;
    decBuf[2290] = 256'h8b05800576056705470530051a05ff04f504f204ef040605230536055c058b05;
    decBuf[2291] = 256'haa05d105f50515063c0660066d068b06a606b806d406e706f20608071c072907;
    decBuf[2292] = 256'h43075c0771079d07c807f00728085d088d08d108ff0828094e09620969096e09;
    decBuf[2293] = 256'h690952093d0922090909fa08f108ee08fa080d0920093f095409670979098809;
    decBuf[2294] = 256'h80097d09710951093a091409e608c708aa087c085d0841082708190815080208;
    decBuf[2295] = 256'h050808080608130810080a080c080308eb07e007ca07a50796077f0769076507;
    decBuf[2296] = 256'h69076c078607a507c307f607260851088408b408d308060928092f0956096509;
    decBuf[2297] = 256'h73098909a409b509e409140a400a890acf0a0f0b6a0bbf0bf60b3c0c7b0ca50c;
    decBuf[2298] = 256'hd90cee0c010d110d210d1c0d200d2c0d220d310d3a0d3c0d4d0d5c0d620d750d;
    decBuf[2299] = 256'h820d850d8f0d890d730d630d430d0c0de70ca90c5e0c180cd90b7e0b410b0a0b;
    decBuf[2300] = 256'hc40aa90a800a4b0a360a240afc09e309cc09a5098c096b0934090f09de08a608;
    decBuf[2301] = 256'h8108510818080208ed07ce07d407d907dd070408270848087708a208b308d708;
    decBuf[2302] = 256'hee08f20806091009130928093a094b096a099d09cd09060a3a0a6a0aa30ad70a;
    decBuf[2303] = 256'h070b330b4f0b5e0b760b7a0b6e0b6b0b550b350b200b050be50ad90abd0aac0a;
    decBuf[2304] = 256'ha90a9a0a8d0a8b0a800a6a0a560a2f0afc09cc0987094709fd08a3084e080108;
    decBuf[2305] = 256'ha70752070507bf06800646062006f005dd05c105a8059a058505690551053505;
    decBuf[2306] = 256'h0205e004b40482045f0440042404150419041d043104490465049004b704d104;
    decBuf[2307] = 256'hfb0422053c055c057a058d05ad05c205d505ee05fd0512062906450660068e06;
    decBuf[2308] = 256'hba06e10619074e0770079c07b807c807d507d107b607a5078207590731070307;
    decBuf[2309] = 256'hd706bb0697068006620647062f061906f905d305af057c053e05f4049a044504;
    decBuf[2310] = 256'he2036a03f80291021902c70160010201c6008f0049000900cfff8cff4cff12ff;
    decBuf[2311] = 256'hc0fe73fe2dfedafd8dfd47fd08fdbdfc8bfc4bfc12fcecfbbcfb9dfb8cfb7dfb;
    decBuf[2312] = 256'h78fb7cfb80fb99fba8fbbcfbc9fbd5fbdcfbe2fbdcfbd8fbd9fbdafbdefbeffb;
    decBuf[2313] = 256'h04fc1efc45fc73fc9ffcd1fcf4fc2cfd51fd66fd85fd96fda6fdaafdaefda3fd;
    decBuf[2314] = 256'h91fd88fd74fd61fd56fd42fd35fd2efd1ffd11fd09fdf3fcdafcbafc8bfc60fc;
    decBuf[2315] = 256'h22fcd7fb7dfb41fbdefa80fa2bfab2f961f9faf89cf847f810f8caf778f757f7;
    decBuf[2316] = 256'h11f7e4f6baf686f648f60ef6bcf56ff515f5c0f45df41af4c5f38ef35cf32ef3;
    decBuf[2317] = 256'h26f31ff326f32cf33df34cf351f366f362f36df37cf37ff387f3a1f3acf3c1f3;
    decBuf[2318] = 256'hedf3fff31bf43ff456f474f4a7f4bbf4e7f41af53cf55bf58ef5a2f5c2f5e9f5;
    decBuf[2319] = 256'heef5eaf5f6f5e3f5d1f5cef5aff599f596f576f561f55df544f535f532f515f5;
    decBuf[2320] = 256'hfaf4e8f4baf47cf452f400f4b3f359f304f3a1f243f2eff18cf149f10cf1d5f0;
    decBuf[2321] = 256'ha3f075f03cf025f0e7efaeef79ef3beff1eebfee7fee35ee17eed7ed9ded78ed;
    decBuf[2322] = 256'h48ed1ced00eddcecbbecb7eca4ec99eca9ecacecbeece2ecf1ecffec1ded21ed;
    decBuf[2323] = 256'h2bed41ed38ed3bed50ed53ed66ed89edadedd7ed20ee52ee92eeccee00ef30ef;
    decBuf[2324] = 256'h68ef8eefb0efdcefe2eff1ef1bf02cf03bf06ef082f0a2f0d4f0f7f016f154f1;
    decBuf[2325] = 256'h6df183f1b3f1b9f1bff1d9f1cbf1c7f1caf1c0f1c3f1ccf1bff1c1f1d0f1c6f1;
    decBuf[2326] = 256'hc1f1c5f1b2f1a0f19df186f176f17ff172f16ff17af16cf167f165f14ff12cf1;
    decBuf[2327] = 256'h15f1e6f0bbf09ef07bf06df071f06df07ff0a7f0c3f0ddf007f123f132f149f1;
    decBuf[2328] = 256'h3cf140f144f141f144f151f158f16ff19ef1c0f1e0f11ef247f27bf2b9f2e2f2;
    decBuf[2329] = 256'h17f355f37ef3b3f3e3f302f435f465f484f4b7f4e7f412f545f575f594f5c7f5;
    decBuf[2330] = 256'h05f61ef652f682f6aef6d5f60ef724f747f77ff795f7aaf7bdf7c2f7c8f7ccf7;
    decBuf[2331] = 256'hbff7c3f7d5f7d8f7ecf70ef825f854f88cf8a3f8c5f8e4f8eaf8eff8f4f8dff8;
    decBuf[2332] = 256'hd3f8c8f8b9f8b6f8bef8c5f8d4f8eef8fff81bf937f948f964f97ff998f9b4f9;
    decBuf[2333] = 256'hcff9eff90cfa37fa53fa77fa97faadfacffae7fafcfa1ffb3ffb65fb93fbbffb;
    decBuf[2334] = 256'hf2fb30fc69fc9efcdcfc16fd4afd7afdb2fdd8fd08fe34fe50fe7efeaafec6fe;
    decBuf[2335] = 256'hf4fe20ff52ff90ffcaff0e006000ad00f30033016c01a101c301e201ff010e02;
    decBuf[2336] = 256'h1c0231024c026c029202c002ec022a0363038903b903f1031704390458047504;
    decBuf[2337] = 256'h8e04a504b204cd04df04e204f004f804fa04050513051f0538055e057805a105;
    decBuf[2338] = 256'hd405e9051406310640064e065b064f0652064f064c064f0656065d0673068c06;
    decBuf[2339] = 256'h9e06c006ea0606072a07540770079e07ca07da07fe0715082208360840083d08;
    decBuf[2340] = 256'h5108630874089408be08e5081d0952097409ac09e109030a3c0a610a830aaf0a;
    decBuf[2341] = 256'hcb0ae50a050b230b2f0b4e0b630b670b800b9c0baf0bd60b040c300c6e0ca70c;
    decBuf[2342] = 256'hcd0cfd0c290d450d540d590d4c0d480d370d1b0d170d1a0d110d250d370d3e0d;
    decBuf[2343] = 256'h5e0d880d990dbd0dd40de10d030e1b0e1f0e3a0e440e3b0e3e0e360e1c0e180e;
    decBuf[2344] = 256'h0f0efb0d030e130e160e340e6b0e810ebf0ef90e0f0f400f6b0f7c0f960fa40f;
    decBuf[2345] = 256'h9f0fb30fc40fc10fdb0ff40ffd0f221046105d108c10c410db10191142116711;
    decBuf[2346] = 256'h8a11a911af11be11cc11b711bb11b711a111a411a711a011b311c011b911d011;
    decBuf[2347] = 256'hd911d111d911d611bf11c211ae11911185116d1144112811fa10c2108d105d10;
    decBuf[2348] = 256'h0c10eb0fb90f790f710f5a0f460f4c0f520f420f470f320f070feb0ebd0e840e;
    decBuf[2349] = 256'h500e200ee80dc20da00d800d7b0d760d680d750d800d7d0d990da40da80db80d;
    decBuf[2350] = 256'hc00db30dbf0db40d9a0d970d870d6d0d6a0d670d580d6b0d800d890db00dd70d;
    decBuf[2351] = 256'he70d070e1c0e200e320e350e210e190e040ee40dd70dbc0d960d860d660d400d;
    decBuf[2352] = 256'h3a0d2d0d170d1b0d180d0e0d170d1a0d040d010de40cb20c900c570c050cce0b;
    decBuf[2353] = 256'h880b480b1f0bf90ac90ab60ab10a970a930a860a720a680a5f0a3f0a320a170a;
    decBuf[2354] = 256'hf109d709b709900977094d0926090c09ec08ce08c208b808b508c908d608e208;
    decBuf[2355] = 256'h020922092f094a0954095809600953093e09350923090d09ff08ed08d708d408;
    decBuf[2356] = 256'hd708d508e808fa080b092609410953095c095f094d0937091209da08a5086708;
    decBuf[2357] = 256'h2e080808d807ac07900776075f075b07480728070a07e006ad066f063606e305;
    decBuf[2358] = 256'h96055005ec04a90454040704c1036f032203f002b002760251022102f501cd01;
    decBuf[2359] = 256'haa01800159012a01f200be00800036000400c4ff8aff64ff34ff09fff8fedefe;
    decBuf[2360] = 256'hd9fedefee2feecfe02ff10ff23ff38ff46ff4eff55ff53ff4dff45ff39ff32ff;
    decBuf[2361] = 256'h30ff34ff3cff4bff62ff85ffa5ffc3ffdefff6ff060014001700190013000500;
    decBuf[2362] = 256'hf5ffe6ffd4ffbaffa9ff8dff72ff59ff3dff22ff09ffe7fec7febafe9ffe7ffe;
    decBuf[2363] = 256'h6afe3ffe18feeafdb2fd6efd2efde4fc9efc5efc14fccefba0fb77fb51fb3dfb;
    decBuf[2364] = 256'h2afb24fb15fb10fb04fbf0fadffabcfa9cfa76fa48fa1cfa00fadcf9cef9c1f9;
    decBuf[2365] = 256'hc5f9d0f9e6f9fff926fa54fa73fa9bfab4fad5faeafaf6fa00fb09fb0cfb14fb;
    decBuf[2366] = 256'h25fb2bfb31fb48fb51fb60fb77fb81fb89fba1fba4fbb2fbc5fbc7fbc9fbd3fb;
    decBuf[2367] = 256'hcbfbbcfbb2fb98fb65fb43fb0bfbc7fa9afa4ffa1dfaf0f9b6f990f96ef942f9;
    decBuf[2368] = 256'h1bf901f9cef89ef873f829f8e3f7a4f749f7f4f6a7f64df6f8f5c1f57bf54df5;
    decBuf[2369] = 256'h24f5f0f4cdf4bbf49ef485f46ef450f435f41cf4faf3e3f3c5f3a2f382f36df3;
    decBuf[2370] = 256'h51f340f33df334f337f347f352f36cf393f3b6f3e0f313f443f47bf4b0f4d2f4;
    decBuf[2371] = 256'hf1f419f51ef52cf549f545f550f566f574f58cf5b4f5d1f5fff543f671f69af6;
    decBuf[2372] = 256'hdef6f9f622f739f740f746f74cf732f71bf717f7fcf6e3f6daf6c6f6b8f6bbf6;
    decBuf[2373] = 256'hacf6a2f69df684f66cf65cf631f612f6eaf5bcf584f55ff52ef503f5e7f4aef4;
    decBuf[2374] = 256'h7af465f42df407f4e5f3c6f39ef38ff378f363f35ff34df344f347f334f328f3;
    decBuf[2375] = 256'h26f314f308f302f3f4f2f2f2faf2fff214f333f351f383f3c1f3eaf31ff45df4;
    decBuf[2376] = 256'h97f4cbf4fbf41af542f570f58ff5abf5cff5f0f50df640f662f68ef6c0f6f1f6;
    decBuf[2377] = 256'h1cf75af783f7a9f7d9f7ecf7fdf716f812f816f81af808f8f9f7f0f7d8f7c3f7;
    decBuf[2378] = 256'hbaf79df78af77ff75df746f739f70ef7f2f6d9f6aff67cf65af62ef6f0f5c7f5;
    decBuf[2379] = 256'h84f544f51af5d7f4a9f480f45bf438f425f409f4faf3f5f3e0f3d4f3caf3b4f3;
    decBuf[2380] = 256'ha0f393f374f35ff353f349f345f34ef351f36bf391f3abf3d5f312f43cf470f4;
    decBuf[2381] = 256'haef4d7f40cf54af573f598f5c9f5e8f50ff63df669f690f6c9f6fdf62df772f7;
    decBuf[2382] = 256'hb2f7ecf72ff86ff8a9f8ecf81af954f988f9abf9caf9fdf911fa24fa35fa3afa;
    decBuf[2383] = 256'h48fa4cfa48fa4cfa55fa52fa5ffa70fa7bfa8dfaa2faa5fab2fabefaaffa9dfa;
    decBuf[2384] = 256'h8cfa6cfa43fa27faf9f9cdf9b1f98df976f971f966f95bf958f950f94df94bf9;
    decBuf[2385] = 256'h3cf932f925f90df9fcf8e6f8ccf8b3f8aaf896f889f88bf88df89bf8aef8c6f8;
    decBuf[2386] = 256'he8f812f92ef95cf988f9a4f9c8f9f2f903fa26fa47fa5cfa77fa97fab4fad7fa;
    decBuf[2387] = 256'h01fb28fb56fb8ffbc3fb01fc3bfc7efcbefc08fd3afd7afdb4fddafdfcfd1bfe;
    decBuf[2388] = 256'h2cfe3bfe49fe56fe5afe6bfe7bfe89fea6febafed2feeefe02ff1aff2aff2dff;
    decBuf[2389] = 256'h2aff28ff19ff03ffeffed2feb7fe97fe79fe5efe46fe2afe0ffefdfde7fdd3fd;
    decBuf[2390] = 256'hc6fdb1fd9cfd8ffd7afd66fd4efd32fd17fdfefce2fccffcb6fca7fc9efc91fc;
    decBuf[2391] = 256'h8ffc95fc97fcaafcc2fcd8fcf7fc15fd38fd58fd7ffd98fdb9fdd6fdeafdfbfd;
    decBuf[2392] = 256'h0bfe1ffe37fe59fe79feb1fee5fe23ff6dffb3ff050052009800d80012013801;
    decBuf[2393] = 256'h5a0179018a01a401b201c701e201fa011d023d025b028602ad02d102f1020f03;
    decBuf[2394] = 256'h2a0343035203610368036b0364035e03520340032b031703ff02e902d502c802;
    decBuf[2395] = 256'hc102b202b402b902bb02bf02c602c502c602bf02b202a00286026d0251023e02;
    decBuf[2396] = 256'h1e0212020602fc0105020e0220023f025d0278029702b502c802e102f002f302;
    decBuf[2397] = 256'h0003030301030b031703220339035b037c03a203d003fc032e046c049504ca04;
    decBuf[2398] = 256'hfa0426054d0571059105af05c305cd05dd05eb05f305ff0512061f0639065906;
    decBuf[2399] = 256'h7606a906cb06f7062a074c076b078707a107a607aa07a6078d07840770075807;
    decBuf[2400] = 256'h4907400733073a073c073e0751075f076a0779078307820786077c0767075f07;
    decBuf[2401] = 256'h470725070e07f806dd06cc06c206b406b706b906bb06c906d206d306e406f306;
    decBuf[2402] = 256'hf106f606fb06f906fe06fa06ed06f206f406ed06f80600070407170733074707;
    decBuf[2403] = 256'h6d079107b207d807060819084008640869088608920895089f08a708aa08bb08;
    decBuf[2404] = 256'hce08db08ff082209430969098d09ad09d409f709050a230a2f0a2b0a350a320a;
    decBuf[2405] = 256'h250a270a210a170a180a170a0f0a1e0a280a2e0a430a510a590a6e0a770a740a;
    decBuf[2406] = 256'h7b0a790a670a600a510a370a2d0a170a030afb09f409e509ef09f409f309030a;
    decBuf[2407] = 256'h120a140a240a2e0a2c0a3c0a3e0a300a350a310a230a250a1d0a0c0a130a190a;
    decBuf[2408] = 256'h130a220a340a3b0a570a6a0a7c0a980aa30aa70abd0ac00ab80abf0abd0ab30a;
    decBuf[2409] = 256'hb40ab30aab0aba0ac40aca0ae20a020b0e0b390b550b640b850b9a0ba60bb70b;
    decBuf[2410] = 256'hc10bb80bc00bb90bae0bb00bb20ba60bb70bc60bcc0be30bff0b0a0c2a0c480c;
    decBuf[2411] = 256'h530c730c880c8c0ca40ca70c9f0cac0caa0c960c940c880c750c6d0c610c4a0c;
    decBuf[2412] = 256'h4d0c4a0c420c4e0c500c4a0c5a0c5c0c4e0c500c410c230c0e0cf30bbe0ba80b;
    decBuf[2413] = 256'h850b4d0b370b220bf60af10ae10aca0ac60aba0a9b0a960a830a5d0a4d0a360a;
    decBuf[2414] = 256'h070ae809cc09a80991097c0959094b093e092b092e092b092309300932093009;
    decBuf[2415] = 256'h420944093e0948094a0942094c094b093f09440945093f094509480949095609;
    decBuf[2416] = 256'h64096c098509a409b109d409eb09f8090b0a160a130a150a0e0af809f009dd09;
    decBuf[2417] = 256'hc309b909af09a109a309a6099f09a909a40996099409840964094d092f090409;
    decBuf[2418] = 256'he808ba0882085c082c080108d907ab077f0763073507fd06e606b6068a066e06;
    decBuf[2419] = 256'h40062106fa05d605ac059005620536050f05e104b5048d046a0440042f041504;
    decBuf[2420] = 256'hfe03f203e603db03df03dc03d403d603d003be03b703ac039e03950390038c03;
    decBuf[2421] = 256'h90039903a503ba03d403ed0309041c042e0444045204550460045a0458045a04;
    decBuf[2422] = 256'h55044d044f044b0441043d0434042804230415040604fb03e903d803c103ab03;
    decBuf[2423] = 256'h9103790350032903fb02c2027f023f02f501af016f012501df009f0054000e00;
    decBuf[2424] = 256'he1ffa7ff64ff36ffecfebafe68fe31fed7fd9afd4dfd07fdb5fc68fc22fcf4fb;
    decBuf[2425] = 256'hbafb86fb56fb2afb0efbeafacafaacfa91fa78fa5cfa49fa30fa1afa06faf4f9;
    decBuf[2426] = 256'he8f9e2f9dcf9ddf9dff9e1f9eaf9f5f906fa19fa2bfa3cfa5cfa73fa80fa9bfa;
    decBuf[2427] = 256'hacfabcfad0fad8fadffaeafaecfae7faebfae4fae3fae9fae5fae4faecfaebfa;
    decBuf[2428] = 256'he8faedfadffad1fac9fab0fa8afa70fa3dfa0dfae1f9a4f96af944f906f9cdf8;
    decBuf[2429] = 256'ha7f869f830f80af8daf7a2f77cf73ef705f7dff6a1f667f633f6f5f5abf579f5;
    decBuf[2430] = 256'h39f5fff4daf49cf473f44df41df4fef3edf3d3f3bcf3b8f3a4f39af39df394f3;
    decBuf[2431] = 256'h8df398f38ef38cf398f393f395f3a9f3acf3b4f3d3f3e0f3fbf321f445f466f4;
    decBuf[2432] = 256'h94f4b4f4d0f4fef411f52df546f554f569f585f588f598f5acf5b4f5c4f5e0f5;
    decBuf[2433] = 256'he4f5f5f50bf608f610f621f616f60cf611f6f9f5daf5c4f5a1f578f55cf523f5;
    decBuf[2434] = 256'heff4daf4a2f46df44bf413f4edf3cbf39ff36df34af31ef3ecf2c9f291f25df2;
    decBuf[2435] = 256'h2df2f4f1c0f190f157f123f1f3f0c7f094f080f054f038f033f01cf00ff013f0;
    decBuf[2436] = 256'h08f0ffef08f005f007f012f010f015f024f026f036f051f05df075f09ef0baf0;
    decBuf[2437] = 256'hdef01af143f169f1a7f1d0f1f5f133f25df282f2b2f2d1f2f9f227f33af361f3;
    decBuf[2438] = 256'h99f3b0f3d2f30bf421f443f47cf492f4a7f4dff4e7f4fbf41af520f525f53cf5;
    decBuf[2439] = 256'h38f534f538f528f525f523f50df505f507f5f2f4e9f4ecf4e0f4d5f4d7f4c8f4;
    decBuf[2440] = 256'hc1f4bff4a8f493f48af46df45af44ff433f420f415f4fff3fcf304f4fdf308f4;
    decBuf[2441] = 256'h1ef421f433f44df45ff475f48ef4a0f4b6f4d5f4ebf406f52cf546f570f597f5;
    decBuf[2442] = 256'hbbf5eef51ef64af687f6c1f6f6f634f76df7a2f7edf733f861f89bf8def80cf9;
    decBuf[2443] = 256'h46f97af9aaf9d6f914fa3dfa63faa1facafaeffa1ffb4bfb73fb96fbb7fbd5fb;
    decBuf[2444] = 256'hf7fb05fc12fc25fc29fc2cfc35fc32fc39fc40fc3efc3ffc44fc43fc47fc50fc;
    decBuf[2445] = 256'h4cfc4bfc4afc42fc3dfc34fc26fc1dfc12fcfefbf7fbebfbdcfbd2fbcdfbc8fb;
    decBuf[2446] = 256'hc9fbcdfbd1fbdbfbedfbf9fb10fc26fc35fc51fc6dfc85fc9bfcb5fccdfce9fc;
    decBuf[2447] = 256'h05fd24fd42fd65fd85fdb4fde0fd07fe3ffe74fea4fedcfe11ff41ff79ffaeff;
    decBuf[2448] = 256'hdeff090031005f008b00b200d600000127014b017e01a001cc01f30121024102;
    decBuf[2449] = 256'h68028c02ac02ca02dd02f6020c031a032c033d0348035603650370037a038603;
    decBuf[2450] = 256'h8e039903a803b203be03cd03db03e403ef03f703fd030604030406040c040804;
    decBuf[2451] = 256'h07040d040f041604210429043d0454046404780490049f04b904cb04da04ee04;
    decBuf[2452] = 256'h010508051f052f053d05550571057d059505b705cf05ec050f0626064d067006;
    decBuf[2453] = 256'h9106b706db06f20618073c07530771078c079e07b407c807d507ea07fe070608;
    decBuf[2454] = 256'h2008320841085b086d087c089108a308aa08b908c308c108cd08ce08c708d008;
    decBuf[2455] = 256'hd308cc08d408d808d108d508d408c908ca08c608b408ad08a208900889087a08;
    decBuf[2456] = 256'h6c0867085c084e0849084108330835082d082208260820081608220824081d08;
    decBuf[2457] = 256'h2c0836083708460850084b0859085f085e0866086d0869087708800881089508;
    decBuf[2458] = 256'ha208ae08c508db08e408fb080b0914092609320938094a095b095d096f097b09;
    decBuf[2459] = 256'h7d098f099b099909a309a8099d09a409a009920994098f097f097c0976096709;
    decBuf[2460] = 256'h65095f094f0948093e0928091e091609fe08ee08e008c808bf08b6089f089c08;
    decBuf[2461] = 256'h8d087b086f0864084e0846083308230818080a08f707f407e807de07e007db07;
    decBuf[2462] = 256'hcf07d407d007c407c907c507b707c007be07b707c307c807c607d507df07de07;
    decBuf[2463] = 256'hf007f707f907070809080708110810080708110813080f08150814080e081208;
    decBuf[2464] = 256'h0e080008fe07f607e707e107d507c307c107b207a0079d07930781077a076607;
    decBuf[2465] = 256'h4f07450737071a07ff06e706ca06af0697066e06520638060f06f305cf05a505;
    decBuf[2466] = 256'h89056505450527050c05e504cc04b50497048b0473045d044f043c042c041d04;
    decBuf[2467] = 256'h0b04f503e703da03c403bc03a90399038e03840374037203680360035e035903;
    decBuf[2468] = 256'h5303560353035003560359035a03610367036c037703800384038b038f039203;
    decBuf[2469] = 256'h9b039f03a003a503a2039c039b0395038a037e03710361034e033c0322031003;
    decBuf[2470] = 256'hf402d902c702b102980286026a024f0236021a02ff01e001c2019f017f015001;
    decBuf[2471] = 256'h2401fd00cf00a3007b004d002200faffccffa0ff79ff55ff2bff04ffe0fec0fe;
    decBuf[2472] = 256'ha2fe7ffe68fe4afe2ffe17fe07feedfddcfdccfdbefdb6fdaffda4fda6fda8fd;
    decBuf[2473] = 256'ha6fdabfdb4fdbbfdc2fdc9fdd0fdd7fde2fde6fde9fdeffdf4fdfcfd04fe0ffe;
    decBuf[2474] = 256'h1cfe25fe30fe41fe4cfe56fe65fe70fe7afe8afe90fe92fe9bfe9cfe9bfe9cfe;
    decBuf[2475] = 256'h96fe8efe87fe7afe64fe56fe39fe1efe05fee9fdc6fdaffd89fd65fd4efd28fd;
    decBuf[2476] = 256'hf9fcdafcb3fc8ffc65fc3efc10fce4fbbdfb8ffb6ffb48fb1afb07fbe0fac6fa;
    decBuf[2477] = 256'haffa91fa7efa65fa43fa2cfa0efaebf9d4f9bff9a4f992f983f96ef967f964f9;
    decBuf[2478] = 256'h62f960f969f971f97bf98bf995f9a8f9bff9d5f9eff90ffa24fa3ffa5ffa74fa;
    decBuf[2479] = 256'h8ffaaefabbfad6faeffaf8fa0cfb1ffb2ffb3efb54fb5dfb6ffb85fb87fb95fb;
    decBuf[2480] = 256'ha5fba7fbadfbb3fbaefbacfbb0fba8fba2fba5fb9afb8efb90fb81fb6ffb63fb;
    decBuf[2481] = 256'h4bfb2ffb1cfbf5fac7faa8fa81fa52fa27fafff9c7f9a1f971f946f91ef9f0f8;
    decBuf[2482] = 256'hc4f8a8f87af85bf83ff81bf8faf7eef7d3f7c1f7b1f79df78bf77ff76cf75af7;
    decBuf[2483] = 256'h4ef73bf72df726f71cf716f717f719f721f72df738f74cf763f773f787f7a4f7;
    decBuf[2484] = 256'hb7f7d0f7f2f709f827f852f879f89df8d0f8f2f82bf95ff981f9adf9e0f902fa;
    decBuf[2485] = 256'h21fa49fa6dfa84faa2fabdfad5faebfaf9fa0cfb1cfb27fb31fb3dfb3ffb43fb;
    decBuf[2486] = 256'h4afb47fb48fb4dfb45fb3ffb40fb37fb30fb29fb19fb08fbf9fadffac7fab1fa;
    decBuf[2487] = 256'h91fa73fa58fa39fa1bfa00fae0f9c3f9aff990f97af967f94ff939f92af918f9;
    decBuf[2488] = 256'h0cf90af900f9fef803f908f911f921f930f94af963f97ff99af9baf9d7f9faf9;
    decBuf[2489] = 256'h1bfa41fa65fa8efaaafacefaf8fa1ffb43fb6dfb94fbc2fbeefb15fc44fc7cfc;
    decBuf[2490] = 256'ha1fcd1fc0afd3efd6efda7fdccfdfcfd28fe44fe72fe91feaefebdfeddfeeafe;
    decBuf[2491] = 256'hf6fe00ff0aff0cff0fff0dff0bff05fff5feeafedcfec9feb7fea6fe8ffe79fe;
    decBuf[2492] = 256'h65fe52fe42fe2efe1cfe10fe01feeffddffdd4fdc2fdb1fd9efd8cfd80fd69fd;
    decBuf[2493] = 256'h53fd44fd32fd1dfd0efd01fdf5fcebfce1fcd8fcdafcd8fcdcfce5fceffcfefc;
    decBuf[2494] = 256'h14fd28fd45fd60fd80fd9efdc0fde1fd07fe2bfe4bfe72fe95febffedbfe09ff;
    decBuf[2495] = 256'h29ff45ff73ff92ffb9ffddfffeff1b00460062008600b000cc00f00010013601;
    decBuf[2496] = 256'h500170018e01b101d101ef011202320250026b0284029a02ae02bb02c702cd02;
    decBuf[2497] = 256'hd702d502d402d502ce02c802c202bb02b502af02ab02aa02a702a502a4029f02;
    decBuf[2498] = 256'h9d029f02a0029f02a402a602a602ad02b302b602be02c402c502cc02d202d302;
    decBuf[2499] = 256'hdd02e602e502ed02f802fc020603110319032b033b0346035c03700382039d03;
    decBuf[2500] = 256'hbc03d103f40315043204550476049304b604d704f4040f05280538054c055e05;
    decBuf[2501] = 256'h6a0575057b0583058b058d058e05900593059205910592058f058e058c058705;
    decBuf[2502] = 256'h8705820580057f05790571056b05620557054c053d052b051b050305e704d404;
    decBuf[2503] = 256'hbb049f048c046c0457043c0423040104ea03d503b903a80392037e0371036503;
    decBuf[2504] = 256'h5a0358035703550359035b0357035f0360035a035b0355034b0347033e033203;
    decBuf[2505] = 256'h2d0325031c031d031a0315031703180315031a031c031d0327032e032f033903;
    decBuf[2506] = 256'h46034a035b03660370037f038a039403a003ac03ad03b903c203c303c703cd03;
    decBuf[2507] = 256'hcc03d303d403d203d803d903d403d903dd03de03e603ee03f303000412041e04;
    decBuf[2508] = 256'h35044b045f0477048c049b04b804cb04d604eb04fa0402050e0518051e052705;
    decBuf[2509] = 256'h2f05310537053b053c0547054f0553055c05680570057e058a059205a305ad05;
    decBuf[2510] = 256'hb305bf05c805cc05d605d905db05e205e205e005e205e205db05db05d305c405;
    decBuf[2511] = 256'hba05aa05970585056b055205430529051005fa04e604d404c804b904ab04a204;
    decBuf[2512] = 256'h970489048404760468045b044d043b042a041304fd03e903d103b5039a037a03;
    decBuf[2513] = 256'h5d03410322030403f102d102b402a0028f027902650258024702380226021a02;
    decBuf[2514] = 256'h1002fe01f201e701d901cd01c101b401a4019a018801770164014c0136012201;
    decBuf[2515] = 256'h0b01ee00d300bb009f0084006b005500410029001a000600f3ffe3ffd4ffc6ff;
    decBuf[2516] = 256'hbaffaeffa1ff94ff89ff79ff6aff5cff45ff2fff1bfffefee3fec3fea6fe83fe;
    decBuf[2517] = 256'h6cfe4efe33fe1afe0bfef7fde9fdd9fdcafdc4fdb8fdb0fda8fd9efd98fd95fd;
    decBuf[2518] = 256'h94fd91fd96fd9cfda2fdadfdb9fdc3fdcffdd8fde2fdecfdf4fdfafd03fe0cfe;
    decBuf[2519] = 256'h16fe20fe2dfe3dfe50fe63fe78fe92feb1fecffeeafe0aff30ff54ff74ff9aff;
    decBuf[2520] = 256'hbeffe8ff0f0033005d008400a800c800de00f900110121012f0142014e015801;
    decBuf[2521] = 256'h620172017d01870193019b01a501af01b301b801bb01bb01ba01b901b401ae01;
    decBuf[2522] = 256'hac01a6019f0198019001830176016801560140012c010f01f400dc00c0009d00;
    decBuf[2523] = 256'h7c005f00440024000600ebffccffaeff93ff7aff64ff56ff44ff38ff29ff23ff;
    decBuf[2524] = 256'h1aff15ff0bff01fff8feeafedcfec9feb6fea1fe8dfe75fe65fe51fe3ffe2efe;
    decBuf[2525] = 256'h1ffe11fe05fefafdeffde0fdd2fdc6fdb7fda9fd9afd8bfd81fd74fd66fd60fd;
    decBuf[2526] = 256'h54fd42fd3bfd2cfd16fd02fdeafccefcb3fc93fc6dfc53fc2afc02fce9fbbffb;
    decBuf[2527] = 256'h98fb74fb4afb23fbf5fac9faa2fa7efa54fa2dfa09fae8f9c2f9a9f991f974f9;
    decBuf[2528] = 256'h60f948f92cf918f9f9f8dbf8c0f8a0f883f868f848f82af80ff8f7f7e7f7d9f7;
    decBuf[2529] = 256'hc6f7bff7bdf7b7f7b9f7bef7bff7c9f7d7f7e3f7f8f712f82af846f869f88af8;
    decBuf[2530] = 256'hb0f8d4f8fdf825f953f97ff9b1f9e1f90dfa4bfa74faa9fae7fa20fb55fb93fb;
    decBuf[2531] = 256'hcdfb01fc4dfc7ffcbffcf8fc3cfd7cfdc6fd0cfe4cfe96fedcfe1cff66ffacff;
    decBuf[2532] = 256'hecff26005a008a00c300f7001a0145016d019101ba01d601f001100226024102;
    decBuf[2533] = 256'h52026802760289029502a402b202be02c602d302dc02e802ef02f602fa02fd02;
    decBuf[2534] = 256'hfa02f902f702ed02e602dd02d102c902be02b202a7029c029002840277026402;
    decBuf[2535] = 256'h560246023702290219020a020002f801ef01e801e401e001dd01d801d201ca01;
    decBuf[2536] = 256'hc001b301a5018f017a01630147012c010c01ee00cb00ab008500610037001000;
    decBuf[2537] = 256'hecffb9ff89ff5dff36fffefec9fe99fe61fe2cfeeefdb5fd80fd42fd08fdc5fc;
    decBuf[2538] = 256'h85fc3bfc09fcb7fb6afb38fbe6fa99fa53fa13fac8f982f930f9f9f8b3f873f8;
    decBuf[2539] = 256'h29f8f7f7b7f77ef749f719f7edf6c6f698f678f65cf643f62cf61ff60bf601f6;
    decBuf[2540] = 256'hfef5f5f5f3f5f5f5f3f5fdf509f60ef621f639f649f668f68ff6b2f6dcf60ff7;
    decBuf[2541] = 256'h3ff777f7bbf7faf745f88bf8cbf825f97af9c7f921fa76fad9fa37fb8cfbeffb;
    decBuf[2542] = 256'h4cfcb9fc03fd7bfdcdfd34fe92fefffe66ffc4ff31007a00f3004401ab010902;
    decBuf[2543] = 256'h5e02c1021e037303d60334048904d60444058e05eb0540067706d1060e075b07;
    decBuf[2544] = 256'h8d07df071608480875089f08d308f60815093c09600977099509b009c209de09;
    decBuf[2545] = 256'hf109fc090b0a1a0a210a2d0a380a3a0a430a480a430a440a3e0a300a2a0a160a;
    decBuf[2546] = 256'hff09ef09cf09b209970970094c092c09fd08d108aa087c0850081d08ed07b507;
    decBuf[2547] = 256'h72073207f806b40675062a06e40592054505ff04ad0460040604b10364030a03;
    decBuf[2548] = 256'h9d023602d8016b010401a6003900b4ff5bffe9fe82fe0afe98fd31fdb8fc46fc;
    decBuf[2549] = 256'hdffb82fb14fbadfa50fae2f97bf91ef9b0f867f809f89cf752f7f5f6a0f653f6;
    decBuf[2550] = 256'h0df6bbf56ef528f5e8f4aef46af43df414f4dff3bdf39df381f368f35af34df3;
    decBuf[2551] = 256'h41f33ef33bf343f351f35cf378f393f3acf3d4f307f429f462f496f4d4f40ef5;
    decBuf[2552] = 256'h51f591f5ecf528f675f6cff63df786f7e4f751f8b8f816f983f9eaf97dfae0fa;
    decBuf[2553] = 256'h5dfbeffb78fcf5fc88fd11fe8efe20ffaaff4b00e2006b01e9017b0204038103;
    decBuf[2554] = 256'h3404ab044205cc054906db0664070508710822099909300ab90a130ba50b070c;
    decBuf[2555] = 256'h840cf60c5d0dd60d270eac0e050f560fbe0f00105510a210d41014115e117c11;
    decBuf[2556] = 256'haa11d311ea11fe11111217122612221215120912f811d511be118f1164113111;
    decBuf[2557] = 256'hf310b91085103910df0fa30f560fe80e9e0e260eb40d4d0dd40c620cde0b610b;
    decBuf[2558] = 256'hce0a450ac8093609ac080b087407eb064a06b20529058804f1036703c6022f02;
    decBuf[2559] = 256'ha60105016d00e4ff43ffacfe22fe82fdeafc88fce7fb50fbeefa4dfae1f957f9;
    decBuf[2560] = 256'hdaf868f8e4f767f7f5f68ef615f6c4f55df5e4f493f42cf4e9f394f347f301f3;
    decBuf[2561] = 256'hd3f289f257f22af200f2ccf1a9f18af163f149f132f114f109f1f7f0e8f0eaf0;
    decBuf[2562] = 256'he3f0e5f0f8f000f115f135f153f176f1a8f1cbf103f238f275f2c0f206f346f3;
    decBuf[2563] = 256'ha0f3f5f342f4b0f417f575f5e2f549f6c2f654f7b6f733f8c6f84ff9f0f987fa;
    decBuf[2564] = 256'h11fbb1fb49fcd2fc73fd36feb8fe5fff2100d8007e011602c6029c032c04e304;
    decBuf[2565] = 256'hb80582063907df07a1085809ff09c10a440bea0bad0c2f0dd60d6d0ef60e730f;
    decBuf[2566] = 256'h06108f100c119e1101127e12ef123913b21303144d148f14cc14ed141f153a15;
    decBuf[2567] = 256'h4315591560155a155f1546152f151115e614b41484143f14ed13a0134613f112;
    decBuf[2568] = 256'h8e121512a4111f11a2101010860fe50e4e0ec50d240d8c0c030c3e0b870a110a;
    decBuf[2569] = 256'h4e09970820085e07a70601066905b904120450039902f3013001ad00070045ff;
    decBuf[2570] = 256'hc2fe1cfe84fdfbfc5afcc3fb39fbbcfa4afac6f949f9d7f870f8f7f785f71ef7;
    decBuf[2571] = 256'hc1f653f6ecf5a9f53cf5f2f4b0f45bf424f4def39ef375f331f303f3daf2a6f2;
    decBuf[2572] = 256'h76f24af222f2f4f1d5f1b9f195f17ef169f155f152f148f14bf153f15af165f1;
    decBuf[2573] = 256'h7bf189f19cf1bbf1d0f1ebf10af228f24bf275f29cf2caf202f337f375f3bff3;
    decBuf[2574] = 256'h05f445f4a0f4f5f458f5b5f50af66df6e5f637f7bbf739f8aaf812f98af91cfa;
    decBuf[2575] = 256'ha6fa23fbb5fb3efcbbfc4efdfefd75fe0cffbdff3400f60079011f02b7026703;
    decBuf[2576] = 256'hde03750426059d053406e5065c07f3077c08f9088c09150a920a240bae0b070c;
    decBuf[2577] = 256'h790cfe0c570dc90d130e700ead0efa0e2c0f6c0f950fc90fec0f0b101c103610;
    decBuf[2578] = 256'h43104810531050104010381025100210e80fb50f850f4d0f090fb70e800e260e;
    decBuf[2579] = 256'hd10d840d160dcc0c6f0c020c7d0b240bb20a2d0ad4094109b8085f08cc074307;
    decBuf[2580] = 256'hc60613069c0505057c04ff036c03e3024202d6014d01cf003d00b4ff37ffc5fe;
    decBuf[2581] = 256'h40fec3fd31fda7fc2afcb9fb34fbdafa48fae6f969f9f7f890f832f8c5f75ef7;
    decBuf[2582] = 256'h00f7abf648f6ebf596f549f503f5b1f44ef40bf4cef381f33bf3fbf2b1f27ff2;
    decBuf[2583] = 256'h52f218f2e3f1b3f187f16bf147f127f11af1fff0e7f0d7f0c3f0b6f0aff0a0f0;
    decBuf[2584] = 256'h96f098f093f094f0a3f0a9f0bdf0dff0f6f014f146f168f194f1d2f1fbf13ff2;
    decBuf[2585] = 256'h7ff2b8f2fcf23cf375f3c8f315f45bf4adf4faf440f5a4f502f66ff6d6f634f7;
    decBuf[2586] = 256'ha1f708f881f8f3f85af9d2f944fac9fa22fb94fb19fc96fce7fc6cfde9fd5bfe;
    decBuf[2587] = 256'hc2fe3affacff3100ae0020018701ff017102d8023603a3030a046804bd042005;
    decBuf[2588] = 256'h7d05d2051f067906ce061b076107a107eb0731087108bb08ed082d0967098c09;
    decBuf[2589] = 256'hbd09e809040a280a490a5e0a6a0a7b0a7e0a870a8f0a8c0a8a0a880a7f0a770a;
    decBuf[2590] = 256'h6a0a5a0a4b0a310a190afd09d209ab097c0944091009e0089b085b081108cb07;
    decBuf[2591] = 256'h8b074107e706aa065d060306ae054b05ed0499043604bd036c0305038c021b02;
    decBuf[2592] = 256'hb3012001be004100cfff68fff0fe7efef9fd7cfd0afda3fc2bfcb9fb52fbd9fa;
    decBuf[2593] = 256'h67fae3f989f9f7f895f818f8a6f75cf7e4f672f628f6cbf55ef514f5b6f461f4;
    decBuf[2594] = 256'h2af4d0f394f35df317f3d7f29df269f239f20df2daf1b8f199f171f158f14af1;
    decBuf[2595] = 256'h3df131f12ef12bf12ef13bf142f151f16bf17cf192f1b7f1d1f1f1f118f23cf2;
    decBuf[2596] = 256'h65f298f2baf2f2f227f365f39ff3e2f322f46cf4b2f4f2f43cf596f5d3f536f6;
    decBuf[2597] = 256'h79f6cef61bf775f7b1f714f857f8acf80ff952f9a7f90afa67fabcfa1ffb7dfb;
    decBuf[2598] = 256'hd2fb35fc92fce7fc34fd8efde3fd46fea4fee0fe43ffa1fff6ff43009d00f200;
    decBuf[2599] = 256'h5501b20107026a02c8021d038003c30330047a04d7042c057905bf0511065e06;
    decBuf[2600] = 256'ha406f60643077507c707fe0744088408cf08010940097a09af09df090b0a320a;
    decBuf[2601] = 256'h600a7f0a9b0ab50acc0ae10aed0af80afb0a030b010bfe0af80aea0ada0acb0a;
    decBuf[2602] = 256'hb10a990a7d0a520a1f0afd09b8098b094009fa08bb0870081608c10774071a07;
    decBuf[2603] = 256'hc60679060b06c1056305f6048f043104c4033f03e6027402ef0196010401a200;
    decBuf[2604] = 256'h2500b3ff4cffd3fe61fefafd82fd10fda9fc4bfcdefb94fb37fbcafa80fa22fa;
    decBuf[2605] = 256'hcdf980f926f9eaf89df857f817f8ddf7a9f778f74df725f701f7e1f6ccf6b1f6;
    decBuf[2606] = 256'ha6f697f688f686f67ef681f687f68cf694f6a4f6aff6c9f6e2f6fef621f741f7;
    decBuf[2607] = 256'h67f795f7cef7f3f731f86bf89ff8ddf817f94bf997f9c9f909fa53fa99fac7fa;
    decBuf[2608] = 256'h11fb57fb97fbd1fb14fc54fc9efce4fc36fd83fdc9fd1bfe68fec2fe17ff64ff;
    decBuf[2609] = 256'haafffcff49008f00e2002f017501c70114025a02ac020f035203a703f4033a04;
    decBuf[2610] = 256'h8c04d9041f057105be05040644069e06db0628076e07ae07e8073a087108b708;
    decBuf[2611] = 256'hf70841098709c709010a440a840aae0af10a1f0b480b7c0bad0bcc0bf30b170c;
    decBuf[2612] = 256'h2e0c4c0c5f0c710c870c950ca20cae0cb90cbb0cc30cc20cba0cb60ca80c950c;
    decBuf[2613] = 256'h880c6e0c4e0c310c060cdf0bb10b780b440b140bcf0a8f0a550a030ab6098409;
    decBuf[2614] = 256'h1f09dd0888082508c70772070f07b2064406dd05650514058f043504c4035c03;
    decBuf[2615] = 256'hff0292022a02cd017801ff00ae004600e9ff7cff32ffd4fe67fe1dfec0fd6bfd;
    decBuf[2616] = 256'h08fdc5fc70fc23fcf1fbb1fb78fb43fb05fbdcfab6fa94fa81fa65fa4cfa3efa;
    decBuf[2617] = 256'h31fa25fa22fa1ffa1cfa24fa2bfa35fa43fa5afa70fa8afaa9fad0fae9fa1cfb;
    decBuf[2618] = 256'h3ffb6afb9dfbcdfbf9fb37fc60fca3fcd1fc0bfd4efd8efdc8fd0bfe5efe95fe;
    decBuf[2619] = 256'hdbfe2dff64ffaafffcff49008f00e10018015e019e01d8011b025b029502c902;
    decBuf[2620] = 256'h070330036503a303cc0300043e0468049c04da040305380576059f05c405f405;
    decBuf[2621] = 256'h200648066b068c06aa06cc06e4060a0723073b07580773078c07a207bc07cd07;
    decBuf[2622] = 256'he307f7070408150824082a083a084408460852085b085f0866086c086d087408;
    decBuf[2623] = 256'h7708730873087108670866085b084a083b0829080f08fe07db07bb079d077207;
    decBuf[2624] = 256'h4b072707fe06cb06a90670063c060c06e005a20579053505f504bc0478043804;
    decBuf[2625] = 256'hee03a80356030903af025a020d02b3015e01fb009e004900e6ff88ff33ffd0fe;
    decBuf[2626] = 256'h73fe1efebbfd5dfdf0fca6fc49fcdbfb92fb34fbdffa92fa38fafcf9aff969f9;
    decBuf[2627] = 256'h29f9eff8abf87ef844f810f8edf7c1f79af776f74df730f717f700f7f3f6e7f6;
    decBuf[2628] = 256'hd6f6d3f6d6f6ddf6eef601f719f735f760f787f7abf7def70ef846f87bf8b8f8;
    decBuf[2629] = 256'hf2f836f976f9c0f906fa46faa0faddfa2afb84fbd9fb26fc80fcd5fc22fd7cfd;
    decBuf[2630] = 256'hd1fd1efe78fecdfe1aff74ffc8ff15005b00ae00fb0055019101de0124026402;
    decBuf[2631] = 256'hae02f40234036e03a203d3030b043f0462048104b404c804e704040513052105;
    decBuf[2632] = 256'h36054905540564056c057405800582058c05910593058e058a0584057a056e05;
    decBuf[2633] = 256'h5f0551053e0521050d05ee04d004b504960478045d0436041204f203cc03a803;
    decBuf[2634] = 256'h87036a033f031803f402ca02a3027f0255022e020002d401ad017f0153012b01;
    decBuf[2635] = 256'hfd00d2009f006f0043001000d3ff99ff64ff34ffeffec2fe78fe46fe06febbfd;
    decBuf[2636] = 256'h75fd36fdfcfcb8fc78fc3ffcfbfbbbfb82fb4dfb0ffbc5fa93fa53fa09fad7f9;
    decBuf[2637] = 256'h85f94ef908f9c8f87ef84cf80cf8c1f78ff750f716f7e1f6a3f67af646f616f6;
    decBuf[2638] = 256'heaf5cef5aaf589f56cf551f538f528f50ff504f5fbf4f2f4eff4f2f4f0f4faf4;
    decBuf[2639] = 256'h09f514f526f540f552f56ef591f5b1f5d7f505f631f664f694f6ccf601f73ff7;
    decBuf[2640] = 256'h89f7cff70ff859f8b3f808f955f99bf9fff95dfab2fa15fb58fbc5fb2cfc6ffc;
    decBuf[2641] = 256'hdcfc26fd83fdd8fd3bfe7efeebfe35ff78ffcdff1a007400b000fd0043019501;
    decBuf[2642] = 256'hcc01120252028c02c102fe0238035e038e03ad03d403ee030e04240437044904;
    decBuf[2643] = 256'h52045b04620465046304610454044604380425040d04f703dd03be03a0037d03;
    decBuf[2644] = 256'h5d0336031303e902c2029e02740241021f02e701c1019101650133010301d700;
    decBuf[2645] = 256'h990070003b000b00d3ff9eff6eff43ff10ffe0feb4fe81fe51fe26fefefddafd;
    decBuf[2646] = 256'hb1fd89fd70fd46fd1ffd05fde5fcc7fcacfc8cfc6ffc53fc34fc16fcfbfbe3fb;
    decBuf[2647] = 256'hc6fbb3fb9bfb7efb6bfb4cfb36fb23fb0afbf5fae0fac9fab3faa5fa8dfa77fa;
    decBuf[2648] = 256'h69fa56fa41fa33fa25fa10fa07fafaf9e5f9dcf9cff9bff9b4f9aaf99af990f9;
    decBuf[2649] = 256'h82f975f96df960f953f94ff947f940f93cf939f93af93df93ef944f94ff957f9;
    decBuf[2650] = 256'h62f976f985f997f9acf9c1f9d8f9f4f908fa27fa45fa68fa88faaefad2faf3fa;
    decBuf[2651] = 256'h21fb4dfb75fbadfbe1fb12fc3dfc70fcaefce8fc1cfd5afd94fdc8fd14fe46fe;
    decBuf[2652] = 256'h86fed0fe16ff44ff8effd4ff01004c009200bf000a013c017b01b501f9012602;
    decBuf[2653] = 256'h60029502c502f0022303450371039903bc03dd03030427043e045c0477048804;
    decBuf[2654] = 256'h9e04b204c004cb04d204dc04e104e304de04d704d404c704b904af04a2048d04;
    decBuf[2655] = 256'h79046704510437041f040304ef03d003b203970378035a033f031803f402dd02;
    decBuf[2656] = 256'hb70293027c0256023c021c02fe01e301c301ae018b017d016001440133011d01;
    decBuf[2657] = 256'h0301f200e200ce00bc00b000a100930087007b0074006d006700630060005f00;
    decBuf[2658] = 256'h6200650065006a006c0073007c00830089008f0094009c00a800b000b800c100;
    decBuf[2659] = 256'hca00d400e100ec00fa00060111011f012701330140014d0155015f0169016f01;
    decBuf[2660] = 256'h75017c01840189018c019101970199019c019f019f01a001a301a601a501a001;
    decBuf[2661] = 256'h9e019901970192018c0184017f0176016d0167015e01560150014b0143013b01;
    decBuf[2662] = 256'h36012e012b01260122011f011901130112010f010b0108010701050106010a01;
    decBuf[2663] = 256'h0b010a010e0116011e0125012b013501410149015701670171017f018b019a01;
    decBuf[2664] = 256'hac01bd01cc01de01ee01fd0117022902380252026b0280029a02b302c202dc02;
    decBuf[2665] = 256'hf5021103240336034c036603770387039b03b203c203d003e303f30302041404;
    decBuf[2666] = 256'h2004330440044c045b0465046a047904830485049004950496049c04a204a104;
    decBuf[2667] = 256'ha404a604a504aa04a904a404a704a804a404a804a7049f049e049b0497049804;
    decBuf[2668] = 256'h93048b048f048e0488048c048d0488048f04960498049f04a504a704b404c204;
    decBuf[2669] = 256'hc404d304e504e704f60400050905170525052b053d054d055405660576058105;
    decBuf[2670] = 256'h9305a305ae05c005cc05db05ed05f405fa050806150616061e0622061e062106;
    decBuf[2671] = 256'h20061e061d0613060406fa05ee05d905ca05b80599058405610541052305f804;
    decBuf[2672] = 256'hd104ad047a044a041e04ec03ae03850350031203d802950267021d02eb01ab01;
    decBuf[2673] = 256'h61011b01db00a1004f001800d2ff80ff49ff03ffb1fe7afe34fef4fdbafd85fd;
    decBuf[2674] = 256'h48fd0efdd9fca9fc7dfc4bfc28fcfdfbd5fbb1fb9afb7dfb61fb50fb47fb32fb;
    decBuf[2675] = 256'h25fb1efb1cfb1efb20fb28fb32fb3ffb51fb66fb7afb92fbaefbd1fbf1fb0ffc;
    decBuf[2676] = 256'h3afc61fc85fcb8fce8fc14fd51fd8bfdc0fdf0fd35fe74feaefef2fe32ff6bff;
    decBuf[2677] = 256'hafffefff28005d009b00d500180146017f01b401f2011b0250028002b802ec02;
    decBuf[2678] = 256'h0f033b036d039d03bd03ef0312043104580472048904a704ca04e104ed040905;
    decBuf[2679] = 256'h1a052a0538054505510560056a05730578058205860585058805870585058605;
    decBuf[2680] = 256'h85057f057e05780571056f056a05640563055a0550054f0547053c0535052505;
    decBuf[2681] = 256'h17050f05f604e504d504bb04a3048d046d04500434041504ef03d503ab038403;
    decBuf[2682] = 256'h6a0338031503e902b70287025b022802f801c0017c013d010301bf007f003500;
    decBuf[2683] = 256'hefff9dff50fff6feb9fe6cfe12febefd5bfdfdfcc0fc5dfc00fcabfb5efbf0fa;
    decBuf[2684] = 256'ha6fa48faf4f991f94ef9e1f897f854f8fff7b2f76cf72cf7e2f6b0f65ef627f6;
    decBuf[2685] = 256'hf5f5c7f58df559f537f517f5f0f4ccf4bef4a0f495f48af487f48af492f49ef4;
    decBuf[2686] = 256'hadf4cbf4e8f40bf535f55cf58af5c3f5f7f535f67ff6c5f605f760f79df700f8;
    decBuf[2687] = 256'h5df8b2f8fff86df9d4f932fa9ffa06fb64fbd1fb38fcb1fc22fd6cfde5fd56fe;
    decBuf[2688] = 256'hbefe36ff87ffeeff6700b8001f017d01ea0134029102e60233038d03e2031904;
    decBuf[2689] = 256'h5f049f04c8040c05390563058805ab05ca05e60500060d0623062e0632063506;
    decBuf[2690] = 256'h380635062e06230615060606f305db05b905a1057b0557052e050605d804a004;
    decBuf[2691] = 256'h7a043d040304dd039f0366032203e202a90274023602ec01ba017a013001fe00;
    decBuf[2692] = 256'hac0075002f00efffb5ff72ff32ffe7feb5fe63fe2cfefafda8fd71fd2bfdebfc;
    decBuf[2693] = 256'hb2fc6efc2efce4fb9efb5efb24fbe1faa1fa67fa24fae4f9aaf967f927f9edf8;
    decBuf[2694] = 256'hb8f86df83bf8fbf7d2f79df752f720f7f2f6a8f676f648f60ef6daf5aaf571f5;
    decBuf[2695] = 256'h3df51bf5eff4bcf49af46ef447f42df40df4eff3dcf3c3f3adf3a5f392f38bf3;
    decBuf[2696] = 256'h8df383f388f391f398f3aaf3bbf3c9f3e7f30ef427f451f478f4a6f4d2f410f5;
    decBuf[2697] = 256'h4af58df5cdf507f659f6a6f6ecf63ff7a2f7e4f752f8b9f816f984f9ebf948fa;
    decBuf[2698] = 256'hcefa27fb99fb1efc9bfcecfc71fdeefd60fec7fe3fffb1ff1800910002016a01;
    decBuf[2699] = 256'hc70134029c02f9024e03b1030f044b049804f2042f057c05c205f00529065e06;
    decBuf[2700] = 256'h8006ac06d306e306fa060f07230726072907260719070d07fa06e306c606a406;
    decBuf[2701] = 256'h7a0653062406ec05b8057a054005fd04bd0472042c04da038d033303de029102;
    decBuf[2702] = 256'h3702e30196013c01e70084002600d1ff6eff11ffbcfe59fefbfda6fd43fd00fd;
    decBuf[2703] = 256'habfc48fc06fcb1fb64fb0afbcdfa80fa3afafaf9c0f97df93df903f9def8aef8;
    decBuf[2704] = 256'h75f850f820f8f4f7cdf7a9f788f76bf748f731f71bf708f7f0f6e6f6d2f6c5f6;
    decBuf[2705] = 256'hbef6aff6a9f6abf6a3f6a1f6a8f6a4f6a8f6b5f6b6f6bef6d2f6dff6ebf6fef6;
    decBuf[2706] = 256'h10f726f73af74cf76bf789f79cf7bcf7daf7edf713f837f84ef875f8a3f8c2f8;
    decBuf[2707] = 256'he9f818f937f969f99af9c5f903fa2cfa61fa9ffad9fa0dfb4bfb85fbb9fb05fc;
    decBuf[2708] = 256'h37fc77fcc1fc07fd47fd91fdc3fd15fe62fea8fee8fe32ff78ffb8ff13005000;
    decBuf[2709] = 256'h9d00e30035016c01b20104023b029502d10208034e038e03d9030b044a048404;
    decBuf[2710] = 256'hc804f5042f0564058605be05e405060625064d06660687069c06af06c106d006;
    decBuf[2711] = 256'hdf06e706e906eb06ed06eb06e706df06d006c206b2069b0685066b064c062e06;
    decBuf[2712] = 256'h0b06e105ba059605630533050705e004a804730443040b04d60398035f033903;
    decBuf[2713] = 256'hfb02c1028d024f021502e101b101780144010601dd00a800780040001a00eaff;
    decBuf[2714] = 256'hbfff97ff73ff4aff2eff0affe9fed4feb9fe99fe8dfe72fe60fe57fe48fe3bfe;
    decBuf[2715] = 256'h39fe37fe31fe36fe38fe39fe45fe54fe5efe6efe81fe8efea3febdfed6feecfe;
    decBuf[2716] = 256'h0bff21ff43ff64ff82ffa4ffceffeaff1800440060008400b700d90005013801;
    decBuf[2717] = 256'h5a018601b801db0107022e025c027b02ae02d002fc0223033d0367038e03a803;
    decBuf[2718] = 256'hc803e603010420043e045204710486049a04b204c804d604e904f90404051205;
    decBuf[2719] = 256'h1e05260531053d05420547054b054c054f0552055005520553054b054a054705;
    decBuf[2720] = 256'h3f053e053b05320530052a0520051f051b05130512050e05060507050205fa04;
    decBuf[2721] = 256'hfb04fa04f404f804f704f104f704f704f004fe040005fa0406050d0509051405;
    decBuf[2722] = 256'h1f051d052e0538053605460555055b056705760580059305a005a705ba05c805;
    decBuf[2723] = 256'hd305e705f405fb0512061c062406370642064d065b066406690676067f068406;
    decBuf[2724] = 256'h910697069806a606ab06ad06b706bb06ba06c206c706c406cc06cd06c606d206;
    decBuf[2725] = 256'hd306c906cd06ce06c606c706c606bd06be06bd06b506b606b306ab06aa06a706;
    decBuf[2726] = 256'h9f06a306a0069b06a306a0069906a306a406a006a606a906aa06b306b506b106;
    decBuf[2727] = 256'hbd06c206c106ca06d106cd06d806dd06d906e406e806e706ed06f106ee06f406;
    decBuf[2728] = 256'hf106ed06f306f006e806ee06e906dc06da06d506c606c006b406a20691067e06;
    decBuf[2729] = 256'h6c0656063c0624060e06e905c505a4057e0550053105fe04ce04a20470044004;
    decBuf[2730] = 256'h1404e103a3037a0337030903cf028c025e022402e101a10167013301f500bb00;
    decBuf[2731] = 256'h870049000f00daffaaff72ff3eff0dffe2feaffe7ffe60fe38fe0afeebfdcffd;
    decBuf[2732] = 256'hb5fd9efd89fd75fd6bfd62fd59fd56fd54fd56fd58fd61fd6cfd80fd92fda7fd;
    decBuf[2733] = 256'hbcfddefdf5fd1bfe3ffe5ffe8efebafee1fe0fff3bff6eff9effd6ff0b004800;
    decBuf[2734] = 256'h8200b700f5003f017101b101fb012d026d02a702ea022a0364038903c7030104;
    decBuf[2735] = 256'h350465049e04c304f3041f0546056a059405b005d405f4050a0625063d064d06;
    decBuf[2736] = 256'h610673067f068e0698069a069f06a306a206a3069d0694068c067f0671066306;
    decBuf[2737] = 256'h4f063d0628060e06ee05d905b6059605780555052c050f05ec04c2049b046c04;
    decBuf[2738] = 256'h41041904f503c303a003680342031203da02a60275024a021702d9019f016b01;
    decBuf[2739] = 256'h3b01f600c8007e0038000b00d1ff7eff47ff01ffc1fe88fe44fef2fdbbfd75fd;
    decBuf[2740] = 256'h23fdecfca6fc54fc1dfcd7fb85fb38fbf2fab2fa68fa22facff998f93ef902f9;
    decBuf[2741] = 256'hb5f86ff81df8e6f78cf74ff702f7bcf67cf642f60ef6c2f590f550f517f5f1f4;
    decBuf[2742] = 256'hc1f489f472f442f423f4fcf3d8f3c1f3abf390f37ff375f367f35ff361f357f3;
    decBuf[2743] = 256'h55f361f366f373f387f394f3aef3cdf3e3f306f438f45bf487f4b9f4e9f422f5;
    decBuf[2744] = 256'h65f5a5f5dff522f674f6c1f607f747f7a2f7f7f744f88af8eef831f99ef9e8f9;
    decBuf[2745] = 256'h46fa9afae7fa41fb96fbf9fb57fcacfcf9fc53fda8fdf5fd3bfe9ffee2fe37ff;
    decBuf[2746] = 256'h84ffcaff0a0054009a00da00240156019601bf01f4012402500277029b02bb02;
    decBuf[2747] = 256'hd902ec02fe0214031c032403300332032c03310329031f0312030103eb02dd02;
    decBuf[2748] = 256'hc002a50285025f0231021202ea01b2018c014f011501e000a20058001200d2ff;
    decBuf[2749] = 256'h88ff42fff0fea3fe5dfe0bfea8fd65fd10fdadfc6afc15fcb2fb55fb00fbb3fa;
    decBuf[2750] = 256'h59fa04faa1f943f9eef88bf849f8f4f791f733f7def67bf638f6e3f580f53ef5;
    decBuf[2751] = 256'he9f49cf456f404f4b7f371f31ef3d1f29ff260f226f2f1f1b3f17af154f124f1;
    decBuf[2752] = 256'hf8f0dcf0aef082f071f04ef036f02af016f005f0fbefedefeaeff2efebefedef;
    decBuf[2753] = 256'h00f0feef0ef02ef03cf051f074f08bf0b2f0e0f00cf133f16bf1a0f1def117f2;
    decBuf[2754] = 256'h5bf29bf2e5f217f369f3b6f3fcf34ef4b1f4f4f449f5acf5eff55cf6a6f603f7;
    decBuf[2755] = 256'h58f7bbf719f886f8edf830f99df905fa62fab7fa30fb81fbe9fb46fcb3fc1bfd;
    decBuf[2756] = 256'h78fdcdfd30fe8efecafe2dff8bffe0ff2d008700c30010015601a901e0012602;
    decBuf[2757] = 256'h65029f02d40204033c0371039303bf03e6030a042a044804630475048b049904;
    decBuf[2758] = 256'ha104a804ae04b004a8049f0495048604700456043d042104f703db03ac038103;
    decBuf[2759] = 256'h4e031e03e602b10273023a02f601b6016c013a01e8009b0055001500baff65ff;
    decBuf[2760] = 256'h18ffd2fe80fe33fed9fd84fd37fdc9fc80fc3dfcd0fb86fb43fbeefa8bfa48fa;
    decBuf[2761] = 256'hf3f9a6f960f920f9d6f890f850f817f8e2f7a4f77bf746f716f7f7f6d0f6acf6;
    decBuf[2762] = 256'h8bf66ef653f648f638f62af627f61cf619f61ff625f62df63af647f65cf676f6;
    decBuf[2763] = 256'h8ef6b0f6daf6f6f624f75df791f7c1f7f9f72ef86cf8b6f8fcf83cf986f9ccf9;
    decBuf[2764] = 256'h1efa6bfab1fa03fb50fbaafbfffb4cfca6fcfbfc5efda1fd0efe58feb6fe0aff;
    decBuf[2765] = 256'h6dffb0ff1d006700c5001a016701c10116026302a9020d035003a503f2033804;
    decBuf[2766] = 256'h7804d2040f0546058c05cc05060649067706c106f30621074a077e07ae07ce07;
    decBuf[2767] = 256'h000823084e0876088f08b008d608e50806091b09360948095e096c097e098a09;
    decBuf[2768] = 256'h8c099a09a0099e09a209a10998099509920985097b096f0959094b0933091e09;
    decBuf[2769] = 256'h0f09f208cf08b8089b08780857083a080f08f307c507990772074e071207e806;
    decBuf[2770] = 256'hc30685065c062706e905c0057d054f051505e104950463043504eb03b9038c03;
    decBuf[2771] = 256'h52031d03df02a602800242021902e501c2018a01640142011601ef00cb00ab00;
    decBuf[2772] = 256'h950073005200450032001a0016000800fbfff9fffbfff9ff01000d0014002600;
    decBuf[2773] = 256'h37004a0067008a00a100c700f500140147017701a301d60113024d028202cd02;
    decBuf[2774] = 256'hff023f038903cf030f045a04a004df043a057705c4050a065c06a906ef062f07;
    decBuf[2775] = 256'h7907d30710085d08a308e3081c096009a009d9091d0a5d0a860aca0af70a200b;
    decBuf[2776] = 256'h550b770b970bbe0bd80b010c1d0c2d0c440c590c5d0c6e0c780c750c780c7a0c;
    decBuf[2777] = 256'h740c760c690c570c500c410c230c170c030ce40bc60bab0b8b0b6e0b4b0b180b;
    decBuf[2778] = 256'hf60ad60aa40a740a540a160aed09c8098a0961092c09fc08c4088f085f083308;
    decBuf[2779] = 256'h0108c3079a07650735070907d706a6067b0648061806f905c60596056a054305;
    decBuf[2780] = 256'h1505f504ce04a0048104590435041504ef03cb03b403960373035c0347032403;
    decBuf[2781] = 256'h0d030003e502d302be02a902a2028c027e0276026a025b025902540249024402;
    decBuf[2782] = 256'h43023a023b023e023a023c02420247024d0255025d026c0276027c029002a202;
    decBuf[2783] = 256'hae02c502db02ef020703230336034f0371038803a603c103da0302041e043804;
    decBuf[2784] = 256'h620489049804c204e90403052d05490562058c05b305cd05ed0514062d064e06;
    decBuf[2785] = 256'h74068306a406c106dd06f50611071d0735074b075407660777077d078b079007;
    decBuf[2786] = 256'h8f0796079207890786077b076e07650753073e0729071207f606db06b4069006;
    decBuf[2787] = 256'h70064a061b06f005bd058d0561052305ea04b50469043704f803ad0367032703;
    decBuf[2788] = 256'hdd0297024502f8019e0161011401ba007e001b00d8ff83ff36ffdcfe9ffe3cfe;
    decBuf[2789] = 256'hfafda5fd58fd12fdc0fc73fc41fceefba1fb6ffb30fbe5fab3fa73fa3afa05fa;
    decBuf[2790] = 256'hd5f99df977f947f91bf9f4f8d0f8b0f892f877f85ef849f834f822f81bf810f8;
    decBuf[2791] = 256'h06f808f806f808f812f818f822f831f83ff856f86cf886f89ef8baf8ddf8fdf8;
    decBuf[2792] = 256'h24f948f971f999f9bcf9eff91ffa4bfa7efaaefae6fa1bfb59fb82fbb6fbf4fb;
    decBuf[2793] = 256'h2efc62fca0fccafc0dfd3bfd74fdb8fde6fd1ffe54fe84feb0feeefe17ff3cff;
    decBuf[2794] = 256'h6cffa5ffcaffedff1800400064008400a200bd00dc00f2000d01250135014301;
    decBuf[2795] = 256'h50015c0167016d016f01730175016e016801640157014b014001290113010501;
    decBuf[2796] = 256'he800c500ae0090006e004d0027000300d9ffb2ff84ff58ff26fff5fecafe8cfe;
    decBuf[2797] = 256'h52fe2dfeeffdb5fd80fd43fdf8fcc6fc86fc4dfc18fccdfb87fb59fb0ffbc9fa;
    decBuf[2798] = 256'h9bfa51fa0bfacbf991f94ef90ef9d4f891f863f819f8e7f7a7f76df739f708f7;
    decBuf[2799] = 256'hc4f696f66df638f6faf5d1f5acf57cf55cf535f507f5f4f4cdf4a9f492f47cf4;
    decBuf[2800] = 256'h61f450f43af42cf424f413f40df40ff409f40bf413f414f41ff433f43bf450f4;
    decBuf[2801] = 256'h70f485f498f4bff4d8f402f529f54df580f5b0f5dcf51af654f688f6c6f600f7;
    decBuf[2802] = 256'h43f783f7cdf713f853f89df8e3f836f983f9c9f91bfa7efac1fa15fb78fbbbfb;
    decBuf[2803] = 256'h10fc73fcb6fc0bfd58fdb2fd07fe54fe9afeecfe39ff7fffbfff09004f008f00;
    decBuf[2804] = 256'hc900fd003b017501a901d90105022d0250027a029602b002d002dd02f0020203;
    decBuf[2805] = 256'h0503080310030d030303f902e902da02c802a9028b0270024a022602fc01d501;
    decBuf[2806] = 256'h9d01680138010001cb008d0043001100bfff88ff42fff0fea3fe5dfe1dfec2fd;
    decBuf[2807] = 256'h86fd39fddffca2fc3ffcfcfba7fb70fb16fbdafa8dfa47faf4f9bdf977f938f9;
    decBuf[2808] = 256'hedf8bbf87bf842f80df8ddf7b1f773f74af725f702f7d7f6baf6a1f68af66cf6;
    decBuf[2809] = 256'h59f647f637f62ff627f620f61ef624f622f62af63ef645f656f669f67cf696f6;
    decBuf[2810] = 256'hb5f6d3f6f6f61ff73cf76af795f7c8f7f8f724f857f894f8cef803f94ef994f9;
    decBuf[2811] = 256'hc2f90cfa52fa92fadcfa22fb74fbc1fb07fc5afca7fc01fd55fda2fde8fd3bfe;
    decBuf[2812] = 256'h9efee0fe35ff98fff6ff33009600f30030019301f00145029202d8022a038d03;
    decBuf[2813] = 256'hd00325047204b8040a0557058905db0528065a069a06e506170756079007b607;
    decBuf[2814] = 256'he6071e08440866089208b908d308f30808091c0934093e094c09540951095809;
    decBuf[2815] = 256'h56094a094109340921090909ed08d208b9089108690845081308e207aa077607;
    decBuf[2816] = 256'h3807fe06bb067b063006ea05980561050705b20465040b04b7036a031003bb02;
    decBuf[2817] = 256'h5802fa01a5014201e50090004300d5ff8bff2dffd8fe75fe33fedefd7bfd38fd;
    decBuf[2818] = 256'he3fc96fc50fcfefbb1fb7ffb3ffbf5fac3fa83fa49fa24fae6f9bcf997f975f9;
    decBuf[2819] = 256'h55f939f920f908f9f3f8e8f8ddf8d4f8cbf8cef8cbf8d6f8e0f8e9f8fbf80bf9;
    decBuf[2820] = 256'h23f93ff95af979f9a0f9c3f9e4f913fa3efa71faaffad8fa0dfb4afb84fbc8fb;
    decBuf[2821] = 256'h08fc41fc85fcc5fc0ffd55fd95fddffd25fe77fec4fef6fe48ff95ffdbff2d00;
    decBuf[2822] = 256'h7a00c00013016001a601f80145028b02cb0215035b039b03e5032b046b04a504;
    decBuf[2823] = 256'he80428057205a405e4051e0652069006b906ee062c0755077b07ab07d607fe07;
    decBuf[2824] = 256'h2208420868088c08a308c108dc08ee080409180925093509400946094f095409;
    decBuf[2825] = 256'h5209590955094d094c09410932092c091d090509fc08e208c308b6089b087408;
    decBuf[2826] = 256'h5b083a081408fa07d1079e077c0750072907fa06cf069c067a0641060d06dd05;
    decBuf[2827] = 256'ha505700540050805d304a3046b0436040604ce03990369033103ee02c0028602;
    decBuf[2828] = 256'h52022f02f701c301920167013f011101e500b300900065003d0024000300ddff;
    decBuf[2829] = 256'hb9ffa2ff7cff6cff4cff37ff1cff0afffbfee6fed9fecdfec7feb9feb0feabfe;
    decBuf[2830] = 256'ha7fea8feaafea6fea9feaffeb5febcfec3fed0fedbfee6fef8fe0dff1bff28ff;
    decBuf[2831] = 256'h3eff52ff6aff7fff94ffabffc1ffdbfffaff10002b0043005f007b009a00af00;
    decBuf[2832] = 256'hca00ea00080123014201580173019201a701c301db01f70112022b023a025402;
    decBuf[2833] = 256'h6d027c029102a802b802c602d902e902f8020603120321032f03340340034703;
    decBuf[2834] = 256'h4e0354035c036103640365036403660365035f0360035e035603550352034603;
    decBuf[2835] = 256'h41033a0333032a03200314030c030103ef02e302d902cb02be02b0029e029202;
    decBuf[2836] = 256'h8702750269025b024d0240023202240217020902fb01ef01e301d601c901be01;
    decBuf[2837] = 256'hb401aa019c018c0186017c0170016b01630157014f01470141013d0135012e01;
    decBuf[2838] = 256'h280123011d011b01160114010f01060102010301fd00f600f400f300f200ef00;
    decBuf[2839] = 256'hed00e800e700e300df00da00d900d500d100ce00cb00c700c300be00ba00b500;
    decBuf[2840] = 256'haf00a900a5009f009c00990092008a00870081007a0074006b00610060005800;
    decBuf[2841] = 256'h51004b0045003d003700320027001f001d0014000b0007000000f9fff3ffecff;
    decBuf[2842] = 256'he8ffe3ffddffd3ffcfffccffc6ffc1ffbbffb5ffb4ffafffa9ffa7ffa4ffa1ff;
    decBuf[2843] = 256'h9fff9cff98ff95ff93ff90ff8fff8cff88ff87ff86ff84ff83ff80ff7eff7dff;
    decBuf[2844] = 256'h7aff77ff75ff72ff71ff70ff6eff6bff6aff68ff63ff62ff60ff58ff55ff54ff;
    decBuf[2845] = 256'h4fff4bff46ff42ff3eff36ff2eff2dff27ff1dff1cff18ff10ff0bff09ff02ff;
    decBuf[2846] = 256'hfcfef4feedfeecfee5fedafed5fed1fecafec6fec0febbfeb9feb6feaefea9fe;
    decBuf[2847] = 256'ha6fea1fe9dfe99fe96fe95fe91fe90fe91fe8bfe84fe85fe86fe87fe86fe84fe;
    decBuf[2848] = 256'h81fe84fe84fe84fe88fe89fe86fe8bfe8dfe8cfe91fe92fe92fe97fe99fe9afe;
    decBuf[2849] = 256'h9dfe9efe9ffea1fea2fea1fea4fea5fea6fea7fea7fea7fea7fea8fea7fea5fe;
    decBuf[2850] = 256'ha2fea1fea0fe9afe96fe93fe8bfe84fe83fe7cfe73fe6ffe66fe5afe55fe4afe;
    decBuf[2851] = 256'h3efe36fe28fe1ffe14fe07fef7fdecfddafdcafdbffdadfd9cfd8dfd7ffd6cfd;
    decBuf[2852] = 256'h5ffd4efd3bfd2efd19fd0afdfdfce8fcd4fcccfcb7fca2fc95fc85fc72fc64fc;
    decBuf[2853] = 256'h54fc45fc37fc27fc18fc0efcfffbf0fbe6fbd9fbcefbc4fbb7fbacfbaafba3fb;
    decBuf[2854] = 256'h9dfb98fb91fb8cfb88fb83fb83fb82fb81fb80fb83fb85fb88fb8afb8ffb97fb;
    decBuf[2855] = 256'h9ffba2fba9fbb4fbbafbc3fbcdfbdafbe5fbf3fbfbfb0afc1cfc2dfc3bfc49fc;
    decBuf[2856] = 256'h59fc6cfc7ffc8ffca7fcbdfcd1fce3fcf8fc0dfd24fd3afd54fd6cfd7cfd96fd;
    decBuf[2857] = 256'haefdc4fdd8fdf0fd0cfe27fe40fe56fe70fe8ffea4febffed8fef4fe07ff20ff;
    decBuf[2858] = 256'h3cff57ff70ff86ff9fffb8ffd4ffe7ff00001c002f004800640077008900a500;
    decBuf[2859] = 256'hb800d100e100f5000c011c013001420158016c0179018e019d01aa01bb01c501;
    decBuf[2860] = 256'hd301df01ee01f8010102090216021c0224022b02320236023c02410243024602;
    decBuf[2861] = 256'h4502420241023f023c023a0233022f022b0223021b0216020c020002f501e701;
    decBuf[2862] = 256'hd701c801b601a6019701850170015b014901340120010801f200d800c000a400;
    decBuf[2863] = 256'h88007000540039001900fbffe0ffc1ffa3ff80ff69ff43ff29ff09ffebfec8fe;
    decBuf[2864] = 256'ha8fe8afe6ffe4ffe32fe0ffef8fdd1fdb8fd97fd7afd5ffd46fd2afd0ffdf6fc;
    decBuf[2865] = 256'he0fcccfcb5fc9ffc8bfc78fc63fc4ffc3cfc31fc22fc18fc0bfc03fcfcfbf2fb;
    decBuf[2866] = 256'he9fbe6fbe3fbe2fbe1fbe0fbe0fbe6fbe7fbedfbf5fbfcfb05fc11fc1bfc2afc;
    decBuf[2867] = 256'h3cfc4dfc5cfc72fc86fc98fcaefcc2fcd9fcf6fc11fd29fd45fd60fd80fd9efd;
    decBuf[2868] = 256'hb9fdd8fdf6fd19fe39fe60fe83fea4fec2fee4fe0eff2aff4eff78ff94ffb8ff;
    decBuf[2869] = 256'he1fffdff21004b0067008b00ab00d200f5000d013301570177019501b001cf01;
    decBuf[2870] = 256'hed01080221023d02600277028c02a702c002dc02ef02080317032c033e034f03;
    decBuf[2871] = 256'h6203740380038f039d03a903b803c203ca03d303e003e503ed03f203f603f703;
    decBuf[2872] = 256'hfb03fc03fe03ff03fd03fd03fb03f603f403ee03e203dd03d603cc03c103b403;
    decBuf[2873] = 256'ha7039c038e037f0370035a034b033903240315030303ee02d902c202ac029802;
    decBuf[2874] = 256'h80026402490237021b020002e801cc01b0019f01830168014f0133011001f900;
    decBuf[2875] = 256'hdb00c800af009300780060004a002a001500faffe8ffd2ffb9ffa0ff8aff76ff;
    decBuf[2876] = 256'h5eff49ff3aff2dff1cff0eff00fff3fee1fed6fecbfec1feb8feb0fea9fea2fe;
    decBuf[2877] = 256'h9bfe98fe93fe94fe95fe94fe95fe94fe97fe97fe9cfea4feacfeb5febdfec5fe;
    decBuf[2878] = 256'hccfed8fee0feedfef9fe08ff16ff22ff34ff45ff54ff62ff75ff87ff98ffabff;
    decBuf[2879] = 256'hbdffceffe1fff4ff090017002a003f0053006600760089009c00ac00bf00d200;
    decBuf[2880] = 256'he700f6000801190127013901450154016201720181018f019801a301b001bd01;
    decBuf[2881] = 256'hcb01d101da01e501ed01f401fd01020205020b02100216021a021d021e022002;
    decBuf[2882] = 256'h23022202250224022502240221021f021a02160211020f020a0208020302fd01;
    decBuf[2883] = 256'hf501f201eb01e301db01d401cc01c201b901b001a8019f01990193018c018401;
    decBuf[2884] = 256'h7a016e0162015501490141013901320127011c0113010a010001f900f000e600;
    decBuf[2885] = 256'hdd00d400cc00c300ba00b200ad00a5009e0097008f00870080007a0075006f00;
    decBuf[2886] = 256'h670064005f005900540054004f004d004c004700430042003e003d003e003b00;
    decBuf[2887] = 256'h380038003700380038003600370039003a003d003e003f004100460046004600;
    decBuf[2888] = 256'h4a004d005100540058005c00610067006b006e007200770079007c0080008500;
    decBuf[2889] = 256'h89008c008e00910095009a009e00a200a800ad00b300b600ba00c000c400c500;
    decBuf[2890] = 256'hca00cc00cd00d200d600da00e000e300e400e700eb00ee00f000ef00f200f500;
    decBuf[2891] = 256'hf400f300f500f600fb00fd00fc00fc00fc00fc00fb00fd00f900f600f700f500;
    decBuf[2892] = 256'hf000f100f000ee00ed00e800e600e500e200e000db00d900d800d300cd00cb00;
    decBuf[2893] = 256'hca00c500c100be00ba00b600b100ad00a800a2009e009a00950091008c008c00;
    decBuf[2894] = 256'h8700860084007f007d0078007600730070006e006b0069006400630064006300;
    decBuf[2895] = 256'h6100620061005e005b005b005b005b00580059005a0059005a005c005b005b00;
    decBuf[2896] = 256'h5b005e0062006500660067006800670069006c006d0070007400750077007700;
    decBuf[2897] = 256'h76007700770077007700780079007c007b007a007b007c007900780077007700;
    decBuf[2898] = 256'h7400730070006e006d006a00680062005d00590053004d004a00470043003d00;
    decBuf[2899] = 256'h35002d00260022001a0014000b000200fbfff2ffe6ffdfffd8ffcfffc5ffbbff;
    decBuf[2900] = 256'hb0ffa6ff9cff93ff8eff83ff78ff6fff68ff60ff57ff4cff45ff3eff35ff2dff;
    decBuf[2901] = 256'h22ff1bff14ff0bff03fffcfef8fef2feeafee4fedffedefedcfed7fed5fed0fe;
    decBuf[2902] = 256'hcafec8fec3fec2fec1fec2fec3fec2fec3fec4fec5fec6fec7fec8fec8fecbfe;
    decBuf[2903] = 256'hccfecffed3fed7fedcfee2fee8feebfef1fef3fefbfe03ff0aff10ff18ff20ff;
    decBuf[2904] = 256'h27ff2fff34ff3dff46ff4eff59ff61ff67ff6eff76ff7dff84ff8cff91ff9bff;
    decBuf[2905] = 256'ha2ffabffb5ffbeffc5ffcfffd8ffe1ffedfff6fffaff010007000d0014001a00;
    decBuf[2906] = 256'h22002a00310037003d00410047004c005000530057005a005c00630067006b00;
    decBuf[2907] = 256'h6e006f007000710071007400770078007800790077007600750072006e006d00;
    decBuf[2908] = 256'h6900660063005f005c005c0054004e0047003f003a003300270022001b001400;
    decBuf[2909] = 256'h0e000600f9fff0ffe5ffddffd4ffcbffbeffb3ffa9ff9cff8eff84ff77ff6cff;
    decBuf[2910] = 256'h61ff55ff4aff3fff30ff22ff16ff07fffdfef1fee2fed4feccfebdfeb3fea7fe;
    decBuf[2911] = 256'h9bfe91fe84fe79fe6ffe62fe57fe52fe49fe3dfe36fe2ffe24fe1ffe16fe0ffe;
    decBuf[2912] = 256'h0afe05fe00fefafdf4fdf0fdedfdebfde4fde4fde3fde4fde6fde9fdeafdecfd;
    decBuf[2913] = 256'hedfdecfdf1fdf3fdf8fdfefd02fe07fe10fe17fe1bfe25fe29fe2ffe3cfe44fe;
    decBuf[2914] = 256'h4bfe55fe60fe6bfe74fe7dfe85fe92fe9bfea0feadfeb6fec1feccfed8fee7fe;
    decBuf[2915] = 256'hf9fe00ff0aff18ff21ff29ff31ff3aff43ff50ff5bff65ff72ff7aff81ff88ff;
    decBuf[2916] = 256'h91ff99ffa2ffa8ffb0ffb9ffbdffc0ffc5ffcbffd0ffd6ffd8ffddffe3ffe7ff;
    decBuf[2917] = 256'hecffeeffeffff0fff3fff4fff3fff4fff4fff4fff4fff4fff3fff2ffefffebff;
    decBuf[2918] = 256'he8ffe6ffe1ffdfffdaffd6ffd1ffcbffc3ffbeffbbffb5ffb0ffafffa9ffa7ff;
    decBuf[2919] = 256'ha2ffa0ff9aff93ff8dff85ff80ff79ff73ff6dff65ff5fff58ff50ff48ff3fff;
    decBuf[2920] = 256'h37ff31ff2cff24ff1eff17ff10ff0aff03fffdfef7fef1fee9fee3fedcfed8fe;
    decBuf[2921] = 256'hd3fed1fecbfec8fec5fec3febefeb8feb4feb1feaffeaafea8fea3fe9ffe9efe;
    decBuf[2922] = 256'h9bfe9afe9bfe9afe9bfe9cfe9bfe9efea1fea0fea1fea5fea4fea5fea9feaefe;
    decBuf[2923] = 256'hb0feb5febbfebffec7fecdfed4fedcfee1fee6feecfef2fef9fe02ff09ff0fff;
    decBuf[2924] = 256'h17ff20ff29ff33ff3dff48ff52ff59ff60ff67ff70ff7cff86ff90ff9bffa9ff;
    decBuf[2925] = 256'hb1ffbdffc7ffd1ffdcffeafff2fffeff08000f00180024002c0034003d004400;
    decBuf[2926] = 256'h4e00570060006800710077007f0084008a0094009b009f00a400ab00b300bd00;
    decBuf[2927] = 256'hc100c500cd00d200d600db00dd00e000e400e700ea00ea00eb00ec00ef00ee00;
    decBuf[2928] = 256'hef00f100f100f300f600f500f200f100ef00ec00eb00ea00ea00e900e400e300;
    decBuf[2929] = 256'he300e000df00db00d500d200cf00cb00c500c000ba00b800b300ad00a900a400;
    decBuf[2930] = 256'h9e009a0096008f008d00880082007c0076006e0069006600610060005e005800;
    decBuf[2931] = 256'h5700520049004500410040003f003e003900390038003300340032002d002900;
    decBuf[2932] = 256'h26002200210022001f001e00210022002400250028002c003100320036003900;
    decBuf[2933] = 256'h39003e004000430047004e0054005d0067006d0075007c007f0085008b008e00;
    decBuf[2934] = 256'h95009d00a400b000b800bc00c300cc00d600e200f100fb00070113011a012701;
    decBuf[2935] = 256'h2f013901400146014e01590167017301820190019801a401ab01af01b601bd01;
    decBuf[2936] = 256'hc001c801d501e001ee01fa01050213021b0224022b0235023b0245024c025002;
    decBuf[2937] = 256'h55025a025f0265026b027502810290029a02a602ae02ac02ae02aa02a902a802;
    decBuf[2938] = 256'hab02ab02b002b202b702bf02c402c902d102d502d202d102d202cd02ce02cd02;
    decBuf[2939] = 256'hcb02cb02cb02c402c502ca02c902cb02cc02c602c402bc02af02a7029d029302;
    decBuf[2940] = 256'h8a0282027b027b02760270026c0264025c0255024b023f0237022c0220021802;
    decBuf[2941] = 256'h0a02fe01ef01e501dd01d501d001c601c001b601aa019b018901740160014801;
    decBuf[2942] = 256'h38012a011d0116011801160111010801fb00eb00dc00ca00ba00af009d009600;
    decBuf[2943] = 256'h9000860080007f0077007300740071006a0064005a00530048003e0031002900;
    decBuf[2944] = 256'h22001b001c001b001e00260029002e002f002c002a002900260025002a002900;
    decBuf[2945] = 256'h2b003000310035003b00400046004e0053005a005d005e0060005f005b005800;
    decBuf[2946] = 256'h59005c0064006c0071007a0084008a009000950096009700960097009d00a100;
    decBuf[2947] = 256'ha400ac00b100b400b900bd00c000c600c800c900c800c600be00ba00b300ad00;
    decBuf[2948] = 256'hab00ac00ac00b100b300b400b700b100ab00a600a2009c009b009a009b009e00;
    decBuf[2949] = 256'h9e009800920087007b00770070006a006d006c00680065005f0057004f004000;
    decBuf[2950] = 256'h310027001b0010000e000a00060008000300fcfffafff4ffefffedffe8ffe2ff;
    decBuf[2951] = 256'hdcffcfffc1ffb5ffa9ff9fff9dff9fffa2ffa7ffa4ffa2ff9dff90ff82ff73ff;
    decBuf[2952] = 256'h64ff56ff4dff45ff40ff42ff3eff3bff38ff31ff2fff2cff2aff29ff2bff2cff;
    decBuf[2953] = 256'h2aff25ff18ff0aff01fff3fee9fee7fee9feeafef1fef7fef8fef9fef7feeffe;
    decBuf[2954] = 256'he5fed6fec8febbfeb0feabfeadfeaefeb4febffec6fecdfed3fed4fed9fedafe;
    decBuf[2955] = 256'hd4fecbfec1feaefea1fe9afe98fe9afea6feb5fec3fecffed1fed2fecefec0fe;
    decBuf[2956] = 256'hb4fea9fe98fe8dfe87fe86fe87fe8ffe98fea1feabfeb2feb8febcfeb5feaffe;
    decBuf[2957] = 256'ha9fe9dfe92fe8afe7bfe75fe70fe6bfe6dfe76fe7ffe89fe90fe8ffe89fe7efe;
    decBuf[2958] = 256'h68fe52fe3efe21fe0dfe03fe06fe09fe16fe1dfe28fe32fe30fe32fe2dfe23fe;
    decBuf[2959] = 256'h18fe0bfef0fdd5fdc4fdaefdabfdb3fdbafdc9fdd7fddcfddbfdd6fdc4fdaffd;
    decBuf[2960] = 256'h9bfd7efd6afd60fd57fd59fd67fd72fd81fd8ffd95fd99fd9bfd97fd8efd88fd;
    decBuf[2961] = 256'h7dfd76fd72fd71fd76fd7dfd83fd8bfd91fd92fd9afd9ffda4fdaefdb5fdbbfd;
    decBuf[2962] = 256'hbefdbdfdbbfdbcfdbefdc1fdccfddbfdedfd07fe20fe35fe4afe61fe6bfe79fe;
    decBuf[2963] = 256'h7cfe79fe77fe79fe7bfe86fe9afeb1fecdfee9fe01ff1dff31ff3bff44ff4dff;
    decBuf[2964] = 256'h55ff57ff59ff5bff68ff76ff88ffa7ffcdffe7ff1100220031003f0043003f00;
    decBuf[2965] = 256'h3c003f004d0060007a009900bf00d900f000f400f800ee00e400d600d300d600;
    decBuf[2966] = 256'he000f600100129013f01530160016201640162015d0158015101520156015e01;
    decBuf[2967] = 256'h6b017e018b019c01a201a0019b0190017f01700162015201480142013d013e01;
    decBuf[2968] = 256'h40013e0142014301420141013f0137012f012401190110010701fb00ec00de00;
    decBuf[2969] = 256'hce00c800c200c000c500ca00cb00c700bb00a20083005d002f000f00fefff9ff;
    decBuf[2970] = 256'hfeff13002e004700560059004c0037001700f1ffc3ff97ff7bff6cff70ff85ff;
    decBuf[2971] = 256'ha8ffd2fff9ff130018000b00f0ffc2ff8aff64ff34ff15ff0fff1fff36ff5cff;
    decBuf[2972] = 256'h8affaaffd1ffd6ffd1ffbcffa1ff82ff6cff59ff55ff59ff6dff8affa5ffc4ff;
    decBuf[2973] = 256'hd9ffedfff7fffafffdfffbfffdfffffff9fff0ffe5ffd5ffceffd4ffddfff5ff;
    decBuf[2974] = 256'h1c00400073009500c100dd00e200e700da00bf00ad009e0095009d00b700dd00;
    decBuf[2975] = 256'h0c0144017801a801d401e501e001c0019101650132011e01180134016c01b001;
    decBuf[2976] = 256'h02024f029502b002b8029302700238020402e101db01ec0106022f026202a002;
    decBuf[2977] = 256'hc902df02e602e002c402aa027702470228020c0207020b0229024c0276029202;
    decBuf[2978] = 256'hab02b002a3028002600231020602f501e501e101ed01f901fd01f301eb01d801;
    decBuf[2979] = 256'hcc01c201b801b901b801ad01990173013b010601c9008f0087008000a000c700;
    decBuf[2980] = 256'heb000b0118010501d0007e003100ebffabffa3ffaaffdaff06002d0047004200;
    decBuf[2981] = 256'h2d000200c5ff8bff47ff1aff01ffeafef1fef8fe08ff18ff26ff2aff26ff1cff;
    decBuf[2982] = 256'h06ffecfec5fe97fe78fe67fe62fe79fea8fed4fefbfe0aff06ffe8feb6fe78fe;
    decBuf[2983] = 256'h3efe18fef6fdf0fd01fe25fe57fe7afe99feaafea5fe8efe67fe44fe23fe0efe;
    decBuf[2984] = 256'h0afe15fe2afe3ffe56fe6cfe75fe7dfe88fe8bfe89fe8afe85fe81fe82fe81fe;
    decBuf[2985] = 256'h80fe83fe84fe7ffe7ffe7ffe80fe86fe90fe9cfeaefebafec5fec7fec2feb3fe;
    decBuf[2986] = 256'ha5fe92fe7ffe78fe72fe78fe92fec4fe02ff4dff93ffc0ffd9ffd1ff94ff39ff;
    decBuf[2987] = 256'hccfe64fe07fee2fdd7fd1dfe94fe26ffb0ff09003a000e00b0ff2bffadfe1bfe;
    decBuf[2988] = 256'hb9fd83fdb4fd1bfe94fe26ffafff2d005d004f000c009ffffcfe65fe03fe86fd;
    decBuf[2989] = 256'h75fd67fdaafd17fe7efef6fe68ff94ff87ff4affe7fe6ffefdfd96fd6efd62fd;
    decBuf[2990] = 256'h99fdf3fd48fe95fec7febdfeb5fe81fe51fe25fe09fe04fe08fe0cfe10fef8fd;
    decBuf[2991] = 256'hc9fd8bfd51fd3bfd42fd6dfdc2fd17fe7afebdfec9febefe64fef7fd8ffd17fd;
    decBuf[2992] = 256'hc6fc99fcc2fcfefc77fde9fd6efeebfe1cff48ff3affe6fe6dfedafd51fdd4fc;
    decBuf[2993] = 256'h83fc74fcd1fc57fd1bfe07ffa5fffbff15009eff07ff2ffe66fde3fc9cfcddfc;
    decBuf[2994] = 256'h66fd2bfee2feb7ff470061004a00ddff54ffd7fe65fe1bfe0efe32fe7ffed9fe;
    decBuf[2995] = 256'h47ffaefff1ff15000a00ecffacff72ff3eff29ff3cff63ffa6fff8ff45007700;
    decBuf[2996] = 256'h93009b00750045000000c1ff97ff9fffddff3700bd003a018b019a0172010501;
    decBuf[2997] = 256'h6200cbff69ff57ff88ff0d00ad00700127026e0259021e027d01ba0003008dff;
    decBuf[2998] = 256'h77ffb2ff2f00e2008801f401560244021402ca015101e00096006e0062008300;
    decBuf[2999] = 256'hc9001b016801ae01db01d3019f015301f900a4006d004f006b00b5000f016401;
    decBuf[3000] = 256'hc7010a021602f501af014a01d200810054006200b7003001c20124027d026d02;
    decBuf[3001] = 256'h4102ae01fd005700c0ff5dff6fffe1ffa10058012d02bd02d702c0025302ca01;
    decBuf[3002] = 256'h4d01db00910069005d007e00c40016017901f20143028d02b502a9025c02c601;
    decBuf[3003] = 256'h2e015600c7ff78ff90ff2700d800dd01d1027003c6037703d102e30106017600;
    decBuf[3004] = 256'h5c0074000b0195013502a202b502a30273022902e601da01cf01ed011a023302;
    decBuf[3005] = 256'h2c020902d1017f0148013e016b01d6015b02d8026b03a50394036303de028502;
    decBuf[3006] = 256'h1302e701bf01cb01ec011e025e029702ea024d039003e503f003d2036d03da02;
    decBuf[3007] = 256'h29028301ec00b1000a019d019c029003ac046c058f057005e004f503d8021802;
    decBuf[3008] = 256'h6a014a01a00157022d03f603ad04f4040a05a80407047003bf0248020702f401;
    decBuf[3009] = 256'h29027b02ff02a0030c046f04a404b404a6047e0441040a04d80386033903df02;
    decBuf[3010] = 256'hba02af02e1024603a30311045a044d041004c30355030c03c902bd02b202d002;
    decBuf[3011] = 256'hfd0247038d03f203350471047c0472043204e8038e033903ec02a60279026002;
    decBuf[3012] = 256'h58027b02b3020603530385038e0375033103f202b80292027e0277028802a202;
    decBuf[3013] = 256'hd50205033d0354034d032103d80292025202290212020b020502e901c5019c01;
    decBuf[3014] = 256'h8b019001b90103025d029902a40286024602db0174011601da00cf00d9001801;
    decBuf[3015] = 256'h6301a901fb0132023c023302f901a6012d01bc005400dcffabff7fffa7fffcff;
    decBuf[3016] = 256'ha10047010a028d02750234025c01590065ff88fe6bfe85fe2bff1900f700c001;
    decBuf[3017] = 256'h43025a02ee013e01680065ffb7fe19fe35fe4ffec6fe89ff0b00b200f3002d01;
    decBuf[3018] = 256'h1c01eb00a1000e0085ffe4fe78fe3dfe4ffea0fe60ff1600bd0054018f013601;
    decBuf[3019] = 256'ha300cbffc9fe1afe7cfd5ffde2fd88fe76ff5400e300fd00e6004e009efff7fe;
    decBuf[3020] = 256'h8bfe50feaafe5dff0300c5001401cd00600089ffbffe08fec1fd02fe64fe05ff;
    decBuf[3021] = 256'h9cffffff1000000099ff56ff01fff6fe00ff40ff8affe4ff2100580062005900;
    decBuf[3022] = 256'h3000fbffbdff73ff2dffedfea3fe5dfe1dfe04fe1bfe66fee8fe65ffd7ff2100;
    decBuf[3023] = 256'h2e00f2ff79ff07ff82fe29fe19fe45fea2fe40ff0300ba0060017501ec00e0ff;
    decBuf[3024] = 256'h87fe42fdc7fb2efb5cfb2ffc88fdcdfe9fff1300350097ffcefe17fe71fd05fd;
    decBuf[3025] = 256'h18fd72fde4fd68fee5fe37ff45ff1dfff9fe96fe38fee3fd6afdf9fc91fc34fc;
    decBuf[3026] = 256'hf7fbd6fb08fc7ffc11fd9afd18fe48fe1cfed9fd54fdfafccafcbbfcc8fc05fd;
    decBuf[3027] = 256'h52fd70fd8bfd73fd4dfd0ffdc5fc93fc65fc5dfc83fcb3fcebfc10fd17fddffc;
    decBuf[3028] = 256'h6ffcdcfb53fbfafae9fa33fbc6fb77fc4dfddcfd2bfe13fed2fd49fda8fc10fc;
    decBuf[3029] = 256'h87fb2efbfdfa29fb87fb0cfcadfc44fdcefd03fef3fd6efdaafcbffba2fae2f9;
    decBuf[3030] = 256'h7af999f929fa14fb31fc3dfd31fe90fe74fef1fd1bfd18fc6afbccfa76fac4fa;
    decBuf[3031] = 256'h6afb2dfce4fc5bfd9bfd88fd52fde0fc5cfcbbfb23fbc1fa68fa58fa66faa9fa;
    decBuf[3032] = 256'h2ffbacfb3efca0fcfafc0afdfbfceefcc9fcbefca0fc85fc5cfc27fcf7fbbffb;
    decBuf[3033] = 256'h7bfb4efb24fb0efb07fb26fb64fbbffb14fc61fc93fc8afc50fceefb76fb04fb;
    decBuf[3034] = 256'h9dfa75fa81fae4fa92fb68fc31fdb4fdcbfd5ffdaffc7afb53fa46f9def8bef8;
    decBuf[3035] = 256'h4ef939fa16fbe0fb96fcdefcf3fcb8fc3bfccafb45fba4fa38fad6f9a0f9b0f9;
    decBuf[3036] = 256'hfaf958fac5fa2cfb8afb96fb75fb2ffbb8fa46fadff982f975f980f9c6f92bfa;
    decBuf[3037] = 256'ha3fa15fb5ffb87fb93fb72fb2cfbdafa77fa19fac4f9a3f999f9a2f9ccf9e2f9;
    decBuf[3038] = 256'he9f9d6f9c5f9c0f9d7f917fa8efa00fb49fb71fb4dfbeafa72fa00fab6f9c4f9;
    decBuf[3039] = 256'h31fab5fa33fb84fb75fb32fbadfa30fabef9aff9f2f977fa3cfbf3fb6afc7ffc;
    decBuf[3040] = 256'h44fcc7fb35fbd3fa7afa49fa75fab8fa25fb8cfb05fc56fc82fc90fc83fc62fc;
    decBuf[3041] = 256'h44fc4efc66fc8cfca0fca7fca1fc92fc96fcbdfcfffc64fda6fde3fdeefdbcfd;
    decBuf[3042] = 256'h6afd1dfdc3fc86fc4ffc45fc61fc8afccdfc32fdaafd3cfe9ffe1cff8dfff5ff;
    decBuf[3043] = 256'h38005c0051000b0082ffaafee1fd5efd17fd58fd09fedefea8ff5e0076003500;
    decBuf[3044] = 256'h85ff7ffe8bfdedfc97fc1afdc0fd04ff490070013002de02fe02a702f0014a01;
    decBuf[3045] = 256'h8800d1ff5aff19ffdefef0fe41ff8bffe9ff3e005f0069004d002400efffcdff;
    decBuf[3046] = 256'hbaffc0ffdaff0c004a00a500fa005d01bb010f0230023a023102e7018d012001;
    decBuf[3047] = 256'hf400e600f200290147012c01b0000f004dffcafee2fe4eff4d008701ae026e03;
    decBuf[3048] = 256'h9103f302b6018f0083ffd4fe33ff3600b6011b035f04de04b704c303a7024d01;
    decBuf[3049] = 256'h6500e7ffc1ffe3ff82004b01cd01440285029902630232020602c3019f019401;
    decBuf[3050] = 256'h76017f019801db015202e40295030b047804b2047d042c04a70306036f02e501;
    decBuf[3051] = 256'h68011701260183012102e302cf032d0484046a04f3035b0321030f0380032304;
    decBuf[3052] = 256'hba044305790569051f05c10485047a048404c404ed040305ef04aa044604e803;
    decBuf[3053] = 256'h93039e03e4036d041e05c40530066b06a106900682068f06b306be06b4068706;
    decBuf[3054] = 256'h4d060906dc05e4050a0647068106980691067e066d065e0675069b06b506c306;
    decBuf[3055] = 256'had068306670662068b06e00695074c082209b209cc098509c208d707ba06fa05;
    decBuf[3056] = 256'h4c052c054905cc05a206a4075308300986096c09f50833084807aa0653066d06;
    decBuf[3057] = 256'h140702081e092b0ad90aba0a2a0a3f092208c906e10562058905370615075108;
    decBuf[3058] = 256'h23094a092709c808ff077c0735071f0733076907ba07040846088308e6085e09;
    decBuf[3059] = 256'hd009370a600a3b0aac09fc08f60748076b061406c605de05f3052e068806f906;
    decBuf[3060] = 256'h6107be072b087508b808f5080009f608b6085b08d60735079d068a06bf067207;
    decBuf[3061] = 256'h77086b09490a9f0a1c0a4709d107060656043d033e0210028e02e703e6054a08;
    decBuf[3062] = 256'he5095b0b170b5d0a64088806d804300463044a05710631079a07b9076307e106;
    decBuf[3063] = 256'h990684069706a9067806f4052f051004b602ce01a401cb01790214049d056807;
    decBuf[3064] = 256'h9d08d50808092008f90653053a043b03b0028602ad025b033804c8044b056205;
    decBuf[3065] = 256'h4d05c304ff0314033602a70158017001b1011302900202036903e1035304d804;
    decBuf[3066] = 256'h31054205f8047f048c039802ba012a0110015801c40126025b024b02c6014901;
    decBuf[3067] = 256'hb7002e00f8ff080035009200e7003401a201ec01140251025c027a0283027a02;
    decBuf[3068] = 256'h4602fa017801d700150092ff1bff06ff19ff2bff7dffa9ff9bff8fff6eff50ff;
    decBuf[3069] = 256'h59ff72ff7aff81ff7aff5eff63ff84ffc3ff4c00d6002f013f01f600480072ff;
    decBuf[3070] = 256'h6ffec1fd23fdccfce7fc5dfd20fed7fe4eff8eff54fffafe68feb7fd41fdd4fc;
    decBuf[3071] = 256'he8fc1efdb0fd88fe8bff39009800b5006600c0ffd2fef5fd2bfda9fc32fcc6fb;
    decBuf[3072] = 256'h8bfb79fb89fbb6fb2efcc0fc71fd47fe10ff5eff17ff54fe35fd8ffb76fa43fa;
    decBuf[3073] = 256'h72faedfbb8fd68ff81001a018f0068ffc2fd39fcd4faecf9c2f99bf904fa63fa;
    decBuf[3074] = 256'h2cfbaffb25fc66fc7afc21fccffb68fb40fb4cfb99fbdffb1ffc38fc30fc1cfc;
    decBuf[3075] = 256'h09fc1afc52fca5fc08fd4afd3efdc5fcf2fbb6fa3bf9d6f7eef6c4f684f778f8;
    decBuf[3076] = 256'h13fa2bfb2afcb6fce0fc6dfcbefb20fb90faaafaf2fa5efb99fb63fbb0fadbf9;
    decBuf[3077] = 256'h11f9c3f80af923fa30fb6afce8fc75fc81fbe6f95df892f6d9f5a1f5a0f6e4f7;
    decBuf[3078] = 256'h5ff92afbdbfcf3fd26fe9bfd20fc55fa20f908f8d5f703f8d6f8e2f991fab0fa;
    decBuf[3079] = 256'h93fa11fa6bf9a8f825f8def7c8f752f816f936faf6fa5efb3ffbaffac4f9e6f8;
    decBuf[3080] = 256'h57f871f817f930fa3dfba5fbc5fb35fb4afa6df9ddf88ff8d6f842f97df96bf9;
    decBuf[3081] = 256'hf9f83af883f73bf751f7daf7c3f8dff99ffa08fb28fb98fae1f93bf9cff86cf8;
    decBuf[3082] = 256'h7ef8d0f854f9d1f943fa8dfad0faf4fabdfa4ffaadf9eaf833f8bdf7d2f734f8;
    decBuf[3083] = 256'hd5f86df9cff9e1f98ff9edf856f8f4f729f8fdf839fab4fbb3fc3efdc0fcb3fb;
    decBuf[3084] = 256'heef93df895f7fcf62af7fdf770f81ff97df99af9b4f99df9b2f99ff9d4f905fa;
    decBuf[3085] = 256'h4ffaacfad1fac6fa80faf7f995f93bf96cf90efa27fb81fcc5fd98fe72fe7efd;
    decBuf[3086] = 256'he2fbe9f985f7eaf50af5c6f47ff508f7d3f8fffa74fc40fd7efd46fdadfcc5fb;
    decBuf[3087] = 256'h47fb6dfbd6fbb3fc7cfdcbfde3fd4bfd4cfc12fb40fa80f95df9bcf94bfacefa;
    decBuf[3088] = 256'he6fad0fa20fa79f9b7f868f851f8bdf895f997fa17fce2fd92ff1b011a02ec01;
    decBuf[3089] = 256'h1901c0ffc2fd6efc39fb01fbcefa59fbd7fb4afcb3fcd3fcb6fc67fcf1fb59fb;
    decBuf[3090] = 256'ha9fa32faf1f92cfa85fa38fb0efcd7fcc2fda0fea2ff9600740191010e01aaff;
    decBuf[3091] = 256'h45fea3fc8bfb58fbe3fb0afd16fe0aff2aff9afe7bfd6efcc0fb61fbf1fbdcfc;
    decBuf[3092] = 256'hf9fd05ffb4ff12002f00e1ff9aff84ff70ffa6ffd7ffc8ffa0ff4bffbcfe0bfe;
    decBuf[3093] = 256'h65fdf9fcbefcacfcddfc27fd9ffd11fe5bfe4dfe11fec4fd92fd9bfdb3fdf7fd;
    decBuf[3094] = 256'h49fe96fe04ff89ff71004f0151020003e00250023101d8ff36feadfcaefbc6fa;
    decBuf[3095] = 256'h9cfac3fab7fb13fdb4fe3d00a2012d0257029701a30087ff7afe11fe31fec1fe;
    decBuf[3096] = 256'h78ff1e00b500f000ba004900a6ff0fffd4fee6fef6fee8fea5fe1ffe5bfda4fc;
    decBuf[3097] = 256'h2dfc6efc1ffd83fee8ff8901a202d5020303850212026301440127010d015401;
    decBuf[3098] = 256'h3e012b01f5008300ffffa5ff75ff66ffa9ff2e00cf006601f00125023602b101;
    decBuf[3099] = 256'h10014d0096ff4fff65ffeeffd700f301000368038803bf02d401f6002d001300;
    decBuf[3100] = 256'h2b00970020017a0169013d01fa00a5009a00f400aa013203bb04200608073207;
    decBuf[3101] = 256'hbf0685055e0405031d029e01c5012d020b039b0386042405b4050206bb052305;
    decBuf[3102] = 256'hfd0382021d013500b7ff90fff9ffd60066011d02c3028603a504fe0543076a08;
    decBuf[3103] = 256'hdd08ba081c08e006650566042103a302c9023203d00399045005c70533064606;
    decBuf[3104] = 256'h58064806fe058605d3042d04c103d4032e04e10487051e06a8062507b7076808;
    decBuf[3105] = 256'hde081f09bd08d507790634056204ee038603660310035902e201cd010802f002;
    decBuf[3106] = 256'h0d0419050d062d061006f6050e067a062b0700089008de089708d50752070b07;
    decBuf[3107] = 256'h4c0723082609d509330aa4098408de06e50491035c02240257029c03c3041c06;
    decBuf[3108] = 256'h04078207a9078607660749072f0718070207ee06dc06ac066206cf05f7042e04;
    decBuf[3109] = 256'h77035f03f603f6042f0656071608f30794073e07bc06a4061007e807eb08240a;
    decBuf[3110] = 256'h4b0b0b0c2e0c900bc70adc0980089807c5069f0636061706fa057705a104d803;
    decBuf[3111] = 256'h21030a03a103c7049706c208380a040b420b0a0b710ae60967094109d8087908;
    decBuf[3112] = 256'h23086c07c60603064d05d6046a047d04fa04ad05b206a7078408140962094a09;
    decBuf[3113] = 256'hb3085108f7070808aa08c309d00a0a0cdc0c030d9a0c3b0ce50b620bbc0aa309;
    decBuf[3114] = 256'hfd077406a904f902e00147017501f401b40262033f0442057c064f070e087708;
    decBuf[3115] = 256'h570801087f07370778077708b109d80a980bbb0bdd0adb09a108ce075b077e07;
    decBuf[3116] = 256'h9e07ba0738073206f904d20312037a0358040706b707d00869093b0968085b07;
    decBuf[3117] = 256'had060f06f2050c0624060e06ac052f055c045903ab020d02f0013e02e402a703;
    decBuf[3118] = 256'h5e0476043504ab030b03ca020503c903e90442062a07fc0770084d082d08d707;
    decBuf[3119] = 256'hbd07d407ea07d6077d0789064f058003540149fff5fdc0fcf8fc5dfeb8009d03;
    decBuf[3120] = 256'h55061a086c088c07b005840379012500e7ff1f00b80043011901a600b2ff14ff;
    decBuf[3121] = 256'hf7fe1600bc01b5039105cf05b7042002a6ffc2fcd0fa76fa6dfbe2fcbefeea00;
    decBuf[3122] = 256'h8b03b906dd08070aad0912080606a20363018200b6ff79ff40ff73ff45ff6fff;
    decBuf[3123] = 256'h49ffb1ff10002d007b006400230072ff6dfe79fd9bfc0cfc26fc0efc24fc37fc;
    decBuf[3124] = 256'h02fc32fcb7fca0fdbcfe7cffe5ffc5ff89fe62fd09fc21fb4bfb0bfc8afdeffe;
    decBuf[3125] = 256'h3400b2008c002300c4ffa8fff6ff6d00d900ed00280009ffaffdc7fcf5fb82fb;
    decBuf[3126] = 256'h5ffb00fb70fa22fadaf9c5f9b1f97cf90af968f8d0f76ef7ebf7dff8eafaf5fc;
    decBuf[3127] = 256'hd1fe8bffc3ffc4fe7ffd04fc39fa04f95cf88ff81af9edf9f9fa62fb81fbb8fa;
    decBuf[3128] = 256'hcdf9b0f8a4f781f71ff85bf9d6fad5fba7fbd4fa2ef935f7e1f5a3f5bcf687f8;
    decBuf[3129] = 256'h37fa30fc84fdc2fd1afd81fc3cfb6afaaaf941f9e2f88cf8a1f784f6c4f55cf5;
    decBuf[3130] = 256'hbbf584f606f7bff67bf5c3f2d2f0c2ef70efe6f04af340f421f5edf5a6f6bff7;
    decBuf[3131] = 256'h56fa84fd83007402cf02d801a2fec8fa29f7def3baf157f1fcf04ff199f155f1;
    decBuf[3132] = 256'h18f150f14ff293f3baf4c7f5a4f506f503f40ff332f2a2f1b7f09aef41eeb6ed;
    decBuf[3133] = 256'he0ed86ef60f2dff52af94dfbb1fbecf9acf776f453f2eff195f1e7f1c7f293f3;
    decBuf[3134] = 256'h4cf4f5f45af6fbf784f9b7f92cf9b1f7e6f5b1f409f4d6f3eef273f1dceeadeb;
    decBuf[3135] = 256'h8ae926e936ead1eb72eeebf03df1f3f0aff071f019f17ef220f4a9f576f58ef4;
    decBuf[3136] = 256'hbef20ef1d6f06ff16df349f57ef646f67bf4d3f10ff074eebeee12f0c3f1dbf2;
    decBuf[3137] = 256'ha8f21df24bf124f18df12bf2bbf23df385f31cf41bf555f67cf73cf8d3f7b6f6;
    decBuf[3138] = 256'h10f587f322f2f4f172f27ff32df48cf4c3f33bf2b2f04defc2ee95efeef0d6f1;
    decBuf[3139] = 256'h58f165ef79ec87eae2eac6ed0df209f69ff818f9f4f63cf4c2f1cbf016f1e2f1;
    decBuf[3140] = 256'h9bf2b4f3b3f4f8f5c7f76efa33fccefd83fda7fb00f987f647f467f323f360f3;
    decBuf[3141] = 256'hb8f253f10ef03ceffcef07f2a7f421f7bcf807f93bf88bf672f53ff56df5ecf5;
    decBuf[3142] = 256'h12f635f655f638f61ef606f647f6a9f64af70df85bf8e4f7cbf625f52cf350f1;
    decBuf[3143] = 256'h97f05ef05df1a2f271f49df63ef902fb9efc13fe57fe9efdf6fc91fb4cfa25f9;
    decBuf[3144] = 256'h7ff786f5aaf3faf1c2f127f3def55ef9b8fbdbfd3ffee4fd92fd47fd8bfd44fe;
    decBuf[3145] = 256'hedfebafed2fd03fcd7f9ccf768f571f491f3d5f38ef417f67cf7aaf72cf7d2f5;
    decBuf[3146] = 256'h8ef467f38df3c7f442f6a7f78ff8b6f95cfb55fd4100fa02be0459060f06cb05;
    decBuf[3147] = 256'h1105d904a60478045103ab0142ff02fdf7faa3f9e9f8b1f87ef850f87af83af9;
    decBuf[3148] = 256'he8f9c6fac8fb02fd29fe82ffc7004501d20053ff22fd81fabcf8c6f7a6f8faf9;
    decBuf[3149] = 256'h26fc31fe95003002a6030a06ee08e00aa40c520cb10983068403cc00bcff6aff;
    decBuf[3150] = 256'h1fffdbfe22fe7afd79fe1a00f402ac05260878082d08d906a4058c042703e201;
    decBuf[3151] = 256'h670002ffd4fea6ff9901fd039805e3059f056a0452035302810257021703c503;
    decBuf[3152] = 256'h21051f07fb08270b9d0c690da60d6e0da10d160d440c9d0ac4070b05dd01defe;
    decBuf[3153] = 256'hedfcddfbe7fa9cfa68fb18fd62008e05610ac20ebf125515af171d18b917aa16;
    decBuf[3154] = 256'h0e1503139f105f0e540c6809b006cc023600ccfe5ffe89ff4e01e9025f04a304;
    decBuf[3155] = 256'he104890588068608ea0ace0d4e11991497178919981aa1190117d213af11bd0f;
    decBuf[3156] = 256'h630f100f300ecc0b430808042f01a2ff29ff72009c016103fc040707f309730d;
    decBuf[3157] = 256'hae11aa1541189b1a2d1a031989160113b60fb70cc60a200bbc0c5c0f21111812;
    decBuf[3158] = 256'h37115b0fab0d730d720e2a11e213f214fb13f011040f120db80c9c0f1b135717;
    decBuf[3159] = 256'h0c1991192718df16b4155a15bf138810d40bf1045b00dbfd9dfe0f0271064a09;
    decBuf[3160] = 256'hd70a400cae0c9f0e83122b174d1a021c861c1d1bd5197119cc191e1a941bd81b;
    decBuf[3161] = 256'ha31aaa18be153e12030e2a0b94082b077308650ade0c6710b113b0166819781a;
    decBuf[3162] = 256'hca1a5419001850163815d1151517e518191a511ab81917188e16c31413138a11;
    decBuf[3163] = 256'h590fb80c3f0aa408c3071709bf0bed0ec7125414cc14ce114e0e130a3a07bf07;
    decBuf[3164] = 256'h190a170dd00f2a108f0e590b5a086906c3065e08d409180a5f099709940cff12;
    decBuf[3165] = 256'hc020832e053b6446d24a7b49f040f43630286d1aeb0d8c022afb23f75bf8affb;
    decBuf[3166] = 256'hc304dd0a69107013b0102f09200209f803f459f075f185f8f0fe7106810dec13;
    decBuf[3167] = 256'h6c1b77206221e21e94190012f00a5a0685054706f70698072908a5070e09320b;
    decBuf[3168] = 256'h780f74130b166518ad19d81ae71bde1c931cc71b891be11aae1a6919f2165912;
    decBuf[3169] = 256'hb70ced087b051b06170ac00ee1114f11b00da2069701d7feacff760349086a0b;
    decBuf[3170] = 256'hd80a39070d029bfefbfdb0ff4602af034203500122fefefbd4fa2efbcafc14fd;
    decBuf[3171] = 256'h48fc1dfaa7f8ebf80efc7802b90a7d12911b3a1f8e228c21cc1e4c1c82181015;
    decBuf[3172] = 256'hef11f20d530a0807c00595043b048d046d052905f403fb0197fffcfd47fe9bff;
    decBuf[3173] = 256'hc701d2032605e804cf036a02df01b5015c005efe72fbb9f85ff843fb89ff8603;
    decBuf[3174] = 256'h13059b049c018ffc5bf686f038ebc6e7e5e59ae73aeb57f12cf77afc4d016e04;
    decBuf[3175] = 256'h4707e70a500c2c0a58042dfba2f24eef59f46ffe330df61ae62385251721111d;
    decBuf[3176] = 256'hf716330f270ae701ebf735f11beb37ec46f387fb4b035206920311fcfdf272ea;
    decBuf[3177] = 256'haee2a3dd0dd938d8fad86cdc0ee264ea28f233f7f4f91ef954f582f020ec8eeb;
    decBuf[3178] = 256'h1ced66f040f4d6f63ff8f7f63ef4c5f173f113f461f9b7017b09860e46117110;
    decBuf[3179] = 256'h2b0e5809f704d7ff04fb62f514f041eb61e939ece2f0c5f730fe5b02990188ff;
    decBuf[3180] = 256'ha5f83af264ec16e7a4e3c3e10ee093e00be12fe320e5e5e637e757e67be446e3;
    decBuf[3181] = 256'h7ee3e3e49be71aeb74ede1edf0ebc1e89ee63ae6b4e886ed7bf605ff91049305;
    decBuf[3182] = 256'hd30253fb3af0e4e57fdc65d611d30fd2cfd44fdc68e7b2f434015409b6105e0f;
    decBuf[3183] = 256'h260e9a088a0149f915edb6e16cd47dcbddc93fd1a4da81ea51f536fb00fd20f8;
    decBuf[3184] = 256'hbef008ead0e8b4e7b6e8a1e921ec67ee17ef77eec2ec19e877e229ddf6d620d1;
    decBuf[3185] = 256'h56cde4c903c895c82ccb67cfaad580dbcee001e72ceb7af04df56ef847fbc2fa;
    decBuf[3186] = 256'h68f86af5b1f2c1f34af776fce8ff8800affdf5f689f0b4ea66e5f4e192dddddb;
    decBuf[3187] = 256'h4fdac8daebdcf9e1cbe62deb29efc0f129f371f4d5f410f388ef5cea89e5e7df;
    decBuf[3188] = 256'h1ddcabd88ad5b1d21ad0b1ce44ce35d064d387d540d804dae8dc2fe172e7f3ee;
    decBuf[3189] = 256'h02f6c3f8edf7a7f5f7f497f570f80ffc88fc64fa90f4baeef0ea40ea20ecd6ed;
    decBuf[3190] = 256'h5aee10eb5be63ae3a8e23fe589e8d2e96ee9aae70ee61ae816ec59f284f646f7;
    decBuf[3191] = 256'h35f5d3f0d7ec49ebd1ea88e9d0e637e295dc47d797d6b8d9b4dd5de27ee510e6;
    decBuf[3192] = 256'h8be504e627e8a7ebe2efdef36cf5e4f552f6eef594f5f8f32df084ebe2e59ce3;
    decBuf[3193] = 256'h4ce4eee944f208fa14fffeff7efdb4f9e2f480f0cbee3dedc5ec7ceb8be97be8;
    decBuf[3194] = 256'h29e834ea30ee2df2ccf544f621f413ef41ea20e7b1e751eb8cef65f2fbf474f5;
    decBuf[3195] = 256'h06f5a3f448f4f6f316f33af18aef01ee02edbdeb42eaabe77ce47ee153e063e1;
    decBuf[3196] = 256'h35e6c9edd9f444fb6fff3100e10000ff4bfdbefb45fbd8fa74fa84fbd6fb21fc;
    decBuf[3197] = 256'hddfb23fb7bfaaefaacfc98ff510215041e03e8ff34fbd2f6d6f236efdcec03e9;
    decBuf[3198] = 256'h6ce622e3d9e104e37de506e941ed3ef1e6f588fbd6000a07350b7b0d2b0e8b0d;
    decBuf[3199] = 256'h400fd6114013ad13670f0008e7fc85f5cfee26eb42ec49ef09f289f44bf59bf4;
    decBuf[3200] = 256'hfaf38cf423f75efba10122092d0ec312981352111f0b49057f016eff0e00c301;
    decBuf[3201] = 256'h4802cf018700cefd0afc6ffaf9f8a5f779f56ef3a2f2d7f321f73dfd1303e509;
    decBuf[3202] = 256'h7b0e50149e19101db11dd81a1d14070af2fdd3f571eec9ef72f3fef809fec900;
    decBuf[3203] = 256'h9f01e503f605d707af0a3d0cb50c6d0b7b09d609cc0a420c860c510be808a806;
    decBuf[3204] = 256'hc80594064d071507180464ff02fb06f781f6eaf70efafffbc4fd0400cf037808;
    decBuf[3205] = 256'hda0cb20f4912b213b016f71a1720e9244b29002b73293725f41ec9153e0d0a01;
    decBuf[3206] = 256'hebf889f131f06af1bef4c0f580f856f918fa8afd6c04ad0c7114851d9f23f326;
    decBuf[3207] = 256'hf5270b278b24c1204f1ded1814167e132411000f0f0de009e206f004b506870b;
    decBuf[3208] = 256'h1b132a1ac01e961fcc1bf91657118d0d1b0a3a08cc085009aa0b840f2c144d17;
    decBuf[3209] = 256'h261aa2193918f0168d1632163b150512510dae076805da08bd0ffe17fa210126;
    decBuf[3210] = 256'hc82474216d1e831d0320cd239f2840296726b520671b3415b4126e105d0e7c0c;
    decBuf[3211] = 256'ha3091f09a608ef09520af80914075b044c03d406e20dfb184526a12b412dc72b;
    decBuf[3212] = 256'h6222d7194b1449135e12de14a015f01450147711f2105c125a15da18061ed822;
    decBuf[3213] = 256'hfa25af272126c723ee1f451be416e7125110f70dd40ba90a040b430d0f11af14;
    decBuf[3214] = 256'h081751187b19401b6d1fb025312d3c32d236fc352a2fea26b61a570f01054afe;
    decBuf[3215] = 256'h12fd66007607b70f7b17861c461fc61c801a0e172d157813fd1375147317811c;
    decBuf[3216] = 256'hb422352a402f0032802f322a3d21b318271320100b11e011261476139511990d;
    decBuf[3217] = 256'hf909ae0666059006740a2510f716631d38230a2a76304b36153ac63a253a0635;
    decBuf[3218] = 256'h112ca51e2212c3066dfc66f89ef92aff3a067b0e071409151e1449137f0f0d0c;
    decBuf[3219] = 256'hec0813068f05d908440f301b8f26f12d482f9f2ba3213e182412980c960b800c;
    decBuf[3220] = 256'h560d180ec80e680ffa0f7f10160f830fae102713f9172c1e572219230821661b;
    decBuf[3221] = 256'h1816a612c5107a121a1692164a15ca11ad0b8207b80369048a07860b1d0e950e;
    decBuf[3222] = 256'h720cf208c603540033fd5afad6f94efa97fba400380851139b201d2d3d35b736;
    decBuf[3223] = 256'hb032252af11d92123c0886016cfb18f811f551f2d1f49bf82f0044093f14a11b;
    decBuf[3224] = 256'h572271288d298b28a0277528b327a22581223e1cbd14a90b1f035bfb54f83ff9;
    decBuf[3225] = 256'h69f82bf9dcf9baf6e2f339ef18ec63eaf0eb2bf06ff69aff24082012861b2f1f;
    decBuf[3226] = 256'h4b20491f5e1e331a6916f712d60ffd0c670afe086b095d0b210d180ea20ca608;
    decBuf[3227] = 256'h1c0091f795ed8ee9c7ea53f067f9f201b609bc0c7d0fa70e690f580df6089001;
    decBuf[3228] = 256'h7bf880ed12e9bae7d4edd0f73601c009dc0ad5076a0195fb47f696f577f773fb;
    decBuf[3229] = 256'h25017306450b260d710bbf05edfeadf6e9eee2ebf7ea77ed41f175f79ffb69ff;
    decBuf[3230] = 256'h1a007affc4fd25fadaf6b7f41af5dff667faa3fe9f023f06b7062407fa053504;
    decBuf[3231] = 256'hf601bffe30f95ef2f3eb1de6cfe01fe040e360e8f4ef04f76ffdefff2dffbbfb;
    decBuf[3232] = 256'h9af8e5f660f6d8f621f84bf9a6f941fbb7fc83fdc1fda8fc11fa98f7a1f617f8;
    decBuf[3233] = 256'h03fbbbfd16fed6fb0af86bf420f1d7efadee33ec06e8e6e2d5e076e195e6c9ec;
    decBuf[3234] = 256'h9ef268f619f778f6e7f57df8c8fbebfdc1fc73f7a1f061e80de50fe6cfe84feb;
    decBuf[3235] = 256'h95ed46eea5ed5beffaf245f68df763f6caf128ec5ee80ee9efeaebee79f02eed;
    decBuf[3236] = 256'h9fe7cde061dae1d727da38dc5adf56e3ece519ebadf2bcf952fed20008fdd5f6;
    decBuf[3237] = 256'h55ef49ea89e75ee8a4ea16eef7efacf131f2a9f261f11aedd7e657df4bda36db;
    decBuf[3238] = 256'h61df33e6c9ea49ed87ec15e934e7c6e75cea98eeb8f38af8ecfcc5ff5b02d402;
    decBuf[3239] = 256'h8b01b7fb8bf290e72ee078d9cfd5b3d4acd116cd96c58bc0a0bfcbc329cf07e1;
    decBuf[3240] = 256'haef1d000b606120cb20d2c0fd50d9c0c10070502c4f938f428ed68ea3de6f7e3;
    decBuf[3241] = 256'h85e0a5de13de97de01e049e174e219e2c7e17ce1b0e072e05adf5bded0dd4ede;
    decBuf[3242] = 256'h8ee05fe532ea53ed08ef7bed12ecc9ea9fe944e9f2e87ce718e5d9e223e397e6;
    decBuf[3243] = 256'hb4ec35f444fbdaff05ff3bfb07f532ef68ebf6e7d5e4d8e039ddeed9cbd767d7;
    decBuf[3244] = 256'h77d8b6da2cdc08de3ddfc6e091e241e45ae5bfe6bde821eb4eef4af3eaf653f8;
    decBuf[3245] = 256'h0af752f423f100ef0eedffeb1be90de4dadd04d8bed5cfd772dd44e4d9e8afe9;
    decBuf[3246] = 256'hede8dce63be6f1e799ecbaef4cf0bfee65ec41eaa5ea1eeda7f0f2f315f6b2f5;
    decBuf[3247] = 256'h57f560f4ebf20ff167ee39eb3ae89ee817ebe9ef1cf647fa09fb97f7f5f1a7ec;
    decBuf[3248] = 256'h35e995e84aeae1ec4aeeb7eec6ec4cea68e777e567e45ee5d4e6b0e860ea79eb;
    decBuf[3249] = 256'h46eb01ea83e9f6e901eca2ee66f0b8f0adee39ebeee7a6e697e8c6eb9fef36f2;
    decBuf[3250] = 256'h9ff30df470f480f564f8e3fb2eff7600da0015ff8dfb51f70ef138eb66e4a6e1;
    decBuf[3251] = 256'h26df6ce17de39ee654e8e1e94aeb6eededf029f525f9bbfb15fe83fee6fe8cfe;
    decBuf[3252] = 256'h03fbd7f543ee33e773e448e596ea8bf316fc6aff67fea7fb7cf7b2f340f060ee;
    decBuf[3253] = 256'hceed37ebdee870e8d4e898ead8ec23ed57ec22eb5aeb57eee6f3b8fa2401a403;
    decBuf[3254] = 256'h660455027400bffe43ffbcffdf01d1039505d507e009240af8072d047bfea9f7;
    decBuf[3255] = 256'h3ef168eb9ee7cce2ebe059e0e7e113e746ed71f68bfcdfffe100f7ffcc008e01;
    decBuf[3256] = 256'h00056209170b920a57065b02cd0046011f05c809a80bf3094b05a8ff62fdb2fc;
    decBuf[3257] = 256'h52fde4fd56fc2af758f236ef0ff2caf8e00296093f0d230c1c095c0687054906;
    decBuf[3258] = 256'hf90659065d02abfc5df7ebf34bf300f5a0f8dbfcd7006502ce036103a8002ffe;
    decBuf[3259] = 256'ha6fa4cf8def797fa7afe2c047a09ec0ccd0e5e0fda0e710d4d0bce07920373fe;
    decBuf[3260] = 256'ha0f93ef5acf431f58bf764fbfbfd45016903e806240b67113d17071bb71b9618;
    decBuf[3261] = 256'h9a14e80e9a092806c601eefe60fde8fc30feb001eb05e7097e0cf60cae0bbc09;
    decBuf[3262] = 256'hf80701072106dd051b06a307a00a30107e15f01850180c12e108e6fd84f62cf5;
    decBuf[3263] = 256'h65f629fe3805ce094e0c100dc10d200dd60e6c11b7149018301c8a1ed21f6f1f;
    decBuf[3264] = 256'h401c8c172a130a0e980ab708df054803ee00a6ffd00069054c0cb712371a3e1d;
    decBuf[3265] = 256'h291e531d911c801a5f173f126d0dca07840535065609760e48132915bb153615;
    decBuf[3266] = 256'hbe14e116281b011e851e2b1c771715133c10c1102a1272134812190f8a09c005;
    decBuf[3267] = 256'h7006d20a151196189c1b871c071ac117b01510155a13cd11820ea90a12089a07;
    decBuf[3268] = 256'he2089b0bc90eed10de125815e1182b1c741dd71d5e1bd5177b150e1538164817;
    decBuf[3269] = 256'hf516bf13300e5e07c802f301bd058f0a7211dd175d1a1f1b6f1acf19841b231f;
    decBuf[3270] = 256'h6e224826cc2663258921e11cc019e7166216db164817ac175117ff161f165315;
    decBuf[3271] = 256'h9a1411137a10000e770a1e08d5063907b209840e18162c1fb7277b2f82324235;
    decBuf[3272] = 256'hc232f82e252ac325c7211f1dbd189d132b104a0edc0e7311ae1587181d1b961b;
    decBuf[3273] = 256'h4d1a2319a9166914c9119a0e770c130c6e0c520f98139517341b7f1ea2209422;
    decBuf[3274] = 256'ha323ad22a1202d1d01188f14af124013ce144615d9147514d0140f17711bd424;
    decBuf[3275] = 256'h8b2b342f5030492dde265e241822672107225220bc1d9018bd139c10e60e620e;
    decBuf[3276] = 256'hcb0f3910d50fc60e2a0d4a0c7e0bbc0bd40c6b0f9a129815511860196a185e16;
    decBuf[3277] = 256'hfa130413e413c0157017891856186e174417b717f1186c1a9f1a711a9b1a5b1b;
    decBuf[3278] = 256'h661dc7212926de275026242190197c10d30c7f09810a170f42130c171d19fe1a;
    decBuf[3279] = 256'hd61d5b1ec41f0c21a920991f5a1db91a8a1767157513b11116100a0ea60b6709;
    decBuf[3280] = 256'h8608da09820cb00fd411fe123a11fa0eef0c9b0b540cdd0d0e10191205158518;
    decBuf[3281] = 256'hc01ce0211328e92d2f30df30be2d7b27fa1fe6165b0e5f04a9fd8ff73bf439f3;
    decBuf[3282] = 256'hcff7a4fdfa05f60fad16e5170119fa153a13ba10f80fe70d060c2d098e053403;
    decBuf[3283] = 256'hc602f1036a064f09400bba0df90f051259139f12a610ba0d3b0ad2083f096a0a;
    decBuf[3284] = 256'hc40acd092d074903b3002b014e0395076e0afb0b830b5f09350825077807c207;
    decBuf[3285] = 256'hf60646056c02edfe93fc4bfbe7faf7fbdbfe5a02a505a308ce09280ad6098b09;
    decBuf[3286] = 256'h4709010a390aa0095b088907c906ec068a073307ac05620245fc1af8d4f584f6;
    decBuf[3287] = 256'h65f861fcf8fe52019a027001abff22fcd8f8d9f5e8f3d8f22bf3a0f404f7e9f9;
    decBuf[3288] = 256'h2ffe4f032108830c380eb40d8808f400dff755ef91e786e29be170e232e3a4e6;
    decBuf[3289] = 256'h06eb02efa2f2ecf5ebf831fd2d01d605f708890904099b079d04e4012000ceff;
    decBuf[3290] = 256'h83ff2ffe88fb0ef92af6fff4a5f49cf57cf6c0f694f433f050e90fe183db7dd8;
    decBuf[3291] = 256'hbcd592d65cda0cdbeddc7fdd0cdf57e2e6e734ed07f2a7f215f27fef16ee5eef;
    decBuf[3292] = 256'h17f245f58ef663f580f1e0ed86ebf4ebacee45f3a7f77ffa04fb9bf99cf6e4f3;
    decBuf[3293] = 256'hb5f0b7edc5eb4ce967e676e4b1e25fe26ae466e8aaee7ff4cdf9defbfef9def4;
    decBuf[3294] = 256'habeed5e887e376e1d6e067e1dadf71de4ddc23db13dac1d90cdac8d98ad952d9;
    decBuf[3295] = 256'h85d983db6fdeb5e2d5e7a8ec0af1e2f367f4eef3cbf112ef2feb98e82fe7e7e5;
    decBuf[3296] = 256'h4ae65ae708e7e8e72ce861e95aeb46ee37f047f107ef3beb93e631e235dea7dc;
    decBuf[3297] = 256'h3edbf6d976d62bd352cfc4cd2ecf2cd23ad70cdc2ddfbfdf3bdfe1dcbdda05d8;
    decBuf[3298] = 256'h8bd595d44ad416d5c6d62fd914dc93dfdee292e7f4ebf0ef99f4baf76ff9fdfa;
    decBuf[3299] = 256'h94f94bf8ccf490f071eb3de5bdddadd642d0c2cd7ccb8dcdefd10ed7e1db02df;
    decBuf[3300] = 256'hb7e033e0d9ddb6db36d8dcd5b9d355d3b0d302d478d5dcd7c0da06df03e3abe7;
    decBuf[3301] = 256'h8ce91eea87e72de50ae36de3e7e5cbe884ebdeebe7ea47e818e5f5e2cae170e1;
    decBuf[3302] = 256'h1de168e1ace1d8e30ee7e8ea90ef71f1dff052ef16ebf6e585e263df8bdcf4d9;
    decBuf[3303] = 256'h9ad752d6eed549d69bd67bd7bfd7f4d8cedbdbe06fe883f19df7f1faeff92ff7;
    decBuf[3304] = 256'h04f33aefc8eba7e8f2e65be410e1eddefbdcecdbe3dc58de44e18be5abeadef0;
    decBuf[3305] = 256'hb4f67efaf0fd4ffd9afb0dfac2f6c3f37def81ebc6e430e006dcc0d9d1dbb1dd;
    decBuf[3306] = 256'h43dec8de4fdee2dd45debfe091e563ea05f04bf25df4fdf48ff513f68bf6f9f6;
    decBuf[3307] = 256'h07f5d9f1ffed60eaf7e8aee7d9e807ec06ef85f2dff428f6c4f51ff6ccf5adf6;
    decBuf[3308] = 256'h89f8bdf966facdf972f7e9f39ff07bee18ee72ee69ef49f07defcded63eb7fe8;
    decBuf[3309] = 256'h8ee67ee519e7bae953eeb4f2b1f650fa9bfdbeffb001bf02b6030104250202ff;
    decBuf[3310] = 256'h29fb92f829f796f7faf79ff7a9f672f399eff9eb90ead9eb91eedff3a9f71bfb;
    decBuf[3311] = 256'hfbfc8dfd09fd72fe4b02f406560b0b0d860c3c098704e5fe9ffc8efa2efb9cfa;
    decBuf[3312] = 256'h0ff9c4f5ebf14beee2ec75ec9fedafee4af0ebf283f725fd7302a7087c0e4612;
    decBuf[3313] = 256'hf712971305136f10330c1407e000b5fcebf83bf8dbf8b4fb4afe860282062b0b;
    decBuf[3314] = 256'h4c0e0110740e380a18054600e4fbe8f751f5f7f2d4f0a9ef4fef33f241f774fd;
    decBuf[3315] = 256'h9f01e50335035401c2003e00c5ff3300cfff75ff7efec9fe1d00cd01c6039204;
    decBuf[3316] = 256'h4b058305e8064309830b8e0d5a0e1d0e740d410d700d9a0d400c890942054601;
    decBuf[3317] = 256'ha6fd2efd9cfd8dff520191035d07060ca8117a18101d901f5220a11f011f281c;
    decBuf[3318] = 256'h92194716b8106a0b9706760308049505ef075c083207b8041d0393048f08d20e;
    decBuf[3319] = 256'ha8147218221941178c15081571169418861a2b1aec172014770f160b3d08af06;
    decBuf[3320] = 256'h280770089b095f0bfa0c700e3c0ff50f2e106110a511201351155d17b118611a;
    decBuf[3321] = 256'hea1b811eaf21ae2466270c2727241a1fe7181113470fd50bf4093f08a9055e02;
    decBuf[3322] = 256'h15017901a704370a8d12511a61212124f624b022de1dbc1ae4175616cf161718;
    decBuf[3323] = 256'h4219511aa31ac3196f18bf16c614ea12c70fc80c4909ef0682067308c10d1716;
    decBuf[3324] = 256'hdb1def26982aec2dea2cff2b2a2b682a182bb82b262b902836265d22c61f7b1c;
    decBuf[3325] = 256'h331bcf1a2a1bc51c661f4923e92643298b2aef2a75289125d922aa1f621ec51e;
    decBuf[3326] = 256'h8a206e23262636278827122646257b2655299b2d97312e34a63439340e339530;
    decBuf[3327] = 256'h9e2f282e4c2c932b5b2b5a2c582e3430e4316d33d23474364d39cd3c273f4a41;
    decBuf[3328] = 256'h2040f13cf339733628332a30712d8e29ee2595234c223e242128c12b0b2f0a32;
    decBuf[3329] = 256'h6d327d3318352337973ae23de040d242e1434642a53fc23b2238e733eb2f422b;
    decBuf[3330] = 256'h21284825bb235222e42148225723f224fe26ea29302e5033833904410f46fa46;
    decBuf[3331] = 256'h2446de436c404b3db93c353ccc3acd37c032ed2d8b29b3263727af27f8285b29;
    decBuf[3332] = 256'h0129f8292e2de23185374f3b9e3a7d373a310f28841ff819ed142d125711110f;
    decBuf[3333] = 256'hc20f6210f4108a13e415e218d41a4d1de91ec91f0d20541fcb1dce1a19167710;
    decBuf[3334] = 256'h290b56063503800104026e039105830728078d05ec0209ff72fc09fb9bfac6fb;
    decBuf[3335] = 256'h8afd81fe36fe7afeb8fed1ff360191032c050c06c8050f05f6039102f000f7fe;
    decBuf[3336] = 256'h1bfde6fb5dfac4f9dcf8b9f682f384f092eeedee1af381fa9101fc077c0aba09;
    decBuf[3337] = 256'he70445fff7f9c4f399ef4bead9e6f8e467e4f4e54ee871ea2aeda3efe3f1c3f2;
    decBuf[3338] = 256'h07f3caf292f25ff2eaf265f4fcf62afa29fd53fe44fdbbf980f583f1edee65ef;
    decBuf[3339] = 256'h89f1cff5ccf962fceafbebf817f3ece9d2e30edc02d76dd297d1d5d086d166d3;
    decBuf[3340] = 256'h63d70bdceee259e92feff9f26bf68cf91efaa2fa48f86ff4bdeeebe756e32bdf;
    decBuf[3341] = 256'h69de19df79de0bdf74dc1adad2d86ed833da60de5ce2fce556e8c3e8d2e60de5;
    decBuf[3342] = 256'h29e2a9de6eda72d6c9d1a8cecfcb4bcbd2ca1bcc7ecc8ecd85ce90d07cd334d6;
    decBuf[3343] = 256'h44d7f2d651d422d1ffced4cde4ce24d12fd373d335d3fdd262d41ad727dc99df;
    decBuf[3344] = 256'h39e03ddc94d7f2d128ce17ccb7cc26cc98ca20ca68cbafcf15d72ae0b4e878f0;
    decBuf[3345] = 256'h7bf1baee8fea41e50edf8ed77ed03dc8b1c2aabfc0beeabd28bd17bb36b981b7;
    decBuf[3346] = 256'h18ba53be96c46cca36cee6ce46ceb4cd42cf8cd241d762da5edef5e05ee2a7e3;
    decBuf[3347] = 256'h98e5f3e557e421e16ddc0bd80fd478d1f0d139d3f1d5d5d96bdcd5dd42de18dd;
    decBuf[3348] = 256'he9d9a1d804d97edb4fe022e543e8f8e974e90be89de701e8c5e9bcea71eaa5e9;
    decBuf[3349] = 256'h68e910ea0ded9cf2eaf75cfb3dfdabfc15faacf83ef830fa13fec5031b0c1716;
    decBuf[3350] = 256'h2b224b2aad31b4355d3941383a354f34cf310d311e33be3374350a38643a883c;
    decBuf[3351] = 256'h793ef3407b44a7497a4edc52d8566658ed578057e3573e58d9594f5b935b5e5a;
    decBuf[3352] = 256'hf557105558529350f84eed4c894aa547ec447342c542d044cc48ec4dbe52e055;
    decBuf[3353] = 256'h95571057c653ec4f564dfc4ab34950498b475e433e3e4a35bf2cfb24e71bcd15;
    decBuf[3354] = 256'h7912720f5d103211f411a51204124f10c20e490edc0d780d4a0a9505b2fe72f6;
    decBuf[3355] = 256'he6f0d6e940e56bdfa1dbced66cd2dad168d3c2d5c0d8ebd971d744d324ce52c9;
    decBuf[3356] = 256'hf0c43bc3adc153bf7abbe3b889b641b5a4b5ffb508b5fdb211b01fae10adabae;
    decBuf[3357] = 256'h4cb17ab49eb6c8b7d8b873bae9bb4dbee8bf9dbfc1bd23ba84b639b3ccb2bdb4;
    decBuf[3358] = 256'hecb7c5bb5cbea6c1cac3bbc535c8bdcb17ce16d107d3ccd4c3d5a3d6f7d71adb;
    decBuf[3359] = 256'hf3de93e2cee6caea58ecb2eed5f000f25af251f306f3d2f307f570f7f9fa2500;
    decBuf[3360] = 256'h9703b80691091e0b970b290b710842051f03f401b90342077d0b560ed10d770b;
    decBuf[3361] = 256'h9e070705ad021b03b702a8011ffef3f8c0f295ee4fec9eeb3fecd0ec55edeceb;
    decBuf[3362] = 256'h7eebc6e84ce60de46ce1f2dea0de80dfd4e0f7e31be60ce867e8cbe695e3bcdf;
    decBuf[3363] = 256'h13dbb1d6b5d216cfbccc4ecc24cbc9ca77ca01c915c65dc3e3c048bf93bfe7c0;
    decBuf[3364] = 256'h97c200c59cc6e6c6b2c7f0c798c831c903c934c711c481beafb744b119add3aa;
    decBuf[3365] = 256'h84ab24acfdae93b1fcb220b566b986be1ac62acd95d3c0d706da56d934d65cd3;
    decBuf[3366] = 256'haacd5cc829c2a8baa2b7b7b6e2baacbedfc45fc7a5c956caf6cacfcd77d219d8;
    decBuf[3367] = 256'he3db55dff6df87e015e28de2fbe2d0e138dd55d6eacf14cacec71ec7bec773c9;
    decBuf[3368] = 256'hf8c961cba9cc29d055d588db5ee130e8c6ec46ef08f0f7ed95e975e4e1dcd1d5;
    decBuf[3369] = 256'h66cfe6c7dac245be1abad4b7c3b5a1b282adafa84da451a0cd9f26a225a5a4a8;
    decBuf[3370] = 256'hefab13aecbb019b66fbea3ca41d904e71af73c06ff13ee1c0e257c29d32a9b29;
    decBuf[3371] = 256'h0f240821731cf2193019421ba31fc3249629f72df4318133fa336734cb342535;
    decBuf[3372] = 256'h2e342332272e072995253626322af531b939ce42e8483c4c424fae55835bd963;
    decBuf[3373] = 256'h6569676a7d69fd66b7640664a6645c66e066496892694a6c2e70d674797abf7c;
    decBuf[3374] = 256'hd07e2f7e9e7d107ca77a8478cb755273b6716c71d0735877b279d67b727b637a;
    decBuf[3375] = 256'h107ac6791a7b4e7c877cbc7a1d777572d36c09693664d45f91591152fc487240;
    decBuf[3376] = 256'hae38a2330d2f8d2cc3285125ef20f31c41177713a50e830b8707e8038e014500;
    decBuf[3377] = 256'h70019e0478080e0b680d450bc5078a0346fd71f723f28fea7ae161db9dd38dcc;
    decBuf[3378] = 256'hcdc94cc706c5b7c557c6e9c67fc9cacca3d043d47ed87bdc1ae055e42ee7ceea;
    decBuf[3379] = 256'h46ebd9eae7e86ee677e5c2e5aee82dec68f065f404f86df9b6fae0fb3bfcd6fd;
    decBuf[3380] = 256'h21fe65fe1effa700a4033309810e1616251d91236629b42ee834bd3a0b403f46;
    decBuf[3381] = 256'h144ce6525159275ff9658f6a0f6dd97089712a72bb723772ce706070c470d371;
    decBuf[3382] = 256'h6e734f7493745e736571896fd06e086f077035700e6f686d4f6c1c6cbe6d9770;
    decBuf[3383] = 256'h8972e372ff6ff26abe64e95ea35cf25b525bc05a455bdc5993586957ef540b52;
    decBuf[3384] = 256'h8b4e5f492c43563d083836331430182c6726951f2919a911a20ee20bb70cf50b;
    decBuf[3385] = 256'h450b64096805b7ff69fa96f534f17feff1eda7ea83e804e5c8e0ccdc2dd9e2d5;
    decBuf[3386] = 256'hbfd3cdd154cfb8cd18cb34c795c359bf5dbbbdb764b5f6b4e8b6acb8ecbaccbb;
    decBuf[3387] = 256'h98bcdfbb17bcb0bcf5bdc4bf7dc0b5c01cc07bbe62bd63bcd8bb02bc29bc91bc;
    decBuf[3388] = 256'h6fbdabbe7ac022c305c7a5cae0ce00d472d752d908db7ad902d9b9d71dd82cd9;
    decBuf[3389] = 256'hc7da3ddc91ddc6defedefddffbe16fe5abe9caee3cf29ef677f9fbf992f825f8;
    decBuf[3390] = 256'hfaf6a0f63bf846fabafd050128035304f803b80182fea9fa09f7bff376f24cf1;
    decBuf[3391] = 256'hf1f0faef85ee99ebe0e867e6cbe4ebe31fe366e2dde0acdea1dcd5db12dc2bdd;
    decBuf[3392] = 256'h5cdfd2e08ee059dff0dc67d92cd52fd187cc25c829c492c129c0bcbf1fc02fc1;
    decBuf[3393] = 256'h25c270c23cc3f5c32ec4c7c4dfc364c299c06dbeccbb08ba6cb8f7b61bb56ab3;
    decBuf[3394] = 256'h71b1a5b0ecafb4af4db0d8b0ffb158b3fab482b64db807b93fb972b9d0b7d7b5;
    decBuf[3395] = 256'hebb26caf30ab58a8caa652a675a8f5ab4fae97af34af6fad2fabbaa9eea8b0a8;
    decBuf[3396] = 256'h08a809a70aa5a6a267a05b9ef79bb8998196a892088f9f8de88e2e934e98e29f;
    decBuf[3397] = 256'hf2a65dad33b305ba46c242cca7d513e396ef34fe0908f810d815461a9d1bd61c;
    decBuf[3398] = 256'hf21df41e8a235f29292d3b2f1b318a30f32da82af4255220041b311610137e12;
    decBuf[3399] = 256'h03136c144518ee1c90226229a33167397640b7487b508b57f65dcc631a692b6b;
    decBuf[3400] = 256'h8b6ab2672466cb6382621f627962cb6241642d67ad6ae86ee4728476ce79f27b;
    decBuf[3401] = 256'h1c7d777d257d447c5879127516716d6c8c6a1e6bac6cf66fd0736676cf776277;
    decBuf[3402] = 256'hfe768574ea7249701a6d41699864b65d4a57ca4fba484f42cf3abf33292f5329;
    decBuf[3403] = 256'h05249420321c12173f125d0bf10471fd61f6f6efcbeb7de6abe149dd70dae3d8;
    decBuf[3404] = 256'h79d7e7d711d9d6da71dc51dda5dedadf12e079df7bdd07dadbd408d066ca18c5;
    decBuf[3405] = 256'h46c0e4bbc4b652b331b07caeeeac85ab18ab7bab40ad24b0a3b3eeb6c7ba5ebd;
    decBuf[3406] = 256'hc7beebc0a3c387c72fcc91d08dd424d77dd9a1db92dd57dff2e068e2bce36ce5;
    decBuf[3407] = 256'hd6e715ea4ced6fef28f256f555f8d4fb0f000c04b408160d1211b214de19501d;
    decBuf[3408] = 256'hb1218a2421279927e2284529552a942c60300935ab3a7d411346e84bb24f2453;
    decBuf[3409] = 256'h45561e59ac5a335aeb58f9563555f552155249518f50e74fe84e474dbe4bf349;
    decBuf[3410] = 256'hbe488648b94844496b4a2b4b4e4bef4aec496c4807476645dd43ac41763e9c3a;
    decBuf[3411] = 256'hfd36c232c52e2f2cd529fb255321b11b63169011ee0b2408b2049101b8fe2afd;
    decBuf[3412] = 256'hd1fa88f9ecf991f988fad3fa8ffad5f94cf81bf67bf34cf029ee70ebace96ce7;
    decBuf[3413] = 256'hcbe49de1c3dd24dae8d510d382d119d086d023d07dd02bd0e0cf9ccfdacff3d0;
    decBuf[3414] = 256'h58d2f9d312d5abd5c3d49cd3f6d16dd008cfc3cd9dcc90cb10ca11c929c8ffc7;
    decBuf[3415] = 256'h72c8f2c989ccb8cf91d328d672d996dbf9db09ddffdd75dfc9e0fee136e2d1e0;
    decBuf[3416] = 256'hd3de5fdb14d8f1d5c6d46cd4bed409d5d5d50ad792d85dda05dd7edfbee1c9e3;
    decBuf[3417] = 256'h1de552e64be89fe9d4ea5decf6ecdeed08ee48ed54ec37ebdee999e81ee753e5;
    decBuf[3418] = 256'h27e31ce1b8de78dc02db26d96dd855d7f0d508d535d40fd432d4d0d426d5a9d5;
    decBuf[3419] = 256'h1fd68bd615d7d9d7f4d74dd709d651d399d01fcee0cb3fc97ac784c639c605c7;
    decBuf[3420] = 256'h31c9d1cb00cf48d0acd09ccf01ceb6cdfacdabcf14d2f8d4ead6aed800d94bd9;
    decBuf[3421] = 256'h07d9c9d8b1d74cd607d5e4d2d8d074ce35ccbfca7bcab9ca41cc72ce7ed0e2d2;
    decBuf[3422] = 256'h21d52dd791d975dc66de2be07de09ddfc1dd95db8ad9ced987da10dca9dc1edc;
    decBuf[3423] = 256'ha6d9c3d523d2bad04cd03ed26cd56bd8eadb35df0fe3aee6f9e941eb6cec5ceb;
    decBuf[3424] = 256'hc1e94be8f7e635e7dde710e828e705e5cfe1d0dedfdc1adbc8da13dbdfdb1cdc;
    decBuf[3425] = 256'he4dbe5da44d94bd76fd5b5d40dd4dad308d4ded31ed3e5d169d09ece6acd71cb;
    decBuf[3426] = 256'h1dca63c9bbc822c83ac76bc5bac332c233c177c2efc43dca9bd5fae050eb64f7;
    decBuf[3427] = 256'h84ffe6069c0db61342194d1e0d218d234f24c127a229c22e9433b636b23a3f3c;
    decBuf[3428] = 256'hc73b7e3a54398f3799364e360a364836f03657362936fb36a138eb3b0842de47;
    decBuf[3429] = 256'h2c4d9e50bf5374550b58655a885c415fba61fa6305666968f26b3c6f60711874;
    decBuf[3430] = 256'h92762d78387a147cc57ddd7e447e467ce27959760f731070916c466923673165;
    decBuf[3431] = 256'h2264746429646d64b4639b623661955f0c5ea75c625b3c5ae2589e577a554452;
    decBuf[3432] = 256'h454f384a65450341e43b72389136b8332b32d12fd22c1a2aeb263722d51dd919;
    decBuf[3433] = 256'h3015cf108b0ab604e4fd78f7f8efedea57e6d7e391e180dfe0de4edec0dc66da;
    decBuf[3434] = 256'h43d88ad511d376d100d034cf7bce43ceaacd1ecd4cccf2ca51c938c839c752c6;
    decBuf[3435] = 256'h27c69bc6bdc6ddc6fac6abc635c6c9c58ec50bc6ffc60ac9aacbd9cefcd027d2;
    decBuf[3436] = 256'h36d32dd40dd5e9d691d9bfdc99e041e562e85fecf5ee4ff173f364f5def766fb;
    decBuf[3437] = 256'h9200c6069b0ce911bc165e1c28209a23bb267128fe29582cc62cb72e7c301732;
    decBuf[3438] = 256'h2234fe35ae37a739933c13405e433747d74a304d544f7e508e5185526553a953;
    decBuf[3439] = 256'hf052475248516050e24fbc4fdf4fbf4f694fb24edc4d134d904c194cd94bd94a;
    decBuf[3440] = 256'h14496d468942ea3eae3ab2361333aa31862f952dd02bec28332605232b1f951c;
    decBuf[3441] = 256'h4a194c1693131a11350e440cca092f08b90675063806e006df070d088f07e905;
    decBuf[3442] = 256'h9f0264fe44f9d2f570f1bbef1cecb2eab4e7c2e5b3e4bce3dce288e153e05ade;
    decBuf[3443] = 256'h06dd56db1edb51dbdcdbaedc22dd44dd64dd47ddf9dcb2dc46dce3dbf5db67dc;
    decBuf[3444] = 256'h44dd1fdf83e11ee394e4e8e5a1e6d9e60ce73ae70de8cde807ea2aec36ee9af0;
    decBuf[3445] = 256'hd9f24ff493f455f41df450f4dbf4abf6d7f80dfc0bffc401880324056e052a05;
    decBuf[3446] = 256'h6805a0059f06e4070b09170a0b0be90b250d4c0e590fc10fa20f120f5b0e140e;
    decBuf[3447] = 256'hd30d980d3f0d4b0c570bf80a4e0b390c950d7d0eff0d0c0c20096706ee035202;
    decBuf[3448] = 256'hdd0099005b002300f0ff08ff35fe29fdeffb1cfba9fa12fbb0fb40fc89fb24fa;
    decBuf[3449] = 256'h27f74ef3aeef64ec40ea88e7c3e528e448e37ce2bae2f2e2bfe2d7e15ce091de;
    decBuf[3450] = 256'he0dc58db59da14d999d7ced5a2d32cd270d2aed237d49cd584d602d729d791d7;
    decBuf[3451] = 256'h2fd8bfd80dd925d910d938d86ed7b8d641d62bd68dd62ed7f1d710d983d960d9;
    decBuf[3452] = 256'h02d9c5d74ad64bd563d439d446d53ad657d763d857d9f5d9bfda76db4bdc4edd;
    decBuf[3453] = 256'hb7ddd6ddbadd9adc8edbdfda41dad1daf0db96dd8fdf6be1a0e249e316e32ee2;
    decBuf[3454] = 256'hafe13ce15fe17fe10ee2f4e17ee1bbe09cdfdcde2ddeceddb2dd98ddf1dc03dc;
    decBuf[3455] = 256'h68da6fd80bd6cbd356d202d1c4d01cd083cf9bce74cd1acc79caf0c825c7f0c5;
    decBuf[3456] = 256'hd8c4d9c3aac329c4e9c423c69ec703c901cb65cd49d090d4afd982de65e5d0eb;
    decBuf[3457] = 256'ha6f178f80dfd380102051307f4088609130b7c0ca00e5811d21312161d18e918;
    decBuf[3458] = 256'h27197e1819171b15b7121c11a60f620f1b1034119912f414d817911abf1d9921;
    decBuf[3459] = 256'h382574294c2cec2f36335a351238413b3f3ef840db447b48b64cb35052548d58;
    decBuf[3460] = 256'h8a5c29607463bc64e7658c659664f56130604c5d945a1a58da55cf536b51d04f;
    decBuf[3461] = 256'h2f4db64ad14719459f426040ea3e963de63bec391038e5356f349332ec2f722d;
    decBuf[3462] = 256'he929ae25d5223f20e51d9c1cab1a9b195c17bb142210c10b7d05fdfdedf682f0;
    decBuf[3463] = 256'h02e9f6e361df36db6cd75bd539d284d0eecd94cb95c8ddc5aec28bc099bed5bc;
    decBuf[3464] = 256'h3abbc4b970b8c0b637b538b450b329b2d0b02eafa5ad40acb5ab34ac8dade8af;
    decBuf[3465] = 256'h28b233b487b540b678b6dfb554b52ab550b5b9b596b699b747b864b9bdba5fbc;
    decBuf[3466] = 256'hc8be08c1a9c36dc564c644c798c8c4cafacdafd210d70ddbacdee8e2e4e68ceb;
    decBuf[3467] = 256'h2ff1f9f4cbf92dfe2902c905040a000ebb14261bfc20ce27632ce42eae32bf34;
    decBuf[3468] = 256'h9f365538e2394b3bb93b1c3cc23b143cf43cd03e8140994132426142e2416f41;
    decBuf[3469] = 256'hd84176422544d5455e47c348084a2f4b884ccd4d9f4ec64e174e7c4c134ad347;
    decBuf[3470] = 256'h32456e43d341f2409e3f6a3ee13ce23b403a4738e3355a322e2d5c28fa23da1e;
    decBuf[3471] = 256'h081aa615cd123710ec0cc80a9e09240789057e03a201f2ff69fe6afd82fc5bfb;
    decBuf[3472] = 256'hb5f92cf8c7f682f507f408f367f1deefadeda2eb3ee9a3e797e543e40fe386e1;
    decBuf[3473] = 256'hede005e0deded1dd97dc1cdbb7d973d84cd78cd669d607d7d0d787d82ed99ad9;
    decBuf[3474] = 256'h5fd929d9b7d850d80dd8b8d755d713d71fd782d74ad8fad925dc31de95e08be1;
    decBuf[3475] = 256'h01e355e405e6fee7dae98beba3ecd6eca8ecd2ec45edc5eef6f097f35bf59bf7;
    decBuf[3476] = 256'h7bf847f900fa38fa37fb1ffc9afd65ff91019c03f004a1064907e207ca089d09;
    decBuf[3477] = 256'h100aed090f099a073506aa05d4052d072b097f0a380b900a2b09d00635052a03;
    decBuf[3478] = 256'h4e019dffa4fd40fba5f99af7cef615f64df6e6f614f7eaf6ddf518f4ecf1e1ef;
    decBuf[3479] = 256'h05eed0ec98ec65ec93ecbeece4ec92ed30ee87ee6dee97ed5becdfea14e95be8;
    decBuf[3480] = 256'h43e710e7e1e6b7e644e6dbe5bfe419e390e191e006e030e0f0e0e4e1c1e251e3;
    decBuf[3481] = 256'h37e34ee339e34ce33be3a8e282e15be0b5de9cdd03dd78dcfadbedda28d9fcd6;
    decBuf[3482] = 256'h86d532d470d489d554d77fd98bdb67dd17dfa0e09fe187e205e3dfe230e211e2;
    decBuf[3483] = 256'h2de219e3b4e4ade601e836e9fde8cae83fe86de7ade644e6e5e58fe575e52ee5;
    decBuf[3484] = 256'h18e553e565e575e566e5b8e4b3e3bfe2e2e152e138e150e165e12ae166e07bdf;
    decBuf[3485] = 256'h5ede51dde9dc8adc34dcb1db4dda82d8d1d649d5e4d3fcd229d2b6d1d9d177d2;
    decBuf[3486] = 256'h7ad385d526d809dcb2e054e6a2eb36f346fadbfe5c06670bfd0f28146e167f18;
    decBuf[3487] = 256'h601af11a881de21fbb235b27a52aee2b512c422b0229f726a325f3236a22d121;
    decBuf[3488] = 256'he920132120222b24cb264529852b902d6c2f1c3186336a36e939253e4443b646;
    decBuf[3489] = 256'h184b144fb452ef56eb5a8b5ec662e667586bba6fb6734c76a6781479b078a177;
    decBuf[3490] = 256'h61752b72516ea96947654b61b45e4b5dde5c7a5c205c845a7958155631537850;
    decBuf[3491] = 256'hff4d1b4b6248e945a9439e41c23f113e383b7f3851357731e12e872c632a7228;
    decBuf[3492] = 256'h6227c725bc235821cf1d851ad0152e10e00a0d062affbff8eaf29ced2aea08e7;
    decBuf[3493] = 256'h30e499e13fdf41dcc1d877d578d287d0c2cecbcd81cdb5cc77cc5ecb5fca77c9;
    decBuf[3494] = 256'h51c8ddc775c755c7abc762c897c966cb0ece87d0c7d2d2d49ed5dcd514d6e1d5;
    decBuf[3495] = 256'h0fd68ed64ed7fcd7d9d869d9ecd992da55db40dcdbdd64df2fe1d6e39be57fe8;
    decBuf[3496] = 256'h37ebb1ed3af175f571f911fd5b003504d407100c2f11c418d31f3f26bf2dca32;
    decBuf[3497] = 256'h3539603d2a413b435d4612489f49094b074ef94f725256558156db5689561355;
    decBuf[3498] = 256'h47540a544254db541f564657a058e459635a225b005ba15a9e596458e9568455;
    decBuf[3499] = 256'hf9547a54a15409556855bf55a4559f54655396516a4ff44d184c684a50498547;
    decBuf[3500] = 256'h59454e43ea404e3fd93dfd3b5539dc36af32b22e0a2aa825ac21151fda1ade16;
    decBuf[3501] = 256'h4714fd10d90e210cf20819057000cefa80f5adf08cedd7eb52ebdaea91e967e8;
    decBuf[3502] = 256'ha2e607e591e3c5e288e2c0e259e32ae300e3f4e1ffe064dfdbdd76dc8fdb10db;
    decBuf[3503] = 256'h9dda7ada1bda8cd9d5d82ed86cd7b5d680d505d4d4d1c9cfedcdc1cbe1ca9dca;
    decBuf[3504] = 256'hdbcaf3cbf2cc37ceb2cfe3d184d4fdd63dd948db9cdc4cde65dfcae00fe2e1e2;
    decBuf[3505] = 256'h54e377e3d9e210e28de176e138e2c0e3b9e51de85dea68ecccee67f0ddf1a9f2;
    decBuf[3506] = 256'he7f2aff216f28bf10cf199f076f096f079f0c8f00ff1d1f1f1f24af48ff50af7;
    decBuf[3507] = 256'h09f8f1f8c3f983fa32fb0ffc2cfca9fbd3fa24f9f8f658f4def19eeffeec39eb;
    decBuf[3508] = 256'h9ee9bee87ae8c0e7f9e760e7d4e6aae6eae53ce51fe479e280e01cdedcdb67da;
    decBuf[3509] = 256'h23dae5d91ddab6dae4da0fdbe8da80dae1d952d9cfd8e7d87ed9a5da20dc85dd;
    decBuf[3510] = 256'h10dee6dd26dd60dbb0d927d8c2d67ed5ffd43fd491d371d3e2d2c8d280d214d2;
    decBuf[3511] = 256'h64d1bdd0a4cf98cea3cdc6ccfdcb17cc2fccc6cceccdbfcecccf7ad09ad07dd0;
    decBuf[3512] = 256'hcbd013d1d5d1f5d201d46ad4c9d439d4b6d3ced3e4d3bcd4bed5e1d5c2d5f8d4;
    decBuf[3513] = 256'ha5d3bdd293d26cd21bd3b9d30fd4f5d30dd4f7d380d469d585d6dfd780d999da;
    decBuf[3514] = 256'h32db60db36db76da82d9a5d815d82fd876d864d942da98da49da44d97fd7cfd5;
    decBuf[3515] = 256'h46d4e1d2b2d2dcd250d344d4a0d5e4d608d913db77ddb7df58e2d1e45ae8a4eb;
    decBuf[3516] = 256'h34f182f6b5fc8b025506c709e80cc10f4510ae11d213c315f218cb1c6b20a624;
    decBuf[3517] = 256'ha328392b932d002e642e092e132d072b2b290027f424a0236c22342267224e23;
    decBuf[3518] = 256'h2124c725c0279c29bf2c993038347338703c0f404b442347ba49234b6b4ccf4c;
    decBuf[3519] = 256'hde4dd54ee050cc5313580f5caf5fea639f652d67a56738670d669463af60f75d;
    decBuf[3520] = 256'h7d5b9958e155b252b44f344cea48eb45fa438041403f353d493a583893365334;
    decBuf[3521] = 256'h48325c2fdd2b9228b8241921ce1dd01a1718e914ea11320f6d0d2e0b2209be06;
    decBuf[3522] = 256'hda035b0010fd11fa92f638f43af148efcfeceae932e7b8e41de37ce003de7ada;
    decBuf[3523] = 256'h2fd756d3adce4cca73c7d3c37ac156bf65bda0bb4ebb6ebab2baefba98bb97bc;
    decBuf[3524] = 256'h38be31c00dc239c4afc57bc634c76cc79fc7cdc7f8c76bc8d3c8b1c926cb57cd;
    decBuf[3525] = 256'hf8cf27d325d6ded857dbf2dcfede52e002e28be3bce55de8d6eabaed73f0ecf2;
    decBuf[3526] = 256'h2cf537f78bf8b7fa2dfc09feb000df03b807610c03125117841daf2179254c2a;
    decBuf[3527] = 256'had2eaa325237b43bb03f50439a46be48764bf04d8b4f015145518c50034f064c;
    decBuf[3528] = 256'h2c4896454b420341d83f143e783c6d3a91386536f0342434e633ae33e1336c34;
    decBuf[3529] = 256'h96340935b73598357b35f834233420332c320f31b62f712ef62c912bf029f727;
    decBuf[3530] = 256'h0b2552226f1ecf1a7518521660149c12b70fff0cd009d2061904a001bcfe03fc;
    decBuf[3531] = 256'h20f880f445f049eca9e85ee585e1dcdc7bd87ed4d6cfb5cc23cc95ca1dca8bca;
    decBuf[3532] = 256'heeca49cb3fcc20cd74ce2dcf65cf98cfc6cff0cf17d0aecf4fcfc0ce09ce33cd;
    decBuf[3533] = 256'h6acc7fcba1cad8c955c9afc818c819c7dfc5b8c4f8c3d5c373c403c586c5fcc5;
    decBuf[3534] = 256'hbbc5a8c5ddc54fc62cc749c856c9d5caa0ccccce6dd1e6d326d6c7d840dbdcdc;
    decBuf[3535] = 256'h7cdfabe2a9e562e890ebb4ed6cf0e6f226f59bf6dff6a2f6f9f560f5d5f4fff4;
    decBuf[3536] = 256'h72f521f6fef6c7f7b2f80efab0fb39fd04ff38005101ea01180242021c02f901;
    decBuf[3537] = 256'h5b010501b600100079ffa1fed8fd55fd3dfdd5fdfbfe1f012a0306053b06e306;
    decBuf[3538] = 256'hb00625065205f903b402910085fea9fc7efa72f896f6e6f45df392f167eff1ed;
    decBuf[3539] = 256'h15ec65eabce923e998e86ee848e8dfe780e7f0e6a2e6bae67ce79ce8f5e9f3eb;
    decBuf[3540] = 256'hcfedfbef71f14df306f4aef4e1f4b3f435f4dbf23af141efededb8ec80ec19ed;
    decBuf[3541] = 256'ha4ed77ee9dee34ee57ed1beca0eaa1e95ce835e7dce597e41ce3b7e116e0fdde;
    decBuf[3542] = 256'h64de7cddfedc8bdc22dcc3db19dc9cdcd1dd4cdf17e143e3b8e494e6c9e7e2e8;
    decBuf[3543] = 256'he1e925eba0ec05ee4aef1df0ddf0fff0e0f0c3f0a9f062f0caeff2eef0edfcec;
    decBuf[3544] = 256'h5decceeb4beb46eac6e8fbe64be5a3e470e4fbe479e59fe5c2e5a3e586e5d4e5;
    decBuf[3545] = 256'h7be612e74de7d0e6dce5a2e47be3a2e321e5b8e751ecf3f141f774fdf504040c;
    decBuf[3546] = 256'h70124518931dc723f227382a492c6a2ffc2f9232ec34eb37a33a1d3d133e5e3e;
    decBuf[3547] = 256'h1a3ee53c5c3b9139e1375836593571349c34c2342b354736a137e538b53ae03c;
    decBuf[3548] = 256'hec3ec840f342ff446347a249434c724f70526254db561b59915ae55b105eb160;
    decBuf[3549] = 256'h4a65ec6a3a700c756e79477cd47d4d7edf7db57c3b7ab37668738e6fef6ba468;
    decBuf[3550] = 256'hcb643462da5fb75dfe5a3a595656d6529b4e9f4aed449f3fcc3a6b366e32cf2e;
    decBuf[3551] = 256'h842b86280625bc217320491fee1e401ff61e2a1ef51cfc1a20197916ff137610;
    decBuf[3552] = 256'h2c0d5209b30568026affeafb9ff8a1f55af182eee2ea88e88ae5d1e2a3dfc9db;
    decBuf[3553] = 256'h2ad8dfd406d16fce15ccf2c9c7c8b8c7c1c6e1c58dc4ddc254c155c06dbfeebe;
    decBuf[3554] = 256'hc8be76bf93c0ecc18ec387c5ebc774cbbece73d3d5d7d1db67dec1e00ae234e3;
    decBuf[3555] = 256'h8fe385e4d0e414e552e58ae589e62ae824ea88ec6cef5df122f362f56df749f9;
    decBuf[3556] = 256'hf0fbb5fd990051038006590a020f6413a719d21d2023f227142b102faf32fa35;
    decBuf[3557] = 256'hf838ea3a633d484000437a455e48164b904dd04f45519952ce53e7541a55eb54;
    decBuf[3558] = 256'hc1544e545a537d527a51fa4f2f4e884b0f492a467243f840b93ead3cd13a183a;
    decBuf[3559] = 256'h7039d7380539873860383d381e383b3889384238d637253720367135d3347d34;
    decBuf[3560] = 256'h2f34e733503351321731f32ee82cfc297d263223581fb01a4e165212a00cd608;
    decBuf[3561] = 256'h650503012afe94fb49f86ff4c7ef65eb8ce8ede493e295dfdcdc63da23d818d6;
    decBuf[3562] = 256'hc4d40ad442d40fd49bd4c5d438d5e6d5c4d61ad768d780d796d7a9d7dfd730d8;
    decBuf[3563] = 256'h97d8bfd8b3d83ad847d781d5d1d3d8d184d0d4cebbcd22cd97cc6dcc46ccafcc;
    decBuf[3564] = 256'h0ecd9ecd20ce67cea8ce32cf8bcf1dd0f5d0f8d132d3add412d66dd851db0ade;
    decBuf[3565] = 256'h83e00ce466e664e956ebcfed0ff01af2f6f322f62df809fab9fb42fd41feccfe;
    decBuf[3566] = 256'h4bff71ffdaff78000801f3019102ae02f701930062fec1fbfcf9bdf747f67bf5;
    decBuf[3567] = 256'hc2f419f480f398f2c6f106f112f074ef1def66ee1fee0aeef6ed2cee7deec7ee;
    decBuf[3568] = 256'hefee13ef08effeee3eef78ef9defdbefe3efebef0df020f01af001f0bbef25ef;
    decBuf[3569] = 256'he1ed29eb38e9bee623e5ade3d1e19de014dfafdd6adcefda8ad98cd738d603d5;
    decBuf[3570] = 256'head351d3c6d2f4d1cdd1f0d110d2d9d2c4d362d4f2d440d529d56ad5f3d570d6;
    decBuf[3571] = 256'h02d7b3d7cbd78ad74fd78ad66bd55ed4dfd27ad192d0bfcf99cf01d0a0d069d1;
    decBuf[3572] = 256'h20d267d27dd2b7d25ed20dd2a6d1ddd02ecff9cd00cc24caefc866c767c639c6;
    decBuf[3573] = 256'h0fc682c676c753c856c990ca63cb09cd02cfded085d34ad5e5d65bd827d964d9;
    decBuf[3574] = 256'h9cd935da64da8eda68da73d918d819d6b5d31ad20fd0bbce02ce59cdc0cc92cc;
    decBuf[3575] = 256'hbccc49cc6ccc0dccf0cb0acc52cce9cce8cd22cf49d0efd1e8d3d4d654da8fde;
    decBuf[3576] = 256'hafe3e2e90dee5bf3cdf6eef9eafd8a01d404ae084d0c891085142518601c391f;
    decBuf[3577] = 256'hcf2129244d267727d2272428d9270d27cf269726fe257325a02447230222dc20;
    decBuf[3578] = 256'hcf1f661f861fdc1f9320c82143230e253a274529a92b442d4f2f2b3157338d36;
    decBuf[3579] = 256'h8c39d23dcf417746d94ad54e7552cf54f2561d582c59da588f58c3570a57d256;
    decBuf[3580] = 256'h39565155d6533f51104e374a97466b41983c37383a349b30602c6328bb23591f;
    decBuf[3581] = 256'h5d1bb4165312330dc109a006c7033902d00088ffebffdcfe8afe3ffeebfc3bfb;
    decBuf[3582] = 256'hb2f9e7f736f61ef553f3a3f11af0e9ed73ec1feb6fe956e857e7b6e5bde3e1e1;
    decBuf[3583] = 256'hbedebfdb40d804d408d069cc2dc831c49bc150be2cbc74b9afb7b9b66eb63ab7;
    decBuf[3584] = 256'hf3b70cb90bba4fbbcbbc30be2ec092c2d1c4ddc6b9c860cbd9cd19d0e5d384d7;
    decBuf[3585] = 256'hcfda84dfe5e3e2e781ebbcef95f223f47df6c5f7b7f9c6fa06fd11ff65009a01;
    decBuf[3586] = 256'hb2024b037a03f8036b04a505c9076a0a980d721111155c18351cde203f253c29;
    decBuf[3587] = 256'hdb2c2630ff339636f038ee3b6e3fb84292462849734c4c50e3523d556057c457;
    decBuf[3588] = 256'h1e5871582658e2572957f0565756cc55a5549953d35123502a4e4e4c9e4a1549;
    decBuf[3589] = 256'hb047b2454e436a40b13d383bf8388237b636fd3574340f336e31e52f802e982d;
    decBuf[3590] = 256'hc52c522c5e2b812a7e29fe27ff26bb253f247422c420cb1e671ccc1a2b18b215;
    decBuf[3591] = 256'hcd1215109b0db70a3807ed03ee006ffd24fa4bf6abf261efacea4ae64ee2afde;
    decBuf[3592] = 256'h64db8bd7f4d4a9d1abcef2cb2eca93c8b2c7f6c7b0c858c9bdca5ecc58ce34d0;
    decBuf[3593] = 256'hdbd254d5f0d6fbd84fda08db40db73dba2db77dbebdb53dc31dd33de6ddfe8e0;
    decBuf[3594] = 256'h4de2efe307e56ce654e7d3e7ace744e766e62ae503e4aae265e1e7e00de101e2;
    decBuf[3595] = 256'h5de35be5bfe7ffe9a0ec19ef59f1faf328f727fa6dfe4601e50430082f0be70d;
    decBuf[3596] = 256'h6110a01241150617a11881194d1a8b1ac31af61a6b1a411ace191f19c0186a18;
    decBuf[3597] = 256'h7f17a2162c15c71325129d10380ff30d240c730a7a081606d60361028500d4fe;
    decBuf[3598] = 256'h4cfd4dfcc1fb97fb0afc73fc93fce9fc03fdebfc01fd3cfdddfd9ffe22ff0aff;
    decBuf[3599] = 256'h9efe78fda8fb74faebf852f880f856f87cf814f876f7acf6c1f565f421f351f1;
    decBuf[3600] = 256'h26ef85ec0beacce7c0e5e4e3b0e297e132e0edde72dd73dc8bdb0ddb9adaebd9;
    decBuf[3601] = 256'h8dd970d921d939d97ad9dcd912da43da16dab9d964d917d949d9d2d9f8da1cdd;
    decBuf[3602] = 256'h27df7be02be2b4e3b3e49be56ee6e1e604e7a5e6dbe525e54fe44ce358e2bae1;
    decBuf[3603] = 256'hf1e06ee086e09be025e1e9e138e220e2dfe156e144e1d6e1aee2eae365e5fee5;
    decBuf[3604] = 256'h2de6abe61ee7cde7e9e8f6e930eb02ec75ec24edc2ed52ee3defdbef31f017f0;
    decBuf[3605] = 256'hd0ef64efb3eeddeddbece6eb8beaa3e97ce8bce799e7f8e7c1e849eab2ec97ef;
    decBuf[3606] = 256'h16f342f815fd77019606080a6a0e6612f4133e176219531bcd1db1206a234d27;
    decBuf[3607] = 256'he4292e2d2d301e32e333da342435e03427345f342c34b7348a354a36f836d936;
    decBuf[3608] = 256'h493629351d34573223317a304730d230f9315333ae35ed376339b73a703b193c;
    decBuf[3609] = 256'hb23cf63dc63f6d425046f0493b4d3950f252b654ad55f8554c570558ad58ac59;
    decBuf[3610] = 256'h375a615aee59fa589e57fd559453af50f74d134a744629432b40e43be8374834;
    decBuf[3611] = 256'h1c2f4a2ae825c820561df518d513020fa00ac8072804ce01abffb9fdf5fb5afa;
    decBuf[3612] = 256'he4f808f7d3f52bf5f8f483f555f62ff6c6f56bf46cf208f0c9ed28ebaee86fe6;
    decBuf[3613] = 256'h63e4ffe1c0dfb4ddd8db28da2fd853d6a3d439d255cf9dcc23cae3c743c57ec3;
    decBuf[3614] = 256'h3ec133bfdfbd26bd7ebcb1bcdfbc09bd2fbd52bdf0bd2dbffcc0a3c31dc601c9;
    decBuf[3615] = 256'hbacb33ce17d197d4d2d8cedc77e119e7e3eab6efd7f2d3f673faaefe6300fa02;
    decBuf[3616] = 256'h6304d10434058f05e105c1061508c5092f0c6e0ea511a3145c178a1a891d7a1f;
    decBuf[3617] = 256'hf4213324d426032a012d48312034c0371a3a3d3c2f3ef33f33423e441a46cb47;
    decBuf[3618] = 256'hc449a04b504dd94e3e502651f8516b524952aa51a850284fc34dc54b61492147;
    decBuf[3619] = 256'heb43ec40343e053b07384e35d5329530f42d302c952a1f2953281e2795256423;
    decBuf[3620] = 256'hc420951d971a1717bd14bf11cd0f540db80bad09d107a5059a03be0117ff9dfc;
    decBuf[3621] = 256'h02fb8cf938f888f6fff434f309f1fdee21ed71eb78e924e8f8e5ede301e148de;
    decBuf[3622] = 256'h1adb1bd863d534d236cf7dcc4fc92bc773c4f9c1babfaebdd2bb22ba7ab9e1b8;
    decBuf[3623] = 256'h6cb93fba98bb39bdc2be8dc0c2c14bc34ac48ec50dc6cdc67bc758c8cec999cb;
    decBuf[3624] = 256'hc5cd66d0dfd21fd52ad706d93bdac4dbc3dc07de2edf88e070e1eee161e23ee2;
    decBuf[3625] = 256'h5ee241e25be2d2e2c0e35ee49ae56de679e76ee8c9e9b1ea2cec2bed70ee97ef;
    decBuf[3626] = 256'hf0f035f204f430f63bf817fa43fc4efeb200f202fd046107fd08720a3e0bf80b;
    decBuf[3627] = 256'hbf0b8c0b5e0b340bc10acd09b0080a078105b6030602ed0088ffa0fe79fd20fc;
    decBuf[3628] = 256'hdbfab5f90ef886f621f5dcf3b5f2a8f16ff048ef3bee8ded2eed4bedcded73ee;
    decBuf[3629] = 256'hb8efa0f072f1e5f108f2a9f153f19cf026f0e5efaaef2defbbeedeed82ec3deb;
    decBuf[3630] = 256'h6ee9bee735e6d0e4e8e315e309e2cfe0a8df02de79dc14dbcfd9a8d89cd762d6;
    decBuf[3631] = 256'h3bd52ed4f4d222d2afd146d126d143d15dd1a5d13cd2edd2c2d3ffd4d1d5ded6;
    decBuf[3632] = 256'hd2d7afd83fd9f6d96ddaaedae8dafadaeada16db09db46dbbfdb30dc0edd2ade;
    decBuf[3633] = 256'h37df71e098e1a4e298e376e492e4e1e4f9e4b8e456e4fce349e3a3e2e1e1c1e0;
    decBuf[3634] = 256'hb5dfc0dee3dd53dd39dd80dd43de2edf4be057e14ce229e3b9e33be4b2e4f3e4;
    decBuf[3635] = 256'hdfe4aae438e4b3e336e305e332e3c5e3ebe412e61fe713e8f0e880e9d3ea18ec;
    decBuf[3636] = 256'h3ceedcf00bf409f789fad4fdd2001905f107910beb0d330f5e102212bd13c915;
    decBuf[3637] = 256'hb5186d1b511ff0224a254928012bc62c612ed72fa3305c31043237321f334634;
    decBuf[3638] = 256'h53358c365f37d237af3750378736d0355a35c234fd34333563359035d335ae35;
    decBuf[3639] = 256'hfb3591367f371a39133b773d5c40db432647ff4a9f4ee9510d54fe550e570558;
    decBuf[3640] = 256'h4f580b58ce5725578c56a455d25412541e53c2512050b74d774b414843458a42;
    decBuf[3641] = 256'h5c3f5d3ca53976369d32fd2ec22ac5261d22bb1dbf191f16d512d60f570cfd09;
    decBuf[3642] = 256'hfe064604cc01e8fe30fcb6f976f76bf59ff46af3c2f2c3f1dbf060ef61eec0ec;
    decBuf[3643] = 256'h37eb6ce9bce752e512e372e0f8dd5ddce7da0bd9d6d7ddd501d4d6d135cfbbcc;
    decBuf[3644] = 256'h7cca70c80cc671c491c3c5c20cc2d3c1a0c172c19cc1c3c1e5c184c24dc338c4;
    decBuf[3645] = 256'h55c5aec64fc8d8c909cc14ce78d05dd315d644d942dcfbde29e203e6a2e9deed;
    decBuf[3646] = 256'hdaf179f5b5f9b1fd5001aa03a9066109db0b760dec0ec81078127114d516b919;
    decBuf[3647] = 256'h721ca01f9f221e267828772b682d2d2f6d317833dc351c3891396d3b993d0f3f;
    decBuf[3648] = 256'h6340984140423f438444aa4551474a499e4ad24beb4c1e4df04c714cfe4b504b;
    decBuf[3649] = 256'hb24aaf497548fa462f457f438641223fe23cd73a7338d736373472323230272e;
    decBuf[3650] = 256'hd32c232b9a293528f026752510246f227620121ed21b3119b8167814d7115e0f;
    decBuf[3651] = 256'hc20db70bdb09af070f054a03af01a4ff50fe1bfd92fb2dfa2ff853f627f4b1f2;
    decBuf[3652] = 256'h4df0b2eea7ec43ea03e8f8e594e354e1dedf02decedc45db46da5ed937d82ad7;
    decBuf[3653] = 256'hf1d5cad4bdd3c9d2ecd1cfd1e9d18fd27dd39ad45ad508d667d6f7d6add7b3d8;
    decBuf[3654] = 256'h78daa4dc45df73e272e52ae859eb7ced35f044f1dff22af36ef327f45ff45ef5;
    decBuf[3655] = 256'h46f66df77af86ef98bfa97fbd1fc4cfeb1fff6007102d603770590068f077708;
    decBuf[3656] = 256'hf508b509630a020b910b140c8b0ccc0c7c0d520e8e0fb5100e12f6121d14dd14;
    decBuf[3657] = 256'hd115af16b1176018fe181b190019181903193d19731983191c195318de161315;
    decBuf[3658] = 256'h621369118d0f590ed00c6b0b260aff08f307730674058c046503590264010900;
    decBuf[3659] = 256'hc4fe49fde4fb42fabaf8eff63ef545f3f1f1bcf0a4efa5ee1aee9bed75ed52ed;
    decBuf[3660] = 256'hf3ecd6ec88ece2eb1feb68eac2e9ffe87de8d7e714e75de628e5ade348e24ae0;
    decBuf[3661] = 256'h6ede39ddb0db4bda64d9e5d8bfd8e2d801d9e5d8cad824d862d7abd6a5d56cd4;
    decBuf[3662] = 256'h99d3d9d22bd20bd228d276d21cd389d339d4dfd477d5d9d59ed620d7f6d7bfd8;
    decBuf[3663] = 256'h42d9e8d9d6da74dbb0dcd7dde4ded8dfb5e045e1fce1a2e23ae311e4a1e4f0e4;
    decBuf[3664] = 256'h37e521e5e6e4b1e480e454e47ce4e9e46ee50fe6d1e654e7cbe70be846e858e8;
    decBuf[3665] = 256'h68e85ae832e8f5e7d4e7dee7f9e723e839e817e8dee79be749e728e75ae787e7;
    decBuf[3666] = 256'h03e8ece8c9e93feb0aedbaee43f074f27ff4e3f6c7f947fd82017e051e09590d;
    decBuf[3667] = 256'h5611f5144f174d1a3f1c6d1f912110256a27692a5a2cd42e6f304f311b32d532;
    decBuf[3668] = 256'h0d33da32ab328132a8321033f132d43251324c3158307a2fb12efa2d542d912c;
    decBuf[3669] = 256'h432c2b2c6c2c6b2da52e782fd1305c312f32ef32e3330035a6362f38603a003d;
    decBuf[3670] = 256'h7a3fba415a441f46ba473049844ab94b414da64e8e4fb84f454f0b4ee54cf24a;
    decBuf[3671] = 256'h8e484e46ad437f40803d013ab636dd32342e132bf3252021bf1c9f17cc126b0e;
    decBuf[3672] = 256'h6e0ac605a502ccff2cfcd2f9d4f61bf457f217f076edfdeabde8b2e65ee529e4;
    decBuf[3673] = 256'h81e34ee31fe3a1e2e1e133e116e00adf15de38dda8dcf1db4bdb5dda80d97dd8;
    decBuf[3674] = 256'h43d71cd676d47dd2a1d0facd35cc9acabac9eec8b0c808c809c721c6fac487c4;
    decBuf[3675] = 256'h64c484c4a0c4bbc402c599c598c65ec80eca07cce3cd0fd0b0d229d50dd88ddb;
    decBuf[3676] = 256'hc8dfa1e240e67cea55edf4f03ff418f8affaeafec3016b068d09890d1f106a13;
    decBuf[3677] = 256'h681621199a1bda1de51f4922e523f025cc277c29052b9e2bcc2ba22bc92bec2b;
    decBuf[3678] = 256'h4a2cda2cf42c3c2d512db32d542e422f1f305c312e323b33e933c7345635a535;
    decBuf[3679] = 256'hec35023664369936eb36dc369936fb356435b3349c3486349a3488345734d233;
    decBuf[3680] = 256'h0e332332c730252fbc2cd8295826fe232520851c2b1a5216b212680f690cea08;
    decBuf[3681] = 256'h9f05c60126feebf9eff558f30df0eaedbfecfbea60e9eae71ee76ee5e5e31ae2;
    decBuf[3682] = 256'heedf78de9cdc68db4fdaead8a5d77ed625d53dd46bd3abd242d222d2ccd1b2d1;
    decBuf[3683] = 256'hcad189d175d140d10fd100d1d8d0b4d07dd04bd0f9cfaccf7acf27cf06cffcce;
    decBuf[3684] = 256'he1ce0acf7bcf0dd0e5d0e8d1dcd2f8d305d53fd6bad71fd9c0da49dcaedd96de;
    decBuf[3685] = 256'hbddfcae08fe2bbe4c6e62ae96aeb75edd9ef19f224f488f623f82ffa0bfc3ffd;
    decBuf[3686] = 256'hc8fe2d007201990259034d04eb047b059505ac056c050905b0041e04bc038603;
    decBuf[3687] = 256'h55038203df03040425044304de036603b302ae01ba00dcff13ff28fec9fd39fd;
    decBuf[3688] = 256'hb7fc9ffc33fca9fb2cfb9afa11fa94f9c0f8f7f70cf7b0f56bf4f0f2f1f1adf0;
    decBuf[3689] = 256'h86efe0ed57ec8ceadce8e2e68ee5dee355e256e112e03fdfccde63de04dee8dd;
    decBuf[3690] = 256'h65ddbfdc53dc7bdb78dacad9add854d70fd694d42fd3ead1c3d0b7cfc3cee5cd;
    decBuf[3691] = 256'h56cd07cdc0ccd6cc38cdb5cd47ce1fcfafcf9ad077d140d2c3d269d3aad30cd4;
    decBuf[3692] = 256'h89d4fbd49dd560d617d7edd7efd89ed9bada7adb29dcc7dc1ddd37dd7eddbfdd;
    decBuf[3693] = 256'hfadd54dee6de6fdf10e0d3e021e198e1d9e13be223e37fe420e61ae8f6e92aeb;
    decBuf[3694] = 256'h43ec42edcdeda0eeacef2cf191f232f4bbf520f765f837f9f7f91afa3afa1dfa;
    decBuf[3695] = 256'h37fa4ffa90faa3fab5faa5fa96fa6efa4afae7f96ef9bcf8e6f7e3f6a9f5d7f4;
    decBuf[3696] = 256'h17f4aef38ff3abf3faf341f4adf436f590f522f621f75bf8d6f93bfb39fd15ff;
    decBuf[3697] = 256'h4101e20310070f0ac70cf60ff412e6145f179f19401cb91e9e218f23be26bc29;
    decBuf[3698] = 256'h752cee2e2e3139338d3446357e35b135e035b6358f356c350e35f1343a343533;
    decBuf[3699] = 256'hfb312b307b2ef22cf32b0b2b362ba92bcc2b6a2cc02c0e2db52da22e412f7d30;
    decBuf[3700] = 256'ha431b0323034fb35ab37a439803b313d2a3f0641b6421f455f47004a794c154e;
    decBuf[3701] = 256'h8a4fde5013524b5218528d516650c04e574c7249ba46d642373fec3b3837d632;
    decBuf[3702] = 256'hda2e312ad025b0203e1ddc18e0144011f60d1c0a7d0632033400b4fc5afa5cf7;
    decBuf[3703] = 256'ha3f42af28ff083ee2fed76ecceeb9bebc9ebf3eb1aecc8ece8eccbece5eccdec;
    decBuf[3704] = 256'h0eed70edededc1ee8aef0cf024f0e3ef33efceed69ec6bea07e8c8e5bce3e0e1;
    decBuf[3705] = 256'hace093dffadeccde4ddedadd71dd94dccbdb14db9dda5cda97da14dbe8db24dd;
    decBuf[3706] = 256'hf3de1fe1c0e3eee6ede9a5ecd4efadf34df797fa4cffae03aa07520cb410b014;
    decBuf[3707] = 256'h50188b1c8720302551284d2ced2f38333636b6390f3ce93f7641d043f4455746;
    decBuf[3708] = 256'h6747b9470448484886484d48b4472947ab463846cf4570451a4597442144e043;
    decBuf[3709] = 256'hf3432944dc4453459345f6450746f74506461346074628460a4601460946e445;
    decBuf[3710] = 256'h8a4536459144bb43f2429e415940323f8c3d033c383a0d3801369d335e31272e;
    decBuf[3711] = 256'h042c84283a256021b81c56185a14b10f500b30065d01fbfcfff857f435f15dee;
    decBuf[3712] = 256'hbdea63e840e64ee48ae2efe00ee0bade01dee8dc83db9cdac9d909d9a0d842d8;
    decBuf[3713] = 256'hebd79dd756d740d77bd7f8d7cbd895d94bdaf2da5edb71db60db2fdbc8da4fda;
    decBuf[3714] = 256'hbdd934d9b6d824d8c2d745d7f4d6aad69dd690d6ddd65fd7ddd78fd836d9cdd9;
    decBuf[3715] = 256'ha5daa8db9cdc76de52e07ee21fe598e7d8e9e3ebbfed6fefd9f118f424f610f9;
    decBuf[3716] = 256'hc8fb42fe2601de0358069808380bb20d4d0f5811ac12e1138a14231551157b15;
    decBuf[3717] = 256'h55153215d314b614681450140f14d4139f132d13e312a0121b129e11cb108e0f;
    decBuf[3718] = 256'h130eae0c0d0b84091f08da065f05fa03b6028f01cf00dbff3dff3afe46fd29fc;
    decBuf[3719] = 256'h1cfb6efa51f992f858f7ddf578f433f3b8f1b9f074ef4deef4ec53ebcae965e8;
    decBuf[3720] = 256'h20e7f9e5a0e45be3e0e115e065de6cdc90da64d8c3d5ffd363d2eed022d0edce;
    decBuf[3721] = 256'h45ce46cd5ecc8bcb65cbb6ca57ca01cab3c9cbc90bca95ca36cbcdcb08cc3ecc;
    decBuf[3722] = 256'hafccf9cca7cd7dce0ccfc3cf99d0efd0a6d11dd25ed223d2edd13bd1c4d0d9d0;
    decBuf[3723] = 256'hedd08ed17cd259d35cd496d511d776d817da30db2fdc74ddf2ddb2de60df41df;
    decBuf[3724] = 256'h5ddf77df01df16df51df63dfd5df95e017e1bde180e2cee275e30ce447e4e8e4;
    decBuf[3725] = 256'haae52de603e7cce74fe8f5e88ce916ea93ea05eb13eb21ebfceaafea7dea50ea;
    decBuf[3726] = 256'hf5e9a0e927e9d6e8aae8d2e83fe9c4e941ea92eadcea04eb59ebfeeba4ec92ed;
    decBuf[3727] = 256'heeee32f002f22df4cef648f92cfcabff05020405bc078109c10bcc0d30101413;
    decBuf[3728] = 256'hcd154618cf1b291e2721e023a4253f27b528f928b2295b2af42a7f2bfd2b242c;
    decBuf[3729] = 256'h012ca22bd92a222a4c298328cc2726276326ac253525c924b624eb241c25be25;
    decBuf[3730] = 256'h5626df26a4278f282d29a32a082c062ee22f0e321934f535a5372e39933a343c;
    decBuf[3731] = 256'hbd3dbc3ea43f774083413242d0422643a342fd41b940173f8f3d5e3b52396636;
    decBuf[3732] = 256'hae33ca2f2b2cef27f3234b1fe91aed164412e20dc308f003cf00d3fc33f9e8f5;
    decBuf[3733] = 256'h0ff278ef1fed20ea68e7eee4aee2a3e0c7de9bdc26db4ad990d8e8d7b5d787d7;
    decBuf[3734] = 256'hb1d7d7d7fad759d822d9a5d91bda5cda49da13dac2d95bd9e2d82fd82ad7f0d5;
    decBuf[3735] = 256'hc9d470d388d261d108d0c3ce48cde3cbfbcad4c915c966c8c8c738c71ec765c7;
    decBuf[3736] = 256'hd2c75bc820c93fca4ccb11cd3dcfddd157d43bd7bbda05dedfe17ee5c9e8a2ec;
    decBuf[3737] = 256'h42f07df47af819fc54005104f0073b0b140fb412ef16eb1a821dbd21ba255028;
    decBuf[3738] = 256'h9b2b742f0b3274339735c236d1376d394d3a193bd23b9a3b013bd33aa83a353a;
    decBuf[3739] = 256'hcd392f396538ae3708379c363a367535be34b9330b336d321632c83181311531;
    decBuf[3740] = 256'h6430ed2f2b2fa82ed22dd02cdb2b802a3b29c0275b26b924312366213a1fc41d;
    decBuf[3741] = 256'he81b381aaf184a174c157013c011560f160d0b0b1f086705ed0264ff0bfd0cfa;
    decBuf[3742] = 256'h54f725f402f249efd0ecebe9fae780e5e5e3dae186e051dfc8dd63dc7bdb00da;
    decBuf[3743] = 256'h01d919d8f2d6e6d566d467d37fd2add186d163d144d161d146d15ed1cad154d2;
    decBuf[3744] = 256'hf5d2b7d33ad4e0d4a3d58ed66bd76ed862d900dac9da80db56dc59dd4dde2adf;
    decBuf[3745] = 256'hf4dfdfe0bce1f8e21fe479e5bde690e750e88ae905eb6aec0bee04f0e0f190f3;
    decBuf[3746] = 256'hfaf53af845faa9fc44fee500a902e904f4065809f40aff0ccb0d000fa80fa710;
    decBuf[3747] = 256'h3211b01124124612a512c212dc12f412de12cb12b912c912d812e512d9128c12;
    decBuf[3748] = 256'h46122b12f111ad115b11b610820f5b0eb50c2c0bc70925089c063705f3037802;
    decBuf[3749] = 256'h1301ceff53feeefc4dfbc4f9f9f7c4f63bf5d6f391f2c2f08def04ee9fecfeea;
    decBuf[3750] = 256'he5e980e899e772e618e530e40ae3fde109e12be029df7adedcdd4cddfedcb7dc;
    decBuf[3751] = 256'h76dcb1dcc3dcf3dc3ddd30dd24ddeddca7dc42dce5db5fdbbeda27da76d9d0d8;
    decBuf[3752] = 256'h64d802d8a9d7b9d7aad708d88dd82ed9f1d9a7da1edb8adbc5dbb3dbc4dbd2db;
    decBuf[3753] = 256'haadb9edba9dbc7db3edcf0dcc6ddc9de03e07ee1e3e284e40de672e714e92cea;
    decBuf[3754] = 256'h2beb70ec42ed02eeb1ee10ef66efe8ef00f041f0a3f0fdf06ef1f3f170f243f3;
    decBuf[3755] = 256'h0df4c4f46af501f615f6dff5aef565f522f5e5f4daf4f8f426f560f576f538f5;
    decBuf[3756] = 256'hbcf4d4f3f7f2f4f146f1e7f057f03df0f6efb5efc8efb6ef28f0caf08df1e1f2;
    decBuf[3757] = 256'hdff443f783f9b9fcb7ff370391058f08480bc10d01100c12e81314161f18831a;
    decBuf[3758] = 256'hc31cf91f1d22d5249a263528ab29772aab2bc42cc32dab2ed22fde305e325d33;
    decBuf[3759] = 256'ha23474359b357835da349d3377326a3130305d2fea2e822e622e452ec32dab2d;
    decBuf[3760] = 256'hc12dfb2d9c2e8a2fa7309a32fe343d37743a723df2403c4460465148cb4a0b4d;
    decBuf[3761] = 256'h164f6a501a52335398548055a6561a57f7561956dd540e53e250d74e734c334a;
    decBuf[3762] = 256'h9247194534427c3f983bf937cd32fa2d98299c25fd21c11dc5192616ea11ee0d;
    decBuf[3763] = 256'h4e0a130617026efd4dfa51f6b1f257f00fefe4edd5ecdeeb93ebd7eb15ec4dec;
    decBuf[3764] = 256'he6ec15ed3fed18edf6ec15ed32edb5edccede2eda7ed06ed44ec58eb3ceae2e8;
    decBuf[3765] = 256'h9ee777e66ae576e499e396e2a2e1c5e0c2df88de61dd08dc66da6dd819d7e4d5;
    decBuf[3766] = 256'hccd433d404d42fd408d4b7d4d3d579d702d999db13de52e01ee4bee7f9eb19f1;
    decBuf[3767] = 256'hebf54dfa6dff40046107810cf20f54145018f01b2b202824d028f12bee2f8432;
    decBuf[3768] = 256'hde340137ba397e3bbe3dc93f1d4152426b430444324408449543e7424842f241;
    decBuf[3769] = 256'ha4412d419640e53fe03eec3d0e3d0c3c5d3b803a7d39cf383138a13752370b37;
    decBuf[3770] = 256'h9f3664362f36fe35ef35c7355a35f3342a346133de3208323f31bc30882f612e;
    decBuf[3771] = 256'h072d662bdd291228622669248d226120c01dfc1b18195f1631133210b30c6809;
    decBuf[3772] = 256'h8e05ef01b4fdb7f918f6cdf2cfef16ed9deab8e7c7e5b7e41ce3a6e152e01edf;
    decBuf[3773] = 256'h75dedcddaedd84ddf7dd1ade79de42dff9dfcfe098e14fe2f5e261e3eae38be4;
    decBuf[3774] = 256'h23e5d3e51be630e6f5e578e5e6e484e42ae41ae40be434e470e4e9e47be52ce6;
    decBuf[3775] = 256'h02e792e7e0e727e83de878e8d1e843e98de9eae957eabfea6ceb42ec45ed7fee;
    decBuf[3776] = 256'hfaef5ff1a4f273f423f6acf7ddf9e8fb4cfe8c00970273042406ac071109560a;
    decBuf[3777] = 256'h7d0b8a0c7e0d5b0eeb0ea20f18102e101a10320fd60d350c3c0a6008af06b604;
    decBuf[3778] = 256'hda022a0131ff55fd20fc27fa4bf816f71df541f391f108f03dee08edf0eb8bea;
    decBuf[3779] = 256'ha3e9d3e723e69ae4cfe21fe196dffdde15deebdd12deefdd4edea4def2de39df;
    decBuf[3780] = 256'h4fdfedde94dee1dd0bdd7bdcc4db1edb87da88d94ed8d3d608d557d3cfd104d0;
    decBuf[3781] = 256'hcfce46cde1cb9cca75c969c875c797c6cec517c5a0c409c4f5c34fc480c4acc4;
    decBuf[3782] = 256'h09c546c593c515c692c624c7d5c74cc88dc816c993c966caa3cbcacc23cec4cf;
    decBuf[3783] = 256'hddd0dcd121d39fd35fd499d56bd6c5d709d930dad6db5fddc4de09e030e1f0e1;
    decBuf[3784] = 256'h58e278e222e207e24fe239e274e286e255e20be219e2f4e12be299e2c6e2eee2;
    decBuf[3785] = 256'h5be3a5e338e410e5d9e5c4e6e1e7a0e84fe92ceaf5eae1eb7fec0eed91ed08ee;
    decBuf[3786] = 256'h49ee84eeb9eea9ee9aee72ee1deebaed5dedefeca6ec63ec3eec07ecadeb10eb;
    decBuf[3787] = 256'h78eaa1e911e9c2e80ae923eac9ebc2ed26f00af3c3f53cf821fbd9fd9eff8202;
    decBuf[3788] = 256'h730438061c09d50b030fdd127c16c719c51c7e1f422182236224b62566277f28;
    decBuf[3789] = 256'h4a2afa2bf32dcf2ffb31db322f346d34353402347733f93285321d327f31ef30;
    decBuf[3790] = 256'h6c30382f112e042d842b852a9e291f299229cc2a472c782e19319333d2357338;
    decBuf[3791] = 256'hed3a883c933ee73f134289436545904706495a4a8f4ba74cda4c094d8a4ccb4b;
    decBuf[3792] = 256'hd64a7b49d94750461f441442b03f273cdd3803355b30f92bd9260722a51d8518;
    decBuf[3793] = 256'hb213100e460a7405520233fdc1f95ff563f1c3ed79ea7ae789e5c4e329e2b3e0;
    decBuf[3794] = 256'h5fdf2ade12dd13dc88db09dbe3da06db25dbb5db6cdc12ddaadd0cde1ede0dde;
    decBuf[3795] = 256'hc4dd81dd2cdddfdc5ddce0db4ddb9ddaf7d95fd9d6d835d872d787d66bd55ed4;
    decBuf[3796] = 256'h24d3fdd1f1d042d0e3cf8dcfdbcf52d015d100d21dd3c3d44cd67dd888da74dd;
    decBuf[3797] = 256'h2ce0a6e22fe679e978ecbef097f336f772fb6eff0e034907450bee0f4f144c18;
    decBuf[3798] = 256'heb1b27202324c227fe2bd62e7632d034f336e538a93aa03b803c4c3d063eae3e;
    decBuf[3799] = 256'he13e0f3f393f133f363f563f723f8c3f753f5f3f243fef3e7d3ebd3dd23cb53b;
    decBuf[3800] = 256'h5c3a7439a1382e38c63728375e36a735d23408345233db32183261312d30b12e;
    decBuf[3801] = 256'hb22d112c882abd280d278425b9238d21821f2e1e021c62199d175d15bd124310;
    decBuf[3802] = 256'h5f0da60a2d0849055703de009efefdfb84f9e8f7ddf589f4d9f2e0f07cee3cec;
    decBuf[3803] = 256'h31ea55e8a4e68ce527e485e2fde098df53de80dd74dc0bdcacdb56db3cdb54db;
    decBuf[3804] = 256'h94dba8dbdedbeedbfddb25dc49dc6adcb0dcf0dc4bdda0dd03de7bdeccde34df;
    decBuf[3805] = 256'hacdf3ee0efe095e183e260e32ae4e0e487e549e600e7d6e79fe856e92ceaf5ea;
    decBuf[3806] = 256'h49eceaede3efbff1ebf3f6f55af8f5f996fc5bfe9a00a6028204b6053f073e08;
    decBuf[3807] = 256'h8309aa0a6a0b180cb60c460d940d0b0e770eb20e0b0f3c0f2d0feb0e960ef10d;
    decBuf[3808] = 256'h1b0d180c240b470a7d09920876076906750558049803a40288017b0087ff6afe;
    decBuf[3809] = 256'haafdb6fc9afb8dfa0df9a8f707f67ef419f3d5f159f0f4ee0deee6ecd9eb2beb;
    decBuf[3810] = 256'h4deabee96fe9f8e88ce851e8b1e719e769e693e590e49ce3bfe2bce1c8e06cdf;
    decBuf[3811] = 256'h27de00dda7db62da90d983d8d5d776d720d73ad781d7c2d7d5d7c4d752d708d7;
    decBuf[3812] = 256'hc5d689d668d672d644d61bd604d6d4d5c1d5c7d5a3d567d52dd5ead4ced4e7d4;
    decBuf[3813] = 256'h1cd583d507d661d6f3d6a4d779d843d996da7edba5dcfedd43dfbee023e268e3;
    decBuf[3814] = 256'h3ae447e5f5e594e696e745e861e96eea62ebbeec03eed5ee95ef43f0a2f0f9f0;
    decBuf[3815] = 256'haff156f244f360f46df51bf6f9f688f7a2f7baf779f717f79af608f6a6f570f5;
    decBuf[3816] = 256'h3ff513f5d0f47bf402f450f37af2b1f1faf024f094ef12efcaeeb5ee7aeeafee;
    decBuf[3817] = 256'h01ef68ef16f0ecf0eef128f3f8f423f75afa58fd9f019b053a09850c830f3c12;
    decBuf[3818] = 256'h6a156918211b9b1d7f203823662665291d2c4c2f6f31283437352e360e37da37;
    decBuf[3819] = 256'h9338ac39453a2d3b003c263c493cea3b213b013a5b3862368634d632bd318a31;
    decBuf[3820] = 256'h5c318631f9311c32fc31e031c531dd31a0328b33e734e536c138ed3a8d3d0740;
    decBuf[3821] = 256'h4742e744ac464748bd49114bc14c4a4e15504a516252fb52cd524f5242517d4f;
    decBuf[3822] = 256'hcc4d634b23498346094425416c3e3e3b3f38f933fd2f542bf226af20841c3617;
    decBuf[3823] = 256'h6412c10cf7082504030107fd68f91df644f2a4ee4aec4ce993e61ae47ee273e0;
    decBuf[3824] = 256'ha7dfeedeb6de83deb1dedbde4edffddfdae06ae121e2c7e233e3bde316e467e4;
    decBuf[3825] = 256'h58e4e0e32de328e2eee0c7df6edecddcb4dbe9d9b4d82bd7c6d525d49cd237d1;
    decBuf[3826] = 256'hf2cf77ce78cd90cc6acbaacafbc9dcc932cab5cabacbaecc49ce42d0a6d28ad5;
    decBuf[3827] = 256'h0ad955dc09e12ae44ae9bcec1ef13df6aff911fe31030308650c61100a156c19;
    decBuf[3828] = 256'h8b1efd215f265b2afb2d45314434fc36c1385c3a3c3b083c463c7e3c4b3cc03b;
    decBuf[3829] = 256'h963b893adb39be38b237be36a135e134ed334f33863203325d31f1308f303530;
    decBuf[3830] = 256'hc32f5c2f192ff52e162f702fdd2f7f30173179311a325b32bd3216330633f732;
    decBuf[3831] = 256'hcf324a32cc313a316230602f262eab2ce02a2f29c6268624e521b71eb81b3918;
    decBuf[3832] = 256'hee141511750d3a091a0448ffe6faeaf64af30fef12eb73e738e35fe0c8dd7eda;
    decBuf[3833] = 256'h5ad869d6a4d409d329d25dd11fd1e7d01ad1a5d123d2e3d292d3aed4bbd5f5d6;
    decBuf[3834] = 256'h70d8d5d919db40dc4ddd87deaedfbae0aee18ce2e2e2fce2b5e249e2e7e16ae1;
    decBuf[3835] = 256'hd7e027e051df88de9ddd80dcc0dbccdaafd956d811d7ead52bd57cd45dd4b3d4;
    decBuf[3836] = 256'h35d53bd675d744d9f4daeddc51dfede08de352e592e79de901ece5ee9ef1ccf4;
    decBuf[3837] = 256'hcbf783fafdfce1ff990213055307f3096d0c080e1310ef11a912511384135613;
    decBuf[3838] = 256'h2f12d510340f3b0d5f0b330928074c059c03a2014e009efe15fdb0fb0ffa16f8;
    decBuf[3839] = 256'h3af68af490f23cf18cef03ee04edc0eb99ea8ce998e8bbe72be7a8e691e6fde6;
    decBuf[3840] = 256'h86e74be836e913eaa3ea26eb6deb82eb6feb39eb08ebbfea61eaf4e9c8e94fe9;
    decBuf[3841] = 256'hbde80ce807e7cde5a6e44de308e28de08edf4ade23ddc9db85dab2d959d814d7;
    decBuf[3842] = 256'h42d6e8d400d4d9d21ad26bd1cdd03dd0bbcfa3cf62cf4ecf60cf91cfdbcf89d0;
    decBuf[3843] = 256'h2fd1f2d111d31ed412d56ed655d77cd83cd930da0edbd7dbc2dc9fdda2de96df;
    decBuf[3844] = 256'h74e003e152e16ae17fe16ce17de18ee17fe18ce198e177e181e1afe1b7e1ece1;
    decBuf[3845] = 256'h37e27de2e2e275e3fee39fe462e5e4e58be64de7d0e717e858e86ce87ee86de8;
    decBuf[3846] = 256'h41e834e840e835e867e870e878e89ee897e884e8a0e8bae8ffe881e922eab9ea;
    decBuf[3847] = 256'h6aeb10eca8eca7ed9beeb8ef5ef157f3bbf5fbf731fb2ffeaf01f904d308690b;
    decBuf[3848] = 256'hc30dc2107a13f415d818911b0a1eee206e24c826eb28a42b682d5f2e3f2f0b30;
    decBuf[3849] = 256'hc4306d310632ee32153488343635953578355e3588344c33253219312430862f;
    decBuf[3850] = 256'h302fad2e662e252ec32d8e2d5d2d312d732df92dbd2e1130b231ac338835b337;
    decBuf[3851] = 256'hbf399b3b4b3dd43e9f404f42d843a345d846f047ef48d749aa4a1d4bb44a164a;
    decBuf[3852] = 256'h4d49c5473c460b446a41f13e0d3c8d3842354432fd2d012a62263621631c0118;
    decBuf[3853] = 256'h05145c0ffb0afe06560235ff38fb99f74ef475f0d5ec7bea7de7c4e400e365e1;
    decBuf[3854] = 256'hefdf23dfe5deaddee0deb2dedcde02dfdfdec0dedcdef7de3edfaadf0ce089e0;
    decBuf[3855] = 256'hdae024e14ce140e109e19be016e076dfb3de30de8addc7dc11dc3bdb72da86d9;
    decBuf[3856] = 256'ha9d8e0d729d7b2d646d632d68cd6fed6a0d7b9d812da57db7bdd86dfeae12ae4;
    decBuf[3857] = 256'h60e75eea17edfaf09af4e4f7befb5dffa8028206210a5c0e3511d5141019e91b;
    decBuf[3858] = 256'h881fd322ac264c2a972d953015346e3692384a3b5a3c513d313efd3eb63fee3f;
    decBuf[3859] = 256'h2140f33f1d40aa3f413fe23e8c3e0a3e933dfb3c723cf53b633b013ba73a353a;
    decBuf[3860] = 256'hb139343960389737ac368f3536344e3327326731b9301b308b2f082f922ecf2d;
    decBuf[3861] = 256'h4c2da62ce42b2d2b272a3329562853275f264225e9234822bf208e1e831c1f1a;
    decBuf[3862] = 256'h3a1782140812240f6c0c3d093f0686030d0184fd39fa3bf782f409f224ef6cec;
    decBuf[3863] = 256'ha7ea68e85ce680e4d0e2d7e083dfd3dd4adc4bdb63dae5d972d994d9b4d90ada;
    decBuf[3864] = 256'h24da3cda27daecd992d962d918d925d94ad9add925dad8da7edb41dcf7dc6edd;
    decBuf[3865] = 256'h31deb3de5adf1ce007e1e5e1e8e2dce3b9e449e5cbe542e683e6e5e61be7ade7;
    decBuf[3866] = 256'h5ee833e936ea70eb97ecf0ed35ef5cf0b5f1faf221f47af5bff6e6f78cf915fb;
    decBuf[3867] = 256'he0fc90fe19007e01c202e90343052a06510711080509e309720af50a9b0bdc0b;
    decBuf[3868] = 256'hf00bba0b280b770aa20965083e0732063e05e203fa02d30113011f00c3fe7ffd;
    decBuf[3869] = 256'h58fcfefa5df944f8dff69bf5c8f4bbf3c7f2abf19ef064ef3dee31ed3dec5feb;
    decBuf[3870] = 256'h96ea13eacce9b6e9a3e9d8e9c8e9b9e9ace957e9dee86ce8e8e747e706e7a4e6;
    decBuf[3871] = 256'h27e6b5e530e58fe4f8e3f9e205e227e125e030df53de50dd5cdcbedbf5da0ada;
    decBuf[3872] = 256'h6cd969d8bad71cd753d69cd525d5b9d47ed490d4a1d4ead463d5b4d5fed55bd6;
    decBuf[3873] = 256'h4fd644d64ed621d608d62dd650d6add65bd702d8c4d8afd98dda56db41dca0dc;
    decBuf[3874] = 256'h30dde7dd2edef0dea7df4ee067e173e267e384e491e53fe6dde6a6e75de863e9;
    decBuf[3875] = 256'h57ea34eb37ec2bedc9ed92eee1eef8eee3eea8ee2beedaed90ed4ded59ed64ed;
    decBuf[3876] = 256'h5aed63ed4aed07edd9ec8fec49ec40ec38ec6cecd3ecb1edcdee27f06bf192f2;
    decBuf[3877] = 256'hebf330f557f64af826fa52fc88ff8602060650092a0dc91014141317921aec1c;
    decBuf[3878] = 256'hea1fa322d125d028882bb72eb531a733203617378d3859399739cf39683a963a;
    decBuf[3879] = 256'h693bdc3bff3b5e3c7a3c2c3cb53b493b4a3a9c393d397438593842380138ed37;
    decBuf[3880] = 256'hdb3749370e37b536433617363f36943639379d38ce3a6f3d333f73417e43d244;
    decBuf[3881] = 256'h83469b470049e849634bc84cb04dd74e974fba4f5b4f924e3e4df94bd649ca47;
    decBuf[3882] = 256'hee454743ce408e3e583b5938da349e307f2b0d286a221c1d4a18a8125a0d8708;
    decBuf[3883] = 256'h2504290089fc4ef852f4b2f077ec9ee908e7bde39ae1a8dfe4dd48dc68db9cda;
    decBuf[3884] = 256'he3d93ad907d936d960d9d3d93cdadada6adbecdb63dccfdc31dd67dd98dd89dd;
    decBuf[3885] = 256'h96dd72dd51dd33dd17ddffdcd9dcc5dc99dc71dc4edc08dc9adb15db75dab2d9;
    decBuf[3886] = 256'h2fd989d81dd809d8f7d749d8ebd8d9d9f5da4fdcf0dde9df4de232e5eae719eb;
    decBuf[3887] = 256'h17ee97f1e1f4bbf851fb9cfe75020c054709200cbf0f0a13e416831ace1da721;
    decBuf[3888] = 256'h3e247928522be82d333156330f36d3376f394f3aa33bd83c803d193e473e723e;
    decBuf[3889] = 256'h983e2f3ed03d073d1c3c3f3b023adc388237e1355834f332ae313330342ff02d;
    decBuf[3890] = 256'h1d2d102cd62ab029a3286927422682258e24f0236023a922d421442159203c1f;
    decBuf[3891] = 256'h7c1e881dab1ca81bb41ad719d4185417ef15ab14db12af10a40ec80c9c0afc07;
    decBuf[3892] = 256'h82054203a20073fd50fb97f869f56af2b2ef83ec60eaa7e72ee5eee2e3e007df;
    decBuf[3893] = 256'hdbdc3ada76d836d6c0d4e4d2afd197d098cf0dcfe3cebccedfceffce1bcf36cf;
    decBuf[3894] = 256'h1ecf08cf1ccf0acf1acf81cfdfcf7dd06bd109d20bd300d4ddd4a6d5c6d685d7;
    decBuf[3895] = 256'h7ad896d9a3dadddb04dd10debfde5ddfb3df01e078e0b9e01be198e1c9e130e2;
    decBuf[3896] = 256'h8ee2e3e272e322e4c9e4b6e594e65de77ce889e9c3ea96ebefecd7eda9eeb6ef;
    decBuf[3897] = 256'haaf088f18af27ef39bf441f65af725f9d5fa5efc5dfda2fe74ff34009d00fc00;
    decBuf[3898] = 256'h52016c0184019901ad0130019e00edffe8feaefddbfccffb95fa6ef914f873f6;
    decBuf[3899] = 256'heaf485f387f1abeffbed72ec0debc8e9f6e836e887e7aae61ae62fe591e401e4;
    decBuf[3900] = 256'h4ae3d4e2bee2aae2e0e231e399e3f6e37ce4d5e426e58de5b6e5c2e5e3e5b1e5;
    decBuf[3901] = 256'h83e58be566e543e518e5c3e40de422e345e242e14ee031df25de31dd14dc54db;
    decBuf[3902] = 256'ha6dac8d939d982d8acd7a9d6fbd51ed51bd46cd38fd2ffd1b1d13ad1f9d00dd1;
    decBuf[3903] = 256'h1fd170d1f5d14ed2e0d291d308d49fd477d540d62bd787d8ccd99bdbd0dc59de;
    decBuf[3904] = 256'h58df9de0c3e1d0e20ae485e5eae68be814ea79eb61ece0ec53ed30edd1ec41ec;
    decBuf[3905] = 256'hbfeb48eb07ebccea4feafee979e9b4e8fde7f8e6bee5ece4dfe376e318e334e3;
    decBuf[3906] = 256'hb7e3bce4f6e571e7d6e81bea96eb61ed8def98f10cf557f830fcd9003a053709;
    decBuf[3907] = 256'hdf0d0011fd149c18d71cb01f59247a27762b162f51332a36c038293a723b9c3c;
    decBuf[3908] = 256'hf73c493dfe3c423d053d3d3d0a3ddb3c093caf3a6b39f037bf354934f532c031;
    decBuf[3909] = 256'h1831e5301331923105322832c6321c336a33403443357d364c38783a833ce73e;
    decBuf[3910] = 256'hcb41bd433646d2474749234b584c714dd64e775090515b531454bc548954fe53;
    decBuf[3911] = 256'hd7523151384fd44c944af4477a453a4304402b3c8b385034302f5d2afc25dc20;
    decBuf[3912] = 256'h091ca7178812160fb40ab8060f02eefef2fa52f708f4e4f12cef67ed27ebb2e9;
    decBuf[3913] = 256'h5ee8a4e7fce6c9e69be619e73fe7a8e707e897e819e9c0e92ceab5ea32eb83eb;
    decBuf[3914] = 256'hebeb48ec6dec4cecf2eb3ceb51ea73e937e810e7b7e515e48de228e1e3dfbcde;
    decBuf[3915] = 256'hafdd76dc4fdb42da08d936d876d753d733d789d775d891d9ebda8cdc15de7adf;
    decBuf[3916] = 256'h78e154e3fbe575e8fdeb48ef22f3c1f6fcfaf9fe9802e305bc095c0db60f8f13;
    decBuf[3917] = 256'h2f17791a781d30205f235d264f28c82a642cd92da52eda2f82301b31a7312532;
    decBuf[3918] = 256'he5324d33ec33423490347834633428348733f0323f326931da3023304d2f842e;
    decBuf[3919] = 256'hcd2dc82c192c7b2bb22a2f2a8929f228b7285d280c28e0279d27602755274b27;
    decBuf[3920] = 256'h54277e27762754271c27ab261926b7251625aa244824a723e4222d22c920fe1e;
    decBuf[3921] = 256'h4e1d551b79194d1742156613b5114c0f0c0d6b0a3d073e04860157fe59fba0f8;
    decBuf[3922] = 256'h72f54ef396f01cee81ec76ea12e877e601e5ade378e2d0e137e108e133e1a6e1;
    decBuf[3923] = 256'h54e231e3c1e378e41ee5b6e566e60de7fae7d8e8dbe914eb3bec48ed3ceedaee;
    decBuf[3924] = 256'h30ef7fef97ef81ef6def5bef2bef1ceff4eecfee98ee52eeeeed76ede3ec5aec;
    decBuf[3925] = 256'h24ec14ec23ec81eceeec37ed7aed9fed94ed9eeda7edafedf3ed45ee92ee14ef;
    decBuf[3926] = 256'hb5ef21f0d1f078f13af2f1f2c7f357f40df5b4f54bf6fcf6a2f765f850f92dfa;
    decBuf[3927] = 256'h30fbdefbbcfc12fd94fd0bfe21fe5cfe91fea2fe93fe85fe18fe76fdb3fc94fb;
    decBuf[3928] = 256'h3bfa99f810f7abf50af411f235f085eefcec97eb52ea2be91fe870e793e690e5;
    decBuf[3929] = 256'h9ce4bfe3f5e23fe2c8e15ce16fe15de18ee1f5e11ee242e28fe2c1e213e3b8e3;
    decBuf[3930] = 256'h8ee491e5cae6f1e74be933eab1ead7eafaea9bea45eaf7e950e9e4e834e85ee7;
    decBuf[3931] = 256'h95e6aae58de480e38ce2afe1ace0fedfe1ded4dd26dd49dc7fdb31dbbada4eda;
    decBuf[3932] = 256'h62da2cda5ddaa7daeada57dbf9db90dc1adddedd61ded8de44df7fdfd8df6ae0;
    decBuf[3933] = 256'hf4e095e182e221e3eae3d5e434e5c4e546e68de6fae683e7dce72ee877e84fe8;
    decBuf[3934] = 256'h13e8b0e71ce793e63ae609e635e6aee6ffe666e78ee721e77fe666e50ce4c8e2;
    decBuf[3935] = 256'hf5e182e15fe17fe1d5e123e23be27ce2dee25be30ee472e53de7e4e913ed11f0;
    decBuf[3936] = 256'h58f454f8f4fb3eff1803ae05f9081c0bd50d031102144818451ce41f2024f826;
    decBuf[3937] = 256'h982a012c242e163025311c32fc32c83382342a35c3359535c2346933c7313e30;
    decBuf[3938] = 256'hd92e4e2ed02daa2dcc2d2b2e0f2e292ee12d1f2d9c2c552ce92b4b2c572db02e;
    decBuf[3939] = 256'haf308b32b634c2369e38d2395b3bc03c623e5b40374262446e464a48fa49134b;
    decBuf[3940] = 256'h464bba4a3c4a96480d47dc44d142f540c93ebe3ce23a3b38c1353832ee2e142b;
    decBuf[3941] = 256'h752739233d1f9e1b53185415d5118a0eb10a1107d602dafe31fa10f737f4a1f1;
    decBuf[3942] = 256'h38f014eeeaecdaeb3fea5fe90be8d6e62de694e5c3e5ede560e6c9e667e7bde7;
    decBuf[3943] = 256'hd7e7efe730e86be8c4e815e95fe9bde9e1e9c0e97ae9f1e8f2e7b8e691e5ebe3;
    decBuf[3944] = 256'h62e2fde0b9df92de38ddf4db79da14d92cd805d7f8d590d5f2d4d5d423d5c9d5;
    decBuf[3945] = 256'he3d63cd8ddd9d6dbb2dddedfe9e1d5e48ee7bcea96ee35f271f66dfa0dfe4802;
    decBuf[3946] = 256'h4406db08160d1211b214ed18c61b651fb022d424fe250e276027ab27ef27b127;
    decBuf[3947] = 256'h7927e026552682252924e42269210420621e4a1de51bfd1a2a1a6a19bc181e18;
    decBuf[3948] = 256'h8e170c176516ce1593155d158e159d15c5153216b7167c1767188319dd1a211c;
    decBuf[3949] = 256'hf41c011eaf1e4d1fa31fbd1f471faf1eff1df91c051ce91adc195c185d171916;
    decBuf[3950] = 256'h9e149f13fd110410280e810b52082f067603fd00bdfeb2fc4efa0ef86df5f4f2;
    decBuf[3951] = 256'h10f057ed93eb53e9dde711e758e6b0e517e58be40de4e7e3c4e3e3e33ae4f1e4;
    decBuf[3952] = 256'hf6e530e757e863e99dea70eb30ecdeec7ced0ceec3ee69ef00f0b1f028f1bff1;
    decBuf[3953] = 256'h21f233f202f29bf1edf0e8eff4ee98ed53ec2cebd3e9ebe8c4e7b8e6c4e525e5;
    decBuf[3954] = 256'h5ce4a5e32fe3c2e2afe2e4e236e39de330e492e433e5f6e5e1e63de8dee967eb;
    decBuf[3955] = 256'h32ede2ee6bf036f2e6f36ff5d4f619f840f999fa3afc53fdb8fefdff7b00ee00;
    decBuf[3956] = 256'hcb00eeffebfeb1fd36fcd1fa30f917f8b2f66ef547f4edf2a9f12ef0c9eee1ed;
    decBuf[3957] = 256'h0eed4eece6eb87eb6aeb1cebd4ea93ea80ea4aea3aea2bea03ea0fea46eaa0ea;
    decBuf[3958] = 256'h56eb0dec12ed06eee4eeadef64f03af103f2baf28ff359f4dbf452f568f57bf5;
    decBuf[3959] = 256'h46f5d4f44ff4d2f340f3b6f281f20ff2a8f14af1c5f024f061ef76ee5aed9aec;
    decBuf[3960] = 256'ha6eb89ea7ce942e8c7e662e51ee4a3e2a4e1bce03de017e080e0dee06ee188e1;
    decBuf[3961] = 256'h71e130e1cee074e084e0cee061e188e2afe308e54de673e780e82ee9cde923ea;
    decBuf[3962] = 256'h0eebebebeeec28ee4fef0ff003f122f106f183f04eef27ee81ecf8ea2de9f9e7;
    decBuf[3963] = 256'he0e647e65fe538e4dfe29ae1cbdf1bde22dcceda99d9f0d857d829d853d82dd8;
    decBuf[3964] = 256'h0ad8ead794d7aed7f5d7b8d80cdaaddb16de56e08ce3b0e52fe989eb88ee40f1;
    decBuf[3965] = 256'h6ff46df7edfa37fe1102b0050a08090bc10d3b107b121b159517d519751c3a1e;
    decBuf[3966] = 256'h7a20852261249625ae264727d2275128c428e72846299c29b6299e295d29fb28;
    decBuf[3967] = 256'hc628542845288828f528d229b02ab22ba72cc32dd02ec42fe130ed316d333835;
    decBuf[3968] = 256'h6437043a7e3c623f1b4294442f463b488f49c34a4c4cb14df64e7150d651be52;
    decBuf[3969] = 256'h90536a53015324522151a24fa34e014d784b134a1548b1457243a63f063ccb37;
    decBuf[3970] = 256'hcf33262fc42ac8262022fe1e021b631709150a128b0e310c32097a060004c101;
    decBuf[3971] = 256'h4b007fff4afe32fd99fc54fb81fa75f93bf868f75cf6adf50ff5b9f49ff457f4;
    decBuf[3972] = 256'h17f48df3a5f2c7f18bf064ef0beec6ec4beb4cea08e935e828e7eee573e4a8e2;
    decBuf[3973] = 256'hf8e06fdf0adec6dcf3db33db85da26da09daefd907daf1d92cda62dad3dab1db;
    decBuf[3974] = 256'h0cdd51deccdfcbe010e28be3f0e491e68ae866ea92ec33efacf191f449f778fa;
    decBuf[3975] = 256'h9bfc54ffcd010d04ae06dc09000cb80e321171137d1559170919021bde1c131e;
    decBuf[3976] = 256'h0c206021102329248e25d226a5276528ce28ed280a29f028d828ee280129ef28;
    decBuf[3977] = 256'hbf287528ac27aa267025f5239022a8212921b62093207420572071202a20e91f;
    decBuf[3978] = 256'h871f0a1f571ee01d9f1d3d1d4f1d3f1d6b1dc91d1e1e551eaf1ebb1eb01ece1e;
    decBuf[3979] = 256'hb21e9a1e831e1c1e3f1d221cc91a27199e17d31523149a12cf101f0f960dcb0b;
    decBuf[3980] = 256'h1b0a02099d07590632052504eb0219020c01d2ff00ffa6fd62fc8ffb36faf1f8;
    decBuf[3981] = 256'hcaf70af7a2f643f65ff67af6c1f62df78ff7e8f75af8c1f804f929f960f96af9;
    decBuf[3982] = 256'h4ef925f9d3f85af8c7f73ef79df606f6a4f56ef53df511f504f510f5d9f493f4;
    decBuf[3983] = 256'h1cf469f394f2caf113f19df031f0a7ef2aefd9ee37eecaed90ed5aed4aed58ed;
    decBuf[3984] = 256'h4bed3fed60ed6aed85edd0eddaede3edfbede5edd0edd7edbaedabed9ded66ed;
    decBuf[3985] = 256'h13edc6ec44ecc7eb56ebd1ea77ea47ea1aea0dea01eab4e95ae9ede84be8b3e7;
    decBuf[3986] = 256'h2ae765e6e3e53ce54ee471e3e1e22ae284e143e1e1e0ace09be08de07fe08be0;
    decBuf[3987] = 256'hace0dee043e1a0e126e2eae26de3e4e3a6e429e5cfe592e67de79ae8a6e99aea;
    decBuf[3988] = 256'h38eb02ec50ec97ec03ed66ed9bed0dee1ceef4ed9fedfaec24ec21ebe7e9c0e8;
    decBuf[3989] = 256'h67e722e6fce43ce448e3e9e292e244e22ce26de281e2b6e208e334e35ce3b1e3;
    decBuf[3990] = 256'hbce302e454e4a1e4fbe468e5cfe548e6bae621e799e72be8b5e879e965ea03eb;
    decBuf[3991] = 256'hcceb4fecc5ec06ed68ed9eedcfedfbedeeedc9ed92edfcec3aecb7ebe1ea18ea;
    decBuf[3992] = 256'h95e9efe883e86fe816e8c5e77be7cde627e639e55ce41fe3f8e1ece0b2dfdfde;
    decBuf[3993] = 256'hd3dd6add0bddeedc09dd20dd8cdd3dde13df4fe0cae12fe3d1e459e6bee760e9;
    decBuf[3994] = 256'h59eb35ed61ef01f27bf4bbf6f1f9effca8ffd602b0064f0a9a0d991018146317;
    decBuf[3995] = 256'h611a531c811fa52196231026ab272129752aa92b522ceb2c192d432d1d2dfa2c;
    decBuf[3996] = 256'hda2cf72ca92cc12cd62cc32cd42c052dd92ce62c3b2d5c2dde2da32e8e2fea30;
    decBuf[3997] = 256'h8b328434e8362839333b973dd73f4d4129435545ca462e496e4b794d554f0651;
    decBuf[3998] = 256'hae514752195246513950ff4e844d1f4c7e4a8548a946f9448f42ab3ff23cc439;
    decBuf[3999] = 256'hc5367f32a62f072cbc289926e023b220b31dc21b93189515dc12f90e620c1709;
    decBuf[4000] = 256'hf4063b047702dc0066ff9afe65fd4dfcb4fb28fbaafa84fa61fa41fa5efa10fa;
    decBuf[4001] = 256'hf8f98cf902f93ef853f736f6ddf498f31df21ef136f063efa3eef5edd8ec7feb;
    decBuf[4002] = 256'h3aea6be8bbe632e567e3b7e12ee063deb3dcb9da65d9b5d79dd69ed512d594d4;
    decBuf[4003] = 256'h6ed4d6d435d5fed5ead606d8acd9a5db81dd29e0ede12de438e614e840ea4bec;
    decBuf[4004] = 256'hafee4af056f2baf4f9f69af914fcf8fe7702d104d007880a020d9d0e1310df10;
    decBuf[4005] = 256'h981140127312ff12d11344146714871431147a13a412db112411ad106c10a710;
    decBuf[4006] = 256'h001193111c129912ea12f9120713e21295123b12ce114911a8101110880fe70e;
    decBuf[4007] = 256'h4f0e9f0dc90cc60b180b7a0a5d0a770aee0ab10b330c7a0c650c030c1a0bfe09;
    decBuf[4008] = 256'ha4086007e505e6045a04dc03b603d903f8034e049d04b504ca04b704a5049404;
    decBuf[4009] = 256'ha304cb04d704a00432045503f90158005ffefbfbbbf945f869f635f58cf459f4;
    decBuf[4010] = 256'h2bf455f47bf4e4f443f526f5d8f431f444f327f21af1e0efbaeefaed91ed32ed;
    decBuf[4011] = 256'h4fed69ed81ed96edaaedbcededed54eee7ee98ef6df037f1b9f101f241f255f2;
    decBuf[4012] = 256'h43f2f2f16df1a9f0f2ef4befb4ee2beef5ed05ee4feec7ee5aef0af052f03cf0;
    decBuf[4013] = 256'h01f0a8ef36ef0aefe2eebdeeb2ee6cee3fee47ee3fee6feec1eef8ee3eefc7ef;
    decBuf[4014] = 256'h50f015f100f2ddf2e0f38ef4edf443f55df516f5aaf421f438f35bf258f164f0;
    decBuf[4015] = 256'h87efbdee07ee90ed24edc2ecb0ece0ec0deda0ed50ee26efb6ef6df0b4f0caf0;
    decBuf[4016] = 256'h8ff0eeef2bef40ee63ed60ecf7eb59eb03eb1deb35eb4beb5eeb29ebf8eaccea;
    decBuf[4017] = 256'ha3eac8ea57ebe0eba5ec5cedd2ede8edfcedc6ed54ededec3fecc8eb88eb9beb;
    decBuf[4018] = 256'hf5ebc8eccbed04ef80f0e5f1ccf29ff379f310f333f230f1b0efb1ee10edf7eb;
    decBuf[4019] = 256'hf8ea10ea3ee97ee8d0e771e71ae700e7e9e655e790e70de89fe801e95ae9cce9;
    decBuf[4020] = 256'hbde97be956e9c7e83ee808e896e76ae75de769e7a0e722e8c3e85ae932ea88ea;
    decBuf[4021] = 256'hd7eaeeeaaeeac1eaf7ea28eb8febeceb11ecf0eb96ebe0ea29ea24e930e813e7;
    decBuf[4022] = 256'h06e612e574e4abe328e3b2e29ce2b0e2e5e257e3bee337e4a8e42de515e632e7;
    decBuf[4023] = 256'h8be88aea66ec0def86f16bf423f752fa50fdd0001a041907d109000dfe0fb712;
    decBuf[4024] = 256'h30151418cd1a461d861f91216d231e25a7260c28f3286f2ad42bbb2ce22d3c2f;
    decBuf[4025] = 256'h2430f630b6311f327e329a324c32053299310f31fd30ed30de3021318e31bb31;
    decBuf[4026] = 256'h3332c5324f33373454356036e037ab395b3be43caf3ee43ffc40fb4186425943;
    decBuf[4027] = 256'hb24454464d48294a554c604eb44fe9509151c4513951bb50614f634d874b5b49;
    decBuf[4028] = 256'hbb46f6441242923e483b4938ca347f31a62d062abb2698241821af1fb11cbf1a;
    decBuf[4029] = 256'h46180616d012d10f520c0709e4062b046702cb0056ff02fe48fda0fca1fbb9fa;
    decBuf[4030] = 256'h3bfa7bf958f978f994f9e3f92afa40fa7bfa45faf4f98cf9c4f8fbf744f79df6;
    decBuf[4031] = 256'h31f6f6f5e5f5d4f5a8f515f53df43af3bbf1f0ef3feeb7ececea3be9b2e74de6;
    decBuf[4032] = 256'h66e5e7e4c1e49ee4bee4dae4f4e43ce5d3e5abe6e7e762e92debdeec66ee97f0;
    decBuf[4033] = 256'ha3f207f546f752f9b6fbf5fd0100650200040b06e707130a1e0cfa0daa0fa411;
    decBuf[4034] = 256'h80133015b916b817fc18cf19421a651a851af5193e193918ff16d815cb14d713;
    decBuf[4035] = 256'hfa12311245116810d80f210f4c0e820d630c0a0b220a4f09dc08b90818093509;
    decBuf[4036] = 256'h1b09a4080d0835076b06b5053e0528058a052b064407ea08e40ac00ceb0ef710;
    decBuf[4037] = 256'h4b127f13b713ea13bc133e13cb121c127e112811d91092102610eb0fb60f640f;
    decBuf[4038] = 256'h380ff50ea00e3d0e8f0d8a0c0b0ba609a707cb05a0039401b8ff8dfd17fcc3fa;
    decBuf[4039] = 256'h13f96af86bf783f605f645f5ddf4bdf413f562f508f69ff629f782f7d3f71df8;
    decBuf[4040] = 256'hb0f861f936fa39fbe8fb86fc15fd64fdabfdc1fdadfd54fd02fd9bfc3efc01fc;
    decBuf[4041] = 256'he0fbc2fbb9fb5efbc0fad3f977f879f69df471f266f08aeed0edb8ec85ec56ec;
    decBuf[4042] = 256'hd8eb18eb24ea47e97de8c6e750e70fe7fbe6c6e6d6e602e70fe74ce741e7fbe6;
    decBuf[4043] = 256'h97e6e9e543e502e5eee424e5b6e567e63ce706e820e837e84de812e8dde7ede7;
    decBuf[4044] = 256'hfce73ee863e858e83ae831e8d6e781e708e755e6dfe59ee53ce52ae53ae52be5;
    decBuf[4045] = 256'h03e5f7e4aae450e4e3e323e338e29ae1d1e082e09ae0b0e0eae044e195e1dfe1;
    decBuf[4046] = 256'h72e223e3f8e335e507e614e74ee820e92dea21ebfeebc8ec7fed25eee7ee9eef;
    decBuf[4047] = 256'h74f077f1b1f2d8f3e4f4d8f5b6f645f794f7acf76bf709f720f604f5aaf309f2;
    decBuf[4048] = 256'h80f0b5ee89ec13eb37e903e87ae67be593e415e43be418e477e407e521e568e5;
    decBuf[4049] = 256'h7ee56ae558e548e51ce50ee563e5f2e5cae606e82de9d3ea5cec5beda0eec7ef;
    decBuf[4050] = 256'h3af0a2f0c2f0a5f057f03ff02af0efefb9ef47efa5eee2ed2ced56ec8debd6ea;
    decBuf[4051] = 256'hd0e9dce8ffe76fe7ede6a5e6bbe6f6e673e705e88fe82fe9c7e977ea1eebe0eb;
    decBuf[4052] = 256'hcbeca9edaceea0effcf09df296f4faf6def997fc5bfe40013103f60491060708;
    decBuf[4053] = 256'h5b09860bfc0cd80e04110f137315b317be199a1bc61d3c1f9020492181214e21;
    decBuf[4054] = 256'h7c21a6211a22c82266232f24e6245d25c9257a26f0268827ea27fc27ec27bf27;
    decBuf[4055] = 256'h9727d4274d28df28b729802a6b2b492c4b2dfa2dd72ea02f57302d31f631e132;
    decBuf[4056] = 256'hfe330b35ff355b379f38c639d33a0d3cdf3c9f3dc23da23d4c3d953c613be539;
    decBuf[4057] = 256'h80388236a6347b326f300b2ecc2b2b29fc25fe224520cc1de81a2f18b6157613;
    decBuf[4058] = 256'h6b111710eb0d750c210bec09d408d507900669055d04dd02de01f6002300b0ff;
    decBuf[4059] = 256'h48ff6afea1fdeafc14fc85fb02fb5cfaf0f98ef910f95ef8b7f7caf6ecf523f5;
    decBuf[4060] = 256'h38f45af3cbf214f29df106f17cf0ffef8def09ef8cee1aee95edd0ec1aec44eb;
    decBuf[4061] = 256'hb4ea66eaadea19ebcaeb70ecdcec3eed74eda5edeeed31ee6eeea5eeebee61ef;
    decBuf[4062] = 256'hf4eff3f0e7f143f32bf4fdf4bdf526f685f6dbf692f797f8d1f94cfb17fdc7fe;
    decBuf[4063] = 256'hc0001402ce027603a9037b0351032a030703e8023e035803cf033b04c4041e05;
    decBuf[4064] = 256'h6f059b05a9059c057b054905e5045204c9036f03dd02a2024902180209021702;
    decBuf[4065] = 256'h3b028802f6025d03d603270471049904a504b004e2043405d905af06eb071209;
    decBuf[4066] = 256'hd209800adf0ac20a740afd093a09b808e20719072e06500587040404bd037c03;
    decBuf[4067] = 256'h69033303e2027b02e7015e01e1006f00eaff6dfffcfeb2fe6ffe32fe3dfe5bfe;
    decBuf[4068] = 256'h9bfee5fe3fff94ffe1ff130041005a0070009300be0007014d017b0194017d01;
    decBuf[4069] = 256'h2401b700150052ff67fe89fd4dfc7bfb6efa05faa6f98af9a4f9ebf9d5f973f9;
    decBuf[4070] = 256'hf6f823f85af7a3f6cdf504f519f43bf339f244f1a6f017f0fcef14f0ffef39f0;
    decBuf[4071] = 256'h4bf05cf04df025f0d0ef6defdaee50eed3ed61edfaecd2ecaeecb9ecd7ec17ed;
    decBuf[4072] = 256'h50ed94ed8bed40edd2ec30ec99eb5eeb28eb39eb82ebaaebe7eb1eec28ec1fec;
    decBuf[4073] = 256'h27ec11ec0aec1dec2dec5cecadece4ec16ed56ed3ded17edccec5eecd9eb80eb;
    decBuf[4074] = 256'h0eebc4ead2ea0eeb9deb4eec24ed26eed5ee73ef03f01df005f0c4ef62ef09ef;
    decBuf[4075] = 256'hd8ee04ef62efffefedf0cbf107f382f4e7f52cf7fef771f894f8b4f85ef843f8;
    decBuf[4076] = 256'hfcf790f72ef7d5f683f675f682f6bff638f7a9f711f853f878f841f8d3f74ef7;
    decBuf[4077] = 256'h89f607f6c0f5d5f537f6d8f670f720f8c6f85ef90efa85fac6fab2fa59fae7f9;
    decBuf[4078] = 256'hbbf9c8f936fa13fb2ffceffce3fd42fe26fea3fdcdfc04fc4dfbd6fac1fafcfa;
    decBuf[4079] = 256'h55fbc7fb10fc39fc45fc3afc44fc4dfc34fc00fc98fbf6fa34fab1f96af97ff9;
    decBuf[4080] = 256'hbaf914faa6fa2ffbacfbfefb47fc8afc96fc8bfc81fc54fc09fcaffb5bfb24fb;
    decBuf[4081] = 256'h56fbccfbc0fcfafd75ffda00c201e9025c03c403e40301041b0433047404fd04;
    decBuf[4082] = 256'h7a054d0650078a08b109570be00c450ee60fff10fe11e612b8132b142015be15;
    decBuf[4083] = 256'h871672171018d9185c19a319b919cd199719a719f1194f1aec1a841be61b3f1c;
    decBuf[4084] = 256'h901cda1c1d1d721dbf1d2d1eb21e521f152034214122c12326256a26e527e428;
    decBuf[4085] = 256'h13293d291729ae2810288027fd26e626d026e4266127d3271c287a289e286728;
    decBuf[4086] = 256'hf92757276926cb25c8241a247c23b3223022b92122214a20811f611e081d201c;
    decBuf[4087] = 256'hf91aed193e19df188918a3188b184b18e81748170316bf149b129010b40e030d;
    decBuf[4088] = 256'h7b0b7c0a940915093c095f097e09d409230adc099b0911090508f90679051404;
    decBuf[4089] = 256'hcf0254015500cafff7fed1feaefecefeb1fecbfee3fea2fe8efe35fec3fd97fd;
    decBuf[4090] = 256'h54fd30fd0ffdf1fcc3fc9afc65fc0cfcb7fb28fb78fad1f93af9b1f857f847f8;
    decBuf[4091] = 256'h56f8b3f820f9c3f95afa0bfb81fb19fc7bfcd4fc26fd8dfd05fe77fefcfe79ff;
    decBuf[4092] = 256'hebff6f00a500f60005012d016a01a101fb016802ed024603b8031f0462046e04;
    decBuf[4093] = 256'h4d04cb03e302c601b9007fff59fe99fda5fc06fc77fb28fb70fbdcfbb4fcb6fd;
    decBuf[4094] = 256'hf0fe17007001b502dc034f047204d40398021c0151ffa1fd18fc19fbd5f956f9;
    decBuf[4095] = 256'h30f953f972f9c9f94bfac2fa03fb8cfbe6fb37fc63fc71fc34fcd1fb3efb66fa;
    decBuf[4096] = 256'h9df9b2f895f788f6daf57bf55ef5adf553f641f75df86af918fab7fa0dfbbefa;
    decBuf[4097] = 256'h77fa89f9acf870f749f6a3f48af3bff18af0e2efe3eeb5ee8aee64eecdee2cef;
    decBuf[4098] = 256'h48ef97efdeefc8ef66efc5ee81ede0eb57eaf2e850e7c7e562e41ee34be23fe1;
    decBuf[4099] = 256'h90e0f2df9cdf19dfd2de91dea5dedade0bdf55df7ddf59df22dfc8de42dea1dd;
    decBuf[4100] = 256'h0add81dc27dcf6db23dc9bdc6eddfeddb5de5bdf9cdffedf34e085e0ece09ae1;
    decBuf[4101] = 256'h11e2d4e28ae331e4c8e451e563e512e5abe418e48ee359e348e392e30be47ce4;
    decBuf[4102] = 256'he4e441e566e59de5f7e533e6ace61ee785e7e3e707e8d0e78ae726e7c8e68ce6;
    decBuf[4103] = 256'hade61be7f8e754e9f5eaeeec52efedf0f9f24df481f52af6c3f6f1f61bf78ef7;
    decBuf[4104] = 256'hf7f756f81ff9d6f97cfa14fb4ffba8fbd9fb40fceefcf3fde7fe43002b01fe01;
    decBuf[4105] = 256'hbd02e0020003aa025b021402fe01120224027502a102ca02ee0225035703a903;
    decBuf[4106] = 256'h0c048404f6047b05f8054906760683065f062806f605c805af05b705cb05eb05;
    decBuf[4107] = 256'h1d066906c3061807390743072707ee06c806c106ed064107ae07160859087d08;
    decBuf[4108] = 256'h5c0802086407a206b705d9044904fb0384034303e1024002d4014b0115010501;
    decBuf[4109] = 256'h14013c0160019701dd015402e60297036d04fc047f05f6053706710683065306;
    decBuf[4110] = 256'h0906e105d5050c06a20664074f086c092c0a200b3d0cb00c5e0dbd0dda0dc00d;
    decBuf[4111] = 256'ha80d100dd60ca00c900cbc0c340da60d660e1d0f930f00103a104c107d108c10;
    decBuf[4112] = 256'h9910be100b1129117b11c8110e12841217137913f61368149414a11495148a14;
    decBuf[4113] = 256'ha8140c15851538160d17d7178d186319f319aa1a501bbc1b461cc31cf31c5b1d;
    decBuf[4114] = 256'hd31d451e051fbb1f62202421db212222ba22f5222a233b2367233f234b234023;
    decBuf[4115] = 256'h5e23b02313245624c3240d25ff24db2462248f23c522da21fd20a72024200c20;
    decBuf[4116] = 256'h22200e20fc1f0d20e01fd31fdf1fa81f121f241ec81cca1a76194b17d5158114;
    decBuf[4117] = 256'h4c13a4120b12801155117c1159113911e3106010ba0ff80ed80d7f0cdd0a5509;
    decBuf[4118] = 256'hf007ab06d8056505fd04dd04870404045e0370029301c9001200cbff8aff9eff;
    decBuf[4119] = 256'hd4ffc3ff7aff1cff66feaffdd9fcd7fb9dfacaf9bef80ff8b0f7cdf71bf8c2f8;
    decBuf[4120] = 256'h84f93bfab2fac8fa65fa7df921f880f6f7f4f8f310f392f21ff2b6f157f101f1;
    decBuf[4121] = 256'hb2f06bf02af017f029f039f048f070f07cf09df093f09cf094f07df069f056f0;
    decBuf[4122] = 256'h0df09fef37efdaee9deebeee04ef7befedef36f079f0b6f0d7f0e1f0eaf0c1f0;
    decBuf[4123] = 256'h8cf085f073f083f0bcf0f0f020f14cf152f157f152f113f1d3f099f037f00ff0;
    decBuf[4124] = 256'hebefcaefd4ef02f02bf06ef0aef0c7f0b0f065f0cfef0cef8aee13eefded5fee;
    decBuf[4125] = 256'hb9ee4befd4ef51f0c3f048f1a1f154f22af3f3f3aaf450f5bcf5d0f577f5c4f4;
    decBuf[4126] = 256'hbff310f333f2ddf1c2f139f2d1f281f327f468f4a3f44af497f392f258f1ddef;
    decBuf[4127] = 256'hdeeef6ed78ed9eed07ee65eef5ee0fefc8ee31ee0aede3eb8aeaa2e9d0e8a9e8;
    decBuf[4128] = 256'hcce82be9f4e9abea22eb63eb76eb64eb75eb83ebe1eb4eecb5ecf8ec65ed92ed;
    decBuf[4129] = 256'hefed75eef2ee64efe8ef42f093f0faf008f1fbf0f0f082f0feef5def6fee92ed;
    decBuf[4130] = 256'h02ed7fec38ec22ec5decb7ec28ed72ed7fed73ed10ed7decf4eb0beb6dea17ea;
    decBuf[4131] = 256'hc9e910ea7cea05ebcaeb81ec27ed93edf5ed07ee38ee64eea7ee14efb7ef4ef0;
    decBuf[4132] = 256'hd7f054f1a6f10df285f2f7f2b7f3a2f4bff5cbf605f8d8f8e4f993faf2fa48fb;
    decBuf[4133] = 256'h96fbddfb4afcacfce1fc33fd7cfdbffdfcfd49fe7bfebbfe05ff73fff8ff9900;
    decBuf[4134] = 256'h3001e1018702f3022e0340032f0321032e033a039d031604a8045805ff056b06;
    decBuf[4135] = 256'hcd06bb06cb06da061d07a20767088609e00a240cf70cb70d1f0ec10d6a0de80c;
    decBuf[4136] = 256'h410c2c0c8e0c2f0d1d0efa0efd0fab10cb10ae106010b90fcc0eee0db20c8b0b;
    decBuf[4137] = 256'h7e0ad009710954093a0982099709ab09bd09ac099e09ab09b709c209e009fc09;
    decBuf[4138] = 256'h140afe09f709e409d309ed09290a940a370bce0b570cd40c460d720dd00df40d;
    decBuf[4139] = 256'h150ef70da50d000d5a0c6c0b8f0aff097c0906091b097d09fb09ee0ae20b810c;
    decBuf[4140] = 256'h4a0dcc0de40dfa0dbf0d420df10ca70c490c3d0c5e0c680c960cbf0cd50c210d;
    decBuf[4141] = 256'h7b0de80da80e930f311034112812c6128f13de13f6130b14f813c213d213fe13;
    decBuf[4142] = 256'h4114df14a2158d16a9170319471a6e1b7b1c291d881dde1dc41dac1d6c1d311d;
    decBuf[4143] = 256'h1f1d501d991d2c1eb61e331fe61f8c20f820a9211f2260229b226622f4215221;
    decBuf[4144] = 256'h8f20a41f061f761ef31dac1d6b1d301d1e1d0e1dff1c421d7f1dcc1d261e4a1e;
    decBuf[4145] = 256'h3f1e491e2e1e051efd1de91dbd1da11d541daf1c091c1b1bfe193e1904183217;
    decBuf[4146] = 256'h7216c315e614e313ef12d311c6108c0f650ea50db10cd40b0b0b1f0a4209b208;
    decBuf[4147] = 256'hfb0755071407d906c806d806c9066b06e605fe04e103d4029b01740067ffb9fe;
    decBuf[4148] = 256'h1bfec4fdaafd92fd52fd17fd76fcb3fb94fa3af999f7a0f5c4f38ff206f1a1ef;
    decBuf[4149] = 256'h16efeceec6ee2eef8def1df06bf0e2f079f1b4f1c6f1b6f131f16df081ef65ee;
    decBuf[4150] = 256'h0bed24ec51ebdeeabbeadbeaf7ea7aebc1ebd7ebc3eb46eb73eaaae98ae87ee7;
    decBuf[4151] = 256'h89e6ebe595e5afe5f6e58ee63ee714e8dde894e90bea21ea0deab4e921e9e7e8;
    decBuf[4152] = 256'hb1e8c1e846e9e7e9d5eaf1ebb1eca5ed04ee21ee3bee23ee0eeefaed0ceefced;
    decBuf[4153] = 256'h0aee18ee3cee5deeb7ee0cef6fefcdeff1effceff2efc4ef9bef85ef70ef8fef;
    decBuf[4154] = 256'he4ef81f044f12ff20cf30ff403f562f5b8f5d3f5bbf54ff5c5f401f4b2f36bf3;
    decBuf[4155] = 256'h55f3b8f358f4f0f479f51af686f6e8f642f731f723f7fbf6a6f66ff651f635f6;
    decBuf[4156] = 256'h3ef672f6bef62cf7cef791f847f91dfaadfafbfa13fbd2fa22fa1cf9e2f767f6;
    decBuf[4157] = 256'h68f580f4aef33bf318f337f354f36ef386f370f384f372f362f318f3d5f250f2;
    decBuf[4158] = 256'haff1ecf06af0c4ef83ef96efccef5ef00ff1b5f178f2faf2a1f3e1f31cf40af4;
    decBuf[4159] = 256'h1bf40cf4fff3f2f313f445f473f4bdf4eff42ff569f570f577f54cf5f7f48af4;
    decBuf[4160] = 256'h05f488f316f392f215f282f1f9f058f0ecefb1efc3eff4ef78f0d2f044f170f1;
    decBuf[4161] = 256'h7df171f166f170f19ef119f2baf2a8f386f44ff5d1f519f65af6bcf615f7a7f7;
    decBuf[4162] = 256'h31f8aef820f987f9e4f939fac8fa52fbf3fbb5fc38fd7ffd95fda8fd73fd21fd;
    decBuf[4163] = 256'hd8fc95fc89fc94fcdafc50fd03fed9fea2ff8d006b01c1010f02f7018b01b300;
    decBuf[4164] = 256'hb1ffbdfe1efe02fe1cfec2fe59ff3100c1007801ef0130026a02a002b002a202;
    decBuf[4165] = 256'haf02a302ae02e0023203ab033d04ee04940557060e07e3077308f6089c09080a;
    decBuf[4166] = 256'h6a0ae70a7a0bdc0b110c220cf50bb20b5e0bfb0ab80a930a5c0a3e0a350a4e0a;
    decBuf[4167] = 256'h730ab10aca0ab40a760afa095909ed088b0879088908b5082e09c009710a170b;
    decBuf[4168] = 256'hae0b380c910c030d4d0d8f0dcc0ded0de30db50d7c0d740db20d2e0e160f3310;
    decBuf[4169] = 256'h3f1179124c130c147414d314b7146814c2132b137a12d4116811051117112811;
    decBuf[4170] = 256'hac114d12e5129513dc131d140a14b0133f13ba1219128211f810c310b2101a11;
    decBuf[4171] = 256'hc7119d12a0139414f3144915fb1425145c13a5122e124412cd12b613d214df15;
    decBuf[4172] = 256'hd31671178e17a8176117f5166b16361646169016581721180d19291ae91a971b;
    decBuf[4173] = 256'hf61bda1b571b811a7e198a186e17ae16ff156115d2144f14d8136c130a13b112;
    decBuf[4174] = 256'h1e129511f4105d10850ff50e3e0e980d010d290c5f0ba90a020a4009bd087608;
    decBuf[4175] = 256'h6008c2083f09d209820aca0adf0a7d0ab809650820075105a10388028901fe00;
    decBuf[4176] = 256'hd400fa001d017c015f0145019f0086ff2cfe8bfc02fb9df9fcf7e3f6e4f559f5;
    decBuf[4177] = 256'h2ff508f571f5d0f526f674f68cf620f66ff53bf414f36ef155f056efcbee4dee;
    decBuf[4178] = 256'h73ee50eeafeecceeb2ee9aee59eed0ed52edc0ec10ec99eb2debf2ea04eb55eb;
    decBuf[4179] = 256'hdaeb57ec2aedbaed3ceeb3eec9eeb5ee5ceecaed19eda2ec0beca9eb73eb63eb;
    decBuf[4180] = 256'h72ebb4ebf1eb28ec5aec3fec15ece1eb7aeb30eb08eb14eb4bebb9eb3eecdfec;
    decBuf[4181] = 256'h76edd8ed55eea7eef0ee33ef88efbfef19f06ef0d1f064f115f28bf223f3acf3;
    decBuf[4182] = 256'h06f436f480f4a8f4fdf476f508f6b9f65ff7f7f780f8d9f80af954f97cf9b9f9;
    decBuf[4183] = 256'h32faa3fa28fba5fb17fc7efcc1fcfefc09fd27fd30fd07fdd2fc94fc4afc18fc;
    decBuf[4184] = 256'h21fc4afc9dfc16fd67fdcefd11fe05fefafdb4fd62fdfffca1fc4cfcfffbcdfb;
    decBuf[4185] = 256'h8efb85fbabfb12fcd2fcbdfd9afe9dff4b00aa00c700ad0066002500eaffb4ff;
    decBuf[4186] = 256'h63ff19ffd6fe81fe60fe2efe4afe84fec7fe19ff50ff5aff3fff05ff95fe02fe;
    decBuf[4187] = 256'h79fdd8fc6cfc31fc1ffc50fc5ffc6cfc78fc6dfc63fc48fc1ffceafbacfb83fb;
    decBuf[4188] = 256'h5dfb64fb6bfb87fba0fbb7fbc4fbd0fbe1fbfdfb28fc5bfc99fcf3fc60fdc8fd;
    decBuf[4189] = 256'h5bfee4fe61ffb3ff1a00420066005b0051004800400047005c0062005d004300;
    decBuf[4190] = 256'h1900dcff91ff37ffe2fec1fea3fed1fe1bff89ff0e006700d900230130013c01;
    decBuf[4191] = 256'h31011301f80011014501ac014f021103fc03da04a30526066d06ae06e9061e07;
    decBuf[4192] = 256'h4f07990711088308cd0810090309e2089c085d08330859089708f10846096709;
    decBuf[4193] = 256'h4909f70868089007c7061006990559056c05a205f3053d068006bc06dd06d306;
    decBuf[4194] = 256'ha6064b06c6054805d7048d048004a404db0435058a05d7051d065d0665066c06;
    decBuf[4195] = 256'h580645064b065a068406c206fb063f077f07b807de070008fa07c7076e071907;
    decBuf[4196] = 256'ha0066f06430636061106da056c05e80447048403cd022702e601d301e4013602;
    decBuf[4197] = 256'h9d02fb020703fc02b6025102f4019f019401ee018b024e0339041705e0052e06;
    decBuf[4198] = 256'h46063006ce059905270518050b052f05a8051a069f061c076d07b707c407b807;
    decBuf[4199] = 256'h970779073907ff06cb069b066f065e0644061b06e8059d052f05c7046a042d04;
    decBuf[4200] = 256'h22046804cc04600510068706f3062e07f806c80660060306f70502065c06e106;
    decBuf[4201] = 256'ha6075c083209fb097e0ac50adb0ac70ab50a850a930ad60a5c0bfd0bbf0caa0d;
    decBuf[4202] = 256'h480ed80e270f0f0fce0e450e800dc90c230cb70b550b1f0bee0afd0a0a0b2f0b;
    decBuf[4203] = 256'h660b840b7b0b410bd00add09e8088d07a5062606b3059005ef057f063607ad07;
    decBuf[4204] = 256'h190854084208f0076c07ef065c06d3057a0549051d052a0536056d05c7050406;
    decBuf[4205] = 256'h5106ab06cf06da06d00690062506a005ff0468049003c70210026a01a700f0ff;
    decBuf[4206] = 256'h4aff87fed0fd2afd68fcb1fb0afb73faeaf9b4f9a4f9b3f9c0f9ccf9abf965f9;
    decBuf[4207] = 256'heef87df8daf76ef70cf7faf6eaf616f724f730f725f7f3f6a1f654f6faf5bdf5;
    decBuf[4208] = 256'h9cf592f5c0f5f9f54cf699f6cbf6b0f665f6f7f555f5bef40df496f355f369f3;
    decBuf[4209] = 256'h9ff310f495f412f564f590f582f515f591f4ccf315f33ff2b0f12df115f12bf1;
    decBuf[4210] = 256'h66f1bff131f298f2f6f232f353f385f38ef397f39ef397f39ef3aef3c8f3fbf3;
    decBuf[4211] = 256'h47f48df4dff416f548f563f57cf583f598f5c4f5e0f504f624f628f61df604f6;
    decBuf[4212] = 256'hd5f58af558f52af522f529f530f543f549f543f536f529f506f5d3f4a3f45ef4;
    decBuf[4213] = 256'h1ef4f5f3dff3f3f32bf460f49ef4d8f4eef4f5f4e2f4bbf48df461f445f440f4;
    decBuf[4214] = 256'h4ef463f47ef49df499f486f46df445f429f438f458f498f4eaf44df590f5cdf5;
    decBuf[4215] = 256'hd8f5baf58cf531f5c4f47af438f42bf462f4a8f41ff5b1f53bf6b8f62af756f7;
    decBuf[4216] = 256'h63f73ff7f2f698f65bf624f62ef680f6cdf64ff7ccf75ff8c1f83ef98ff9bbf9;
    decBuf[4217] = 256'he4f9d7f9b6f984f945f90bf9e5f8b5f896f86ff84bf834f838f843f871f8a9f8;
    decBuf[4218] = 256'hedf83ff9a2f9fff96dfad4fa17fb53fb74fb92fbc0fbfafb3dfca2fc35fdbefd;
    decBuf[4219] = 256'ha6fe84ff87007b011902e202300348030703cc02970246021902f101e501f001;
    decBuf[4220] = 256'h0e023c028602cc020c0335034c035203400324030a030f0313030703e802a802;
    decBuf[4221] = 256'h4402e601910170018e010502b7028d03900484056106f106400787079c078907;
    decBuf[4222] = 256'h5307430752074407500745074f0759078207d4074d08e0089009070a9e0a000b;
    decBuf[4223] = 256'h360b670b760b680b440b230bdd0a9d0a630a200af209d909b409bb09cd09de09;
    decBuf[4224] = 256'hee09e009ba0996096c095b096b0982099f09b309b609a709a4099c09a309c309;
    decBuf[4225] = 256'he3091b0a6d0ad00a2e0bb30b300c810cae0ca00c4b0ce80b550ba50a2e0a9709;
    decBuf[4226] = 256'h5c094a095a09860994096f090c09af0811087a0718079a064906e2058405ff04;
    decBuf[4227] = 256'h8204f0036603e9025702f5019b012a01e0009d00600055005f007b00a400e700;
    decBuf[4228] = 256'h27017201b801e5010e0234023b02410252026c028c02c302070347038003a603;
    decBuf[4229] = 256'hba039b035d03e2026402b2010b017400c3ff7cff3bff00ffeffedefeedfee0fe;
    decBuf[4230] = 256'hecfe0dff17ff32ff19fff4fed2fea6fea0fec4fe09ff8bff09009b00fd005601;
    decBuf[4231] = 256'ha801d401fc01200241028702b502ef0214033703490365037f03a903db032704;
    decBuf[4232] = 256'h6d04ad04d604de04d704d004c004c504d304d704f2040a05270551058405c205;
    decBuf[4233] = 256'hfb054e069b06f5064a0781079f07a8078f075b071d07c20685063806f205e905;
    decBuf[4234] = 256'h02064606aa0622079407fb0759086508700852082408eb07c507b1079e078d07;
    decBuf[4235] = 256'h73075c0747074307550777079707ad0791075d07ec06190650056504c703fd02;
    decBuf[4236] = 256'h4702a001090180000200b1ff67ff3fff33ff3eff34ff2bff23ffeefebefe6dfe;
    decBuf[4237] = 256'h0afe92fd20fd9bfc42fcf0fbc4fbd2fb0efc87fc19fdcafd41feadfee8fefafe;
    decBuf[4238] = 256'hc9fe62fecffd1efd19fc25fb86fabdf96ff928f93df951f986f997f988f960f9;
    decBuf[4239] = 256'hf3f86ef8f1f77ff735f70df719f73af76cf79af7e4f73ef893f8f6f86ef9c0f9;
    decBuf[4240] = 256'h09fa4cfa71fa66fa34faf4f9cbf9c3f9d8f903fa4dfa7ffa9afa81fa4dfa01fa;
    decBuf[4241] = 256'hbbf97bf973f989f9e3f968fa09fba0fb03fc38fc48fc1cfcbffb82fb35fb17fb;
    decBuf[4242] = 256'h20fb49fb8dfbf1fb84fc0efd8bfdfdfd29fe51fe75fe96fef0fe45ffbeff3000;
    decBuf[4243] = 256'h9700da00fe000901eb0099002000afff47ff04fff8fe2fff75ffdaff5200c400;
    decBuf[4244] = 256'h0e0150014401f7009d0018009bff29fffdfed5fee1fe18ff5effb0fffdff1b00;
    decBuf[4245] = 256'h0000b5ff47ffa5fe0efe84fde3fc77fc3cfc2bfc3bfc67fcaafce7fc1efd3cfd;
    decBuf[4246] = 256'h45fd5dfd47fd25fdecfc9afc63fc45fc60fcaafc40fdd8fd61fe02ff43ff7eff;
    decBuf[4247] = 256'h90ff5fff15ffd2fe96fe75fe6bfe74fe8dfe85fe7efe5ffe59fe54fe62fe88fe;
    decBuf[4248] = 256'ha2feb0feb4feb0fe91fe62fe1dfecbfd68fd0afdb6fc7ffc89fca4fcfffc6cfd;
    decBuf[4249] = 256'hf1fd91fefefe60ffb9ffc9ffbbff92ff56ff35ff3fff48ff82ffa7ffbcff90ff;
    decBuf[4250] = 256'h3cffcffe4afecdfd5bfd11fd04fddffcd4fccafcc1fc98fc55fcf0fb78fb06fb;
    decBuf[4251] = 256'hbcfa79fa9efaebfa6dfb0efca5fc2efd64fd95fd69fd40fd1cfd11fd43fda7fd;
    decBuf[4252] = 256'h20fe92fedbfe1eff2aff1fff01ffd4feaafe85fe55fe29fe02fefdfd1dfe5dfe;
    decBuf[4253] = 256'hd3fe45ffacffefff14000900ebffabff71ff2dff12ff0aff20ff6cffc6ff4b00;
    decBuf[4254] = 256'ha500d500e400bc004f00e8ff8aff4dff42ff60ffa0ffdaff0000f9ffcdff79ff;
    decBuf[4255] = 256'h0bffc2fe7ffe5afe7bfeadfedbfef4feecfeaefe64fe0afee6fd07fe61fee6fe;
    decBuf[4256] = 256'h87ff1e008100b600a6005c00c9ff18ff72fedbfd79fd1ffd0ffd1efd61fd9dfd;
    decBuf[4257] = 256'hd4fd1afe36fe3efe27fef7fdb3fd60fd13fdf5fc11fd5bfdddfd7efeeafe4cff;
    decBuf[4258] = 256'h5eff4eff04ffc1fe9dfe66fe70fe8bfec5fe17ff64ff96ffb2ff99ff56ff03ff;
    decBuf[4259] = 256'ha0fe5efe39fe2efe38fe66fe7ffe86fe8dfe55fe11febffd88fd7efd99fde4fd;
    decBuf[4260] = 256'h3efeabfef5fe02ff0effedfecffed8fe12ff73ff2100f700c001ab0289031904;
    decBuf[4261] = 256'hcf044605b20514066e06e00647076f07ac07cd07d70729088c0804099609200a;
    decBuf[4262] = 256'h790aeb0a350b420b360b2b0b0d0b040bfb0a120b420b6e0b8a0ba40b9f0b700b;
    decBuf[4263] = 256'h380bf40ab50a9c0a940aa90ac80ae40ae90af70af30af70a010b110b2b0b5f0b;
    decBuf[4264] = 256'hb20b150c730ce00c290d520d450d0e0ddc0caf0c650c1f0ca80b160b8c0ac809;
    decBuf[4265] = 256'h11099a082e08f3070508f5070308db07b7075407c10610063a057104ba031403;
    decBuf[4266] = 256'h5102cf01290191002f00d6ffa5ffb4fff7ff4b00ae00f1001601f500af004a00;
    decBuf[4267] = 256'hb7ff2effd4fea4feb2fef5fe62ffe7ff6400b600e200d400b00063000900b4ff;
    decBuf[4268] = 256'h67ff21ffcffe6cfef4fd82fdfdfc5cfcf0fb8efb35fbe3fa9afa57fa02fa9ff9;
    decBuf[4269] = 256'h41f9ecf8b5f897f8c5f8fff851f988f9a6f979f91ef999f81bf8ebf7dcf704f8;
    decBuf[4270] = 256'h59f8d2f864f9eef947fab9fa02fb2bfb4ffb86fbccfb30fc8efcfbfc45fd52fd;
    decBuf[4271] = 256'h5efd3dfd47fd50fd8afdcefd20fe83fefbfe8dff1700b80024018601bc018b01;
    decBuf[4272] = 256'h4101c900360086ffe0fe48febffdd1fd22fee2fecdffe900a901120232021502;
    decBuf[4273] = 256'h9201ec00800045007b00cc008c0142021803a803f6033e04280414040204f203;
    decBuf[4274] = 256'he303f103e503f003fa030304fb03e403c203a20370032403ca025d02d8015b01;
    decBuf[4275] = 256'h0a01c000b300d70024019201f9017202c302d202c402a0023d02fa01be01c901;
    decBuf[4276] = 256'h0f027302d10225035c037a035f0336031003e002da02e002da02cd029e024002;
    decBuf[4277] = 256'had012401ca009900c6002301a901260257024802ea0134017d00a8ffdefe5cfe;
    decBuf[4278] = 256'h15fefffd61fedefeb1ff7b00fd00450104017a00d9ff42ffb9fe83fe73fe82fe;
    decBuf[4279] = 256'hdffe34ffadff1f0069005b00d6ffedfed1fd77fc90fb65fb8cfb3afc18fd54fe;
    decBuf[4280] = 256'h26ff9aff77ffd9fe9cfd21fcbcfa78f94df90dfa47fb17fdc7fe50004f012001;
    decBuf[4281] = 256'ha2002f003bff9dfe46fef8fde0fdcbfd90fd36fdc5fc40fce6fbd6fb5bfc43fd;
    decBuf[4282] = 256'h60feb9ffa100cb0058001eff4ffd9ffb16fa7df9abf92afa83fb24fdadfeacff;
    decBuf[4283] = 256'hdbff5cff50fe16fd9bfb9cfab4f98af9fdf9abfa88fb8bfc3afd98fd7cfdc5fc;
    decBuf[4284] = 256'hc0fb40fadbf83af721f688f55af584f544f6f2f6cff799f84ff997f981f946f9;
    decBuf[4285] = 256'ha5f80ef8acf79af70cf8aef89cf979fa09fb23fb0bfbcafa68fa33fa43fa6ffa;
    decBuf[4286] = 256'h97faecfa23fb55fb5efb46fbf3fa64fa8cf9c3f80cf8c5f7daf73df8ddf875f9;
    decBuf[4287] = 256'h4dfadcfa93fb3afca6fce1fccffc9efc54fc2cfc38fc6ffcb5fc07fd6afde3fd;
    decBuf[4288] = 256'h75fe4dff16000101600143018c0058ffddfd78fc90fb11fbebfa54fbf2fb2efd;
    decBuf[4289] = 256'ha9fe0e00af0158022502e00011ff61fd67fb13fad6f97efae3fb9bfe1a026505;
    decBuf[4290] = 256'h88077a09d409de083d060e0310001efe0ffd06fe7bff670220054e0897093309;
    decBuf[4291] = 256'h24084005c00175fe52fceefbfefc3eff740297045007aa07fd07870633050703;
    decBuf[4292] = 256'h91013d00000038009d013e03c7042c065a063006bd05c904ec032203a0022902;
    decBuf[4293] = 256'h920130011e016f011102d4028b030104ec031403d801080058fecffc36fc08fc;
    decBuf[4294] = 256'h86fc93fdcdfef4ffb30091007100a8ff59ff42ff82ff0c001e00ccffeffe15fd;
    decBuf[4295] = 256'hc1fb8cfa54faedfa32fc55fe60003c02f6022e03c9016eff8afc0af9b0f668f5;
    decBuf[4296] = 256'hcbf590f7d0f906fd04002f018901930087feabfc80fa9ff95bf990fa19fc4afe;
    decBuf[4297] = 256'h5500a9016202ba01bb001aff91fd92fc07fc31fc57fc06fde3fdacfe63ff0900;
    decBuf[4298] = 256'h4a005e00e1ff0dff0bfe17fdfafb87fb1efb7dfb46fccefd57ff2201d2027b03;
    decBuf[4299] = 256'h48030302340083fe6bfd38fd20feefff1b02bc043507d0081b09d708a2071906;
    decBuf[4300] = 256'he803dd011101d300ec011d04be0682081e0a680a9c09ec07f3059f046a03c202;
    decBuf[4301] = 256'h2902fa0125024b02f9029703d4044f061a08ca09e30a160b8b0a0f097806ff03;
    decBuf[4302] = 256'h1b01f0ff96ff8c009802fc043b07b1087d093f0997083207d7049702f7ff32fe;
    decBuf[4303] = 256'h3bfd86fddafe8a00840260049405cc053305ef037402a900f8fe70fd3dfd24fe;
    decBuf[4304] = 256'ha0ff6b0196030c05d8059a058204b70206017eff19fe8dfd0cfeccfe4b00b001;
    decBuf[4305] = 256'hf502cb02be01b3ffa8fdccfb8efbc6fb2bfd29ff7d00b201ea0151010d00e6fe;
    decBuf[4306] = 256'h8cfda4fc26fce6fc66fe9700a2027e0437058f0490034b022401b1001a01f701;
    decBuf[4307] = 256'hc002da029302a501490005ff8afd8bfc00fcd5fb95fccffd9fff4f01d802d703;
    decBuf[4308] = 256'ha803810242005efda5fa2cf835f780f7e4f9c8fc47009203b505190609056e03;
    decBuf[4309] = 256'hcd0054feb9fcd8fb1cfc51fdbbff9f0257051c076e078e062a04a10056fd33fb;
    decBuf[4310] = 256'hcffadffbc3fe43028d05b107db0817073304b30068fd45fba8fb6dfdf6003105;
    decBuf[4311] = 256'h2d09bb0a330b100957067402ddff83fd16fd40fe0500450250042c0661072807;
    decBuf[4312] = 256'h290688048f02b30003ff5afec1fd4cfecbfed7ffcc006a01c0010e02b5027703;
    decBuf[4313] = 256'h2e04d404bf04e703ab022f01caff3fffc1fe34ff9dfffcff8b004201e8018002;
    decBuf[4314] = 256'h0903d40221021c01e2ffbbfe48fe25fe44fe61fe7bfe93fefffeb0ffe5000b02;
    decBuf[4315] = 256'h1803f5025702e1007cff38fe65fd8bfdaefd0dfe9dfe54fffaffe800c5015502;
    decBuf[4316] = 256'hd8021f030903a7020602ed00e1ffa7fed4fdaefdd1fdaefe77ff2e007500b600;
    decBuf[4317] = 256'hf10027017801a4017c013f01dc009a00a600c700a9002000f9fe2afdf5fbddfa;
    decBuf[4318] = 256'haafa35fb07fc61fda5feccffbf019b03c705120646051a034effaffb55f90cf8;
    decBuf[4319] = 256'h37f9b0fbf0fdfbff5f02fb037005c40602075a06290488010eff73fd28fd6cfd;
    decBuf[4320] = 256'ha1febaffb900a101cb01a4013c011f00c6fe24fd9cfb03fb8efb09fd3aff4501;
    decBuf[4321] = 256'h99025203aa02450147ff6bfd36fc1dfbeafa19fbebfbf8fcecfd8afe6efe1ffe;
    decBuf[4322] = 256'h79fde2fc7ffc6efcdffcbdfdd9fee6ffda00ba00f1ff69fe00fc65fa84f9c8f9;
    decBuf[4323] = 256'hfdfa66fda6ff1c017002ae02e6024d02c201ef00e2ffa9fed6fdb0fd5efebaff;
    decBuf[4324] = 256'hfe002502ff010b0170ff57febefdecfdbffe18005d013002a3025103ef034604;
    decBuf[4325] = 256'hf703f2022d0101fff6fcb2fce6fdc0003f047b08540bd80b600b6108a905c501;
    decBuf[4326] = 256'h3800cffe61fe8cff5001eb026104b505ea06b206b305b503c90010fe4cfc55fb;
    decBuf[4327] = 256'ha0fb6cfc1cfea5ff3e000f0091ff84fe4afd24fc17fb23fa85f9a1f98dfae8fb;
    decBuf[4328] = 256'h8afda2fe3bff0dff3afe7bfdccfcadfc90fc41fc2afc14fc4ffc14fdfffd9dfe;
    decBuf[4329] = 256'h2dff12ffcbfee1fe43ff2b0009015f01a80044ff79fd44fc9cfbcffbb7fcddfd;
    decBuf[4330] = 256'h9dfec0fea1fe84fe6afeb1fe1dff7ffffcff4e009700a5006800d9ffdafea0fd;
    decBuf[4331] = 256'h79fcb9fb0bfbebfa42fb2dfcc8fdc1ff2502c003a004d4032d01fffd00fb9dfa;
    decBuf[4332] = 256'hacfb90fe49010d03bb024501e1fe46fd66fcaafc6cfc34fc9bfbc9fb9cfcdcfe;
    decBuf[4333] = 256'hc0017804880536052a033e0086fd0cfb71f926f9f2f9a3fb0cfef000a903b804;
    decBuf[4334] = 256'h66045b026fffb6fca7fbf9fb6ffd5b004c0211040805bd04e1023101c7fe2cfd;
    decBuf[4335] = 256'hb6fb82fc32fe0c01c5033e063507ea069605e603cd029a022503f803b8042005;
    decBuf[4336] = 256'h0105ab04f4037d031103d602c402f5022103640388033b03a5026101c0ff37fe;
    decBuf[4337] = 256'h38fd66fd39fe92ff3301bc02ef026402950069fec8fb04fa56faccfbb8fe3702;
    decBuf[4338] = 256'h8205a50709088f050702bcfe99fc6efb33fd72ffa902f10355049002500045fe;
    decBuf[4339] = 256'h69fc34fb8cfa8df95ff9ddf936fbeefd6d01c703eb05c0044702befe73fb2bfa;
    decBuf[4340] = 256'h8efa53fc93fe9e00f201ab02e3024a021c029e01c401e701850215036303ec02;
    decBuf[4341] = 256'ha80107000dfeb9fc00fcc8fbfbfb29fcabfbebfaf7f959f93cf9f3f957fb88fd;
    decBuf[4342] = 256'h2900ee01e4022f03db01afffa4fd40fb49fafff953fb87fc10fedbff1001b801;
    decBuf[4343] = 256'h510280025602960116004bfe1ffc14fa38f803f73bf73af895fa7afdf9005303;
    decBuf[4344] = 256'h9b04380428038d01ecfe73fc33fabdf8f1f7abf8a4fa18fe620161045206ad06;
    decBuf[4345] = 256'h5b06e5040903590160ff84fdd3fb9bfb34fc1cfdeffdc8fdd4fcf7fbdafbf9fc;
    decBuf[4346] = 256'h39ff1d020f046904ce0298ffbefb28f9bff72cf857f9d0fbb4fea6001f031604;
    decBuf[4347] = 256'h610495036901c8fe04fd69fbf3f9aff9edf925fa58fa40fb67fc0dfe25ff58ff;
    decBuf[4348] = 256'h70fea1fc75fa00f9acf7f2f62af729f86ef9e9fae8fb73fc49fcd6fb28fb87fb;
    decBuf[4349] = 256'h89fc4ffe7a005b011701e2ff79fd39fbc3f97ff938fac1fbf2fdfdffd9019302;
    decBuf[4350] = 256'hcb02cc012a00a2fea3fd74fd9efd5efec7fee6fe57fea0fd6bfc44fbebf903f9;
    decBuf[4351] = 256'h30f8a3f8ddf955fccffe0e01ef01ab017600edfe54fe26fe50fe29fef0fc74fb;
    decBuf[4352] = 256'ha9f96cf914fadffb0bfe81ff4d008a005200eb001a0198012501310096fe9cfc;
    decBuf[4353] = 256'h48fb14fadcf975fab9fb89fd3000a9028e05b8065e066705c6024d000dfe97fc;
    decBuf[4354] = 256'hcbfb84fc0dfe0a010904c10686087c099c0848071c05a703630325035d03f603;
    decBuf[4355] = 256'hc8034903d602b302510354048e05b5067507980778075b07aa072008b8084109;
    decBuf[4356] = 256'h2f097d081807e7047203a602e3026c040307320a300d5b0eb50e1a0d790a4b07;
    decBuf[4357] = 256'h270536032602d401b4028003be03f603c303f1037004300524068306f305d404;
    decBuf[4358] = 256'h2d0315027c0107028502f8021b03fc02520371046406c808630a190ac508a205;
    decBuf[4359] = 256'ha302790169006001d602a203d7047f05e40685087f0ad30b950b9c09b0063003;
    decBuf[4360] = 256'he6ffc2fd5ffdb9fd54ffca00a6025604df05de06c607f007ca0790061505e402;
    decBuf[4361] = 256'h43007ffe2cfe0dff7101f90444088c096208e805600215fff2fc8efc53fe3701;
    decBuf[4362] = 256'h7d055608ed0a650b1c0a9d06520379ffe2fc6afcd7fc3bfd95fd8cfed7fe2b00;
    decBuf[4363] = 256'h57028d058b087d0a8c0b960af507c604ed004dfde4fb52fc43febd00a1035a06;
    decBuf[4364] = 256'h690760088007a40578036d0109ff12fec7fd1bffcb00540253038203af02a201;
    decBuf[4365] = 256'h7f015d020c042f077708db086106340238fea1fb29fb4cfd0500330357050f08;
    decBuf[4366] = 256'hd409140c1f0e630eb30c69095b024bfbb6f636f47cf6edf94ffe6f03e106020a;
    decBuf[4367] = 256'h940a0609ac06d3022afe09fb54f9e1fa3bfd1501ab0305064e07ea0626058a03;
    decBuf[4368] = 256'h7f01a3fff3fd2bfe90ffeb01cf04c106d0077e070806b4047f0367026801c6ff;
    decBuf[4369] = 256'haefe15fea0fe6f009b021104550420039701320004002b011e037204af040704;
    decBuf[4370] = 256'ha2025d018b00b1005f013d0240037904f8046b057704dc02720033fe92fb82fa;
    decBuf[4371] = 256'hd5fae0fcccff4b03a505c9072c081d07940359ff5cfbc6f86cf6d9f6cbf8f9fb;
    decBuf[4372] = 256'hd3ff7203bd060608a20729054402c5fe6bfc22fbbffa19fbb5fc95fdd9fd17fe;
    decBuf[4373] = 256'hdffd12fe9dfe1bff8effb1ffd4fed1fd97fc19fc8cfcc6fd41ff0c01c501fd01;
    decBuf[4374] = 256'h640120004dffdafe2bfe0cfe7cfd2efde6fc7efda4fe1f00ea011f03e702e801;
    decBuf[4375] = 256'h47004dfe71fc34fcdcfca7fed30049021503e00176ff37fd96fa86f9d9f9b9fa;
    decBuf[4376] = 256'h0dfcbdfd46ffab0036010c0166ffddfd78fc03fd7efe1501da022c03b601cafe;
    decBuf[4377] = 256'h4bfbe2f974f966fb2afd21fe6cfea0fde6fcaefc47fd2ffe02ffc2ffe5ff46ff;
    decBuf[4378] = 256'h44fe0afd37fcc4fbb8fc53fe4c0018015f0086fd06faacf764f655f884fb82fe;
    decBuf[4379] = 256'h3b014a02530173001fff66febefdf1fd1ffe49fe09ff72ffd3fe24fd01fa03f7;
    decBuf[4380] = 256'h11f521f605f913fee5024707fc088109270728041bff48faa6f460f2b0f190f3;
    decBuf[4381] = 256'hb0f8e4fe0e03d806280607030bff62fa41f7aff634f77efa58feee0057020f01;
    decBuf[4382] = 256'h56fe73fadcf755f89df956fc65fd5cfe7cfd28fc6efba7fbdafbabfb2dfb06fb;
    decBuf[4383] = 256'h6ffbcbfc26ff6601db020f02e4ff18fc78f81ef68cf6b6f730fa70fc7bfebffe;
    decBuf[4384] = 256'h8afd91fbb5f9fcf834f9cdf9b5fadffa1ffa71f912f92ff9e5f92dfac1f9e9f8;
    decBuf[4385] = 256'he6f7c3f7e0f8d3faaffc68fd4ffc84faddf718f622f56cf5c0f6f5f70ef90dfa;
    decBuf[4386] = 256'h98fa1afa73f87af616f420f36af3bef46ff6f7f72af843f7c7f562f4d7f356f4;
    decBuf[4387] = 256'h62f5e2f647f88cf9b2fa3ffa05f98ef65ff361f036ef91ef2cf137f313f548f6;
    decBuf[4388] = 256'h60f7c5f867faf0fb57fb59f95df560f1c1ed48ed47f0c6f302f8fefb83fcfbfc;
    decBuf[4389] = 256'hd7faadf99df84bf800f834f7f7f6def5dff49af3c8f2a1f296f370f5d4f714fa;
    decBuf[4390] = 256'h89fbcdfb0bfc43fc10fce2fb64fbbdf954f714f509f3b5f1f3f19bf29af3dff4;
    decBuf[4391] = 256'h06f612f792f8f7f9dffa09fbe3faeef9d2f85ff8c7f8e4f98afb13fdacfd7efd;
    decBuf[4392] = 256'h02fc6bf9f2f6b2f467f433f5e4f66df86cf9e0f811f76af4a5f253f25ef45af8;
    decBuf[4393] = 256'h7afdec000d049f041103b800b9fd3afae0f7bcf592f4ecf487f6bef9bcfcaefe;
    decBuf[4394] = 256'h08ff11fe06fcb2fa6bfb65fd510042029d02010161fe7dfae7f78df51ff5bcf4;
    decBuf[4395] = 256'h80f6c0f88cfc340155042e07aa0650049bff3afb84f900f969fab1fbdcfcccfb;
    decBuf[4396] = 256'h31fabbf8fff82bfb61fe3b02d1045904110391ff46fc48f91df878f8caf8aaf9;
    decBuf[4397] = 256'h76fab4fa5dfb5cfc5afe3600e6011e021f01c4fee0fb27f9aef600f7e0f744fa;
    decBuf[4398] = 256'h84fc25ffe900e001c002f401c9ffbdfde1fbadfa55fb86fd91ff5d00200026fe;
    decBuf[4399] = 256'h4afc16fb4efbe7fbcffcf9fc86fc1dfc7cfc2bfe4e0171036305080512043103;
    decBuf[4400] = 256'h7503aa04c305f605b10439020bff0cfca9fb03fc43fee400a8029f037f04c304;
    decBuf[4401] = 256'h86044d041a048f031103eb020d03ee02980278011f0037ff61ffba0015035505;
    decBuf[4402] = 256'h6007b408f208ba08bb07760653044702e3ff48fe28ff8c01ba059208290bb10a;
    decBuf[4403] = 256'h6809e9058f036b010801cc02670473064f088c08c5082c08440771064b06b306;
    decBuf[4404] = 256'hd306b606ff052a05270478035903e90308056106a6072109200a080b320b720a;
    decBuf[4405] = 256'hf308c2064c058004390532079609310b120cce0b1d0a2408d0061706bf062408;
    decBuf[4406] = 256'hc609de0aab0a200af9083a088b076c07c2077908ad09290bf40c1f0f2b117f12;
    decBuf[4407] = 256'hbc1284128511e40f0a0d8b095f04ed008bfcf9fb90fead04820ad00f4213e213;
    decBuf[4408] = 256'h2d12970f1e0f8c0fef0fff100810fd0d990bfd09b309070bb70c5f0dc60cc80a;
    decBuf[4409] = 256'h6408c90614077809000d4b106f1299133f134812fd11b911f7112f1296115110;
    decBuf[4410] = 256'h820ed20c290c280d6d0e400f660f2c0e5d0c310ae6093a0be10dc5116415be17;
    decBuf[4411] = 256'h51175f153112320f7a0c6a0b180bf80b4c0d810e0a10a310d110a7108110a410;
    decBuf[4412] = 256'h421145127e13fd13d6139d122111221051107811841261128710130dd8082207;
    decBuf[4413] = 256'hb008eb0c2f13af1ab61da01e201c56182312f80d2e0a7e091e0ab00a340bad0b;
    decBuf[4414] = 256'h1a0c7e0cd80c730ee90fc5117e122713c013ee1318148b146814ca131b12740f;
    decBuf[4415] = 256'hfa0cbb0aaf08f308280a910c760f2e12891292115c0e820ae3066a068e08d40c;
    decBuf[4416] = 256'hf411661506165114b110580e340c0a0baf0a14099e07c20584050d07a4091e0c;
    decBuf[4417] = 256'hb90dd90c750a90076606c0060009a10b650d130d9d0b390955069d032301d100;
    decBuf[4418] = 256'hb1019d04e408e00c6d0ee60ee70b68080e06c5042905ed064007f506a105f103;
    decBuf[4419] = 256'h6802cf015a022d03ec032605a1060608ee08c4081e072505c102ca011502e102;
    decBuf[4420] = 256'h9a0362036302650011ffd3fe5c00f3022206450870091509d50635040601e3fe;
    decBuf[4421] = 256'hf1fc01fe9cff3d020104f804ed02010048fd39fc2ffdfb009b04e5072e090308;
    decBuf[4422] = 256'hd504d6011eff59fd07fd52fd96fdd3fd0cfea5fe8cff5f006c01a602cc034004;
    decBuf[4423] = 256'h9103b70153ff13fd08fbc4faf9fb81fde6fe72ff9ffeacfcd0fa9bf9d3f96cfa;
    decBuf[4424] = 256'h0efc97fdfcfee4ff6200d5003e011e01c800ddffc0feb3fd05fd67fcd7fb20fb;
    decBuf[4425] = 256'h4bfabbf9a1f976faecfbb7fd70fe38fed3fc1cfa9cf642f4faf296f2a6f3e6f5;
    decBuf[4426] = 256'h1cf91afc0cfe66fecbfc2afafcf6d8f4aef3bdf4fdf69ef9adfa5bfae5f8f9f5;
    decBuf[4427] = 256'h08f443f296f20bf46ff6aff8bafa86fb49fbdff8fbf542f37ef187f067f1bbf2;
    decBuf[4428] = 256'hf0f399f400f4bbf294f16ef162f2fdf3f6f5c2f684f6fbf4caf2bff05bee64ed;
    decBuf[4429] = 256'h1aede6ed96effff188f5d3f8f6fa21fcc6fbe2f89bf49ff000eda6ea13eb05ed;
    decBuf[4430] = 256'hc9ee09f1e9f1b5f2f3f24bf218f2d3f0acef53eec8ed46ee9fef9ef17af3aef4;
    decBuf[4431] = 256'he6f4e7f346f2ddef41eeccec88ecbced26f00af3c3f5d2f680f6dff3fcef5cec;
    decBuf[4432] = 256'h11e9eee651e761e8fce972eb4eedfeeef7f0d3f2fff44af57ef4cef284ef39ec;
    decBuf[4433] = 256'h3be949e785e5d7e5b7e61be9a4eceeef12f275f21bf280f00aefc6ee7fef08f1;
    decBuf[4434] = 256'hd3f28cf3e4f24df01eed45e9a5e53ce4aae49be6cae9a3ed3af0a3f15af0a2ed;
    decBuf[4435] = 256'h28ebe9e808e85ce90deb96ec95ed20eef6ed69ee17eff4ef6af1cff2b7f335f4;
    decBuf[4436] = 256'h0ff461f3c6f15cef78ec86eac2e870e8e5e9c1eb69eee2f07df25ef3b2f4eff4;
    decBuf[4437] = 256'h47f47cf2d5efa6eca8e944e954ea38edb8f002f426f689f67af5def3d3f107f1;
    decBuf[4438] = 256'hc0f1d9f2a4f4d9f581f64ef60af5e6f2dbf0ffeec1ee69ef9af1d1f4cff788fa;
    decBuf[4439] = 256'h97fb45fbcff96bf72bf520f3ccf113f1dbf074f1fff1d1f291f340f4def434f5;
    decBuf[4440] = 256'h4ef566f5d2f583f688f736f856f8c6f773f674f498f2dff1a7f10cf30af56ef7;
    decBuf[4441] = 256'h09f954f988f85cf6bcf38df06aee3fede5ec92ecddeca9edd5ef76f2a4f5a3f8;
    decBuf[4442] = 256'h22fc8bfd1efd2cfbfef724f48ef143eefbec5eed23efabf2e7f6c0f956fcdefb;
    decBuf[4443] = 256'hbaf93bf6fff127ef99ed21ed69ee5bf06af1bcf107f2c3f185f1bef157f29bf3;
    decBuf[4444] = 256'h16f515f644f6c5f5b9f4c5f3e7f2caf281f3e6f4b1f661f809f9a2f917f9f0f7;
    decBuf[4445] = 256'he4f6aaf583f4c3f35af33bf357f372f3e8f3d6f4f3f5fff6aef70df829f80ff8;
    decBuf[4446] = 256'hc8f75cf7abf677f5fbf3caf155f089ef4befd4f09ff2cbf4d6f62af8e3f88bf9;
    decBuf[4447] = 256'h24fa53fa7dfa57fa34fa14fabef96ff99af824f7f3f452f243f1f0f0d1f1bdf4;
    decBuf[4448] = 256'h75f7a4faecfb50fc40fb49fad4f808f845f8eef8b9fae5fcf0fe440079012102;
    decBuf[4449] = 256'h8801fd00d6ffc9fe4afd4bfc06fb88fa61fa3efa5efa7bfa95fa3bfb80fcdafe;
    decBuf[4450] = 256'h1a01bb037f05d205f1049d03ed01d500d6ffeefe6ffe49fe3dff170113051009;
    decBuf[4451] = 256'hb80d990f4e11c10f850b8907ea039f0031009500c303c2067a09f40b460c660b;
    decBuf[4452] = 256'h9a0a5c0a940a930b7b0ca50c990b8e09ed067304d80223037704a3064309720c;
    decBuf[4453] = 256'h950e871096114411ce0ff20d420c490a7d093f09c80af90c9a0f5e11fa124413;
    decBuf[4454] = 256'h68113d0f9c0cd70ae1092b0a070c330ea90fed0faf0f260ec10cd90b030c770c;
    decBuf[4455] = 256'h250d020e920e490f1f1021111612b412d0124e1219119e0f390e510d7e0c580c;
    decBuf[4456] = 256'hc10c5f0d620e100ff00e9a0e7b0d6e0cc00b1f0c210da10ea00f2b10ad0fed0e;
    decBuf[4457] = 256'hf90d9a0db70dd10de80dd30d490d5b0dcd0daa0e45105e1191110611df0fd20e;
    decBuf[4458] = 256'h6a0e080fd10fbc101b118b10a00f020f720ec10e380f220f230e5d0c320a9107;
    decBuf[4459] = 256'h81062f060f07eb08930b0c0e4c10c21106124c11530f770d430c9a0b330cd50d;
    decBuf[4460] = 256'h5d0fc210f1101e10120f1d0efe0dc70ee60fa6108310e50fe30e340ed50db90d;
    decBuf[4461] = 256'h6a0d940c580bdd0944091609910af60b970db00e490f1a0f450f6b0fd40fb40f;
    decBuf[4462] = 256'h5e0f3e0e320d3e0cdf0ba80cc70dd40e820f630f260eab0ce00a30098808bb08;
    decBuf[4463] = 256'ha309c90a230c670de30ee20f6d104310cf0f960ec60c9a0a2509e1081e09a70a;
    decBuf[4464] = 256'h720c230e5b0ec20dc40be80937086f086e096d0b490df90ea10f6e0f400f160f;
    decBuf[4465] = 256'h3c0fd30ef60d470c24092606fb045605f10692090b0ca60df10d9d0ced0af408;
    decBuf[4466] = 256'h2808ea0792089109790a4c0b580c920db90ec60f2e100f10460f5a0e7d0d600d;
    decBuf[4467] = 256'he30db90e820f391021105e0f0b0e0d0c310a0508250769079d08070beb0ddd0f;
    decBuf[4468] = 256'hec109a10ba0fde0da90c000c670bdc0a060b2d0b950bb20c720d200e010efe0c;
    decBuf[4469] = 256'h7e0bb309fa083209fd0a290dca0f43123a13ef129b116f0fcf0c550aba086f08;
    decBuf[4470] = 256'h2b086908a1083a09c509440ab70ada0a7b0aeb0997089906bd048803c103f205;
    decBuf[4471] = 256'hbd095d0d98114d13c011660f680caf09a0084d080308bf078a069104b5027702;
    decBuf[4472] = 256'h90038d06660afd0c750d070d4f0a6b06d5037b010e013802b20496074e0ac80c;
    decBuf[4473] = 256'hbf0d090eb50c8a0a7e08a206e905910690071c08f1073207f80525054b05fa05;
    decBuf[4474] = 256'h1607d6073f085f084208c4089a092a0a100adb08b70617049d01a600f100cd02;
    decBuf[4475] = 256'h7405a308c60af10b960b440b39095d073105bb03df01a201da01a5035505be07;
    decBuf[4476] = 256'hfe09de0aaa0bf10a490ae4089f0778061f057e036502cc019e01c4026b04f305;
    decBuf[4477] = 256'h8c065e06e304b202a700dbff21ffcaff2f01d002e9038204530481037402c601;
    decBuf[4478] = 256'h6701bd01dd0236047b054d06c0069d06c00511046a013bfe3dfb4bf9f1f8e7f9;
    decBuf[4479] = 256'h1efd1c00d502990447043c0250ff97fc1efa82f8a2f76ef827f940fad9fa64fb;
    decBuf[4480] = 256'h8efbb5fb63fc80fd26ffaf00ae01dc015e010400c0fe44fddffb3efa25f926f8;
    decBuf[4481] = 256'h55f827f981fa22fcabfddefd53fd2cfc39fa5df8adf605f638f6d9f742facbfd;
    decBuf[4482] = 256'h25006d010a0190feacfbbbf9f6f748f829f97dfa36fbdefb11fc40fcbefc31fd;
    decBuf[4483] = 256'h54fd34fd6bfc80fba3fa13fac5f94ef9b6f854f866f8f8f8d0f99afa7ffaaaf9;
    decBuf[4484] = 256'h34f8cff6e7f565f6bff7bdf921fcbcfd32ff76ff41feb8fc21faf3f6cff4a5f3;
    decBuf[4485] = 256'h4af3e6f4f1f655f94cfa96facaf996f87df74af71cf7f1f67ef68af56ef414f3;
    decBuf[4486] = 256'h2cf25af133f156f1f4f1bef211f456f57df689f738f818f888f79df681f527f4;
    decBuf[4487] = 256'h3ff36df246f2f5f211f404f6e0f715f9ddf8def73cf6d3f338f258f124f258f3;
    decBuf[4488] = 256'h71f4d6f504f632f58cf303f238f07eef27f08cf18af366f59bf643f7aaf665f5;
    decBuf[4489] = 256'h3ff4e5f25af284f244f338f455f561f69bf71af88df8b0f890f8c7f7a7f601f5;
    decBuf[4490] = 256'h08f32cf17cefd4eed3ef2df212f5caf78ff9e1f901f925f7f9f483f32ff276f1;
    decBuf[4491] = 256'h3ef1a5f076f04cf0bff0f9f174f3a5f546f80bfaa6fb5bfb7ff95cf65ef3deef;
    decBuf[4492] = 256'h75ee08ee32ef42f094f0dff023f1e5f0adf0e0f00ef18df100f268f288f2a5f2;
    decBuf[4493] = 256'hbff2a7f292f2a5f270f21ef29af18df081ef8deeefedd2ed54eecbeee1eea6ee;
    decBuf[4494] = 256'h05ee6eed5aedd7ed8aee8fef83f021f1b1f134f27bf23af214f144ef94ed2beb;
    decBuf[4495] = 256'h34eae9e9b5ea66ec5feec3f05ef23ef382f34df2c5f0faee49ed81ed80ee7ff0;
    decBuf[4496] = 256'h5bf20bf4d3f36ef213f0d3ed5dec19ec4eedb7eff7f198f45cf6aff664f688f4;
    decBuf[4497] = 256'h5cf2e6f01af058f001f166f2f1f2c7f207f213f1f3f0bcf144f33df591f64af7;
    decBuf[4498] = 256'h12f779f691f56bf45ef3def179f091ef67ef27f0edf118f424f600f83df805f8;
    decBuf[4499] = 256'h6cf784f609f50af422f3a4f2caf2bef35af553f7a7f8e4f8ccf701f6d5f35ff2;
    decBuf[4500] = 256'h93f14df2f5f2f4f322f4a4f3e4f236f255f2e5f204f45ef5a2f6c9f789f8acf8;
    decBuf[4501] = 256'h8cf8c3f7d8f6bbf5fcf493f4b3f47cf567f6c6f6a9f6f2f5bdf497f3d7f2faf2;
    decBuf[4502] = 256'h98f39af4d4f5a7f667f78af7e9f7ccf7e6f72df843f856f845f8b2f7b3f679f5;
    decBuf[4503] = 256'hfef3fff217f241f24ef313f5c4f6dcf775f88df767f60df582f4acf4b9f57ef7;
    decBuf[4504] = 256'h2ef947fae0fab2fa88fac8f95ff9c1f885f70af6a5f460f3e2f2a1f367f517f7;
    decBuf[4505] = 256'h10f964faa2fafaf961f91cf8f5f69cf5b4f48af44af5c9f694f8c9f971fa3efa;
    decBuf[4506] = 256'h56f9d8f865f8cef82cf983f969f9c2f82bf8c9f722f8f5f8f8f9ecfa0cfbb6fa;
    decBuf[4507] = 256'h96f98af850f7d1f65ef681f61ff7e9f7d4f8f0f9fdfa37fc09fdc9fda6fdc9fc;
    decBuf[4508] = 256'hc6fb8cfa0efa34fae3fac0fb16fcc8fbf2fa63fa48fa4efb13fdc3fe6cff39ff;
    decBuf[4509] = 256'hf4fd25fc74faccf965fa4dfb74fc34fd11fd73fc70fb7cfa9ef948f962f968fa;
    decBuf[4510] = 256'he7fb18fe2300ff01b902f10258027001490089ff21ff7fff49006801c1020604;
    decBuf[4511] = 256'h840411041d03c1017d00aaff84ff7800d40175038e04c1049204c00300035102;
    decBuf[4512] = 256'hf301490200030504f904d6056606b506cc06e206a7062a0677050005c0049705;
    decBuf[4513] = 256'h470772097e0bd20c940c7b0b160ad208a8086709a10a740be70b7e0be00a8a0a;
    decBuf[4514] = 256'ha40a4a0b380c160d6c0d1e0d180cde0a0c0a4c09b509d10ade0b5d0dc20e4e0f;
    decBuf[4515] = 256'h20104710980fbb0e0c0de00ad5088107be07b7091b0c000ff1100112ae11f911;
    decBuf[4516] = 256'h2d11ef104710ae0f690e970d8a0c220c410c970c7d0c360cca0b8f0b0c0c000d;
    decBuf[4517] = 256'h800e4b107f11b711ea111912ef111512f2115411c4104210fa0f3b109d10d310;
    decBuf[4518] = 256'hc3103e109d0f310f930f58104311a2111211be0f1d0e040d9d0de20e06111113;
    decBuf[4519] = 256'h6514a314db14a81479144f14dc132e13501287116d117212f21357153f161516;
    decBuf[4520] = 256'h5515a614481464141b15f1150e16bf15ea14e71338131913a913c8148815f015;
    decBuf[4521] = 256'h1016ba1537159114fa1397133e130d13c412ec124113e613bb1485159f158715;
    decBuf[4522] = 256'hc4140d14f6130b1495147d151b16711657161016a415691510157d14cd132713;
    decBuf[4523] = 256'h6412e1119a112e11f310e11032111012ab133415991681170217f61576141113;
    decBuf[4524] = 256'h2912ff11721220137c146415df167817a7178016da14e11205114b10f410bf12;
    decBuf[4525] = 256'h6615df17d6188b18af168414e3111e1071105111b51350155b179f17e616ce15;
    decBuf[4526] = 256'h0314ce12b5111c1104122b13841426163e17711789160e1543138a12c2122714;
    decBuf[4527] = 256'h8216c218381af4193a1941176515b5139c1269123b1265122513d3137114c814;
    decBuf[4528] = 256'hae14371474138912ac11551107114e11111230133d147715a1157b154114c612;
    decBuf[4529] = 256'hfb104a0fa20e6f0e570f7e102412ad13ac14da140714151239100d0e2d0d710d;
    decBuf[4530] = 256'ha50e9e10f211ac12e412e511fd10820fb70d820cda0b410b6f0bed0b470de80e;
    decBuf[4531] = 256'h7110d6110412de109e0e710a98070a069205b6076e0ae80c830e380e6c0d400b;
    decBuf[4532] = 256'hcb097708bd071507e2065706810641077b084a0a7f0b270cf40bb00a34096907;
    decBuf[4533] = 256'hb905a104a2031603ec025f03df04aa065a0873090c0a8109ae080807ef058a04;
    decBuf[4534] = 256'ha303d0025d02f4015302e3029a03e10375034e022b0020fe54fd16fd2efef9ff;
    decBuf[4535] = 256'h25029b036704ae0395026400eefe12fdd5fc0dfd0cfeadff36019b0283035903;
    decBuf[4536] = 256'h4c02cc0001ff51fd39fca0fb71fb9bfbc2fbe5fbc5fb35fb7efa79f9cbf86cf8;
    decBuf[4537] = 256'h89f8a3f819f95af947f911f97ff8f5f79cf76bf7b5f77ef880f9bafa8dfb67fb;
    decBuf[4538] = 256'hfefaa2f901f878f679f5eef46cf579f6b3f785f8acf8fdf7a1f6a3f4c7f292f1;
    decBuf[4539] = 256'hcbf1caf26bf4f4f58df65ef68cf5e6f35df25ef1d3f0a9f0cff038f1d6f19ff2;
    decBuf[4540] = 256'h8af367f4bef4a4f45cf4c5f33cf306f3b5f26bf2f3f11ff11df06eef0fef2cef;
    decBuf[4541] = 256'hafef55f018f166f11ff187f0afefe6ee2feee8edd2ed35eed5ee42efa4efd9ef;
    decBuf[4542] = 256'ha9ef5fef01ef94ee2dee05eeb0ed63ed45ed05edcbeca6ec68ec3fec55ec77ec;
    decBuf[4543] = 256'hd5ec68eda3ed6eeddbecb5ebe6e9b1e898e7ffe68ae7b1e857ea50eca4ed5eee;
    decBuf[4544] = 256'h26ee27ed85ebfce9fde8cfe84de95aea4eeb2bec82ecd0ecb8ec4cec9cebc6ea;
    decBuf[4545] = 256'hc3e989e8b7e743e766e704e8cee8ede9adea16eb77ea02e937e70be595e3c9e2;
    decBuf[4546] = 256'h82e30be53ce748e924ebddeb15ec7ceb94eac1e902e90de86fe78ce743e8a7e9;
    decBuf[4547] = 256'h72eb22edcbed98ed53ecd8ea73e9e8e86ae890e8e2e7c5e6b8e5c4e4a5e46ee5;
    decBuf[4548] = 256'h59e636e7c6e7ace765e74fe78ae707e879e84de8b9e7e2e618e696e5dde5cbe6;
    decBuf[4549] = 256'he7e741e985ea04eb77eb9aebb9ebd6ebbceba4eb38eb39ea45e928e868e700e7;
    decBuf[4550] = 256'h1fe7afe766e80ce922e9c0e8fbe7dce61ce6f9e558e694e764e998ea41eb74eb;
    decBuf[4551] = 256'h8ceab9e946e998e839e856e870e887e81fe9a8e96dea58ebb7eb0decf3ebaceb;
    decBuf[4552] = 256'h96eb82eb4deb1cebd2ea75ea38ea6feac9ea67ebfeeb12ecdceb6aebabea28ea;
    decBuf[4553] = 256'h40eaacea84eb86ec35ed94edb0ed96ed7fedebed26ee7feeb0ee83ee26eeb9ed;
    decBuf[4554] = 256'h16ed7fecf6eb0deb6feadfe92eea33ebf8eca9ee32f0cbf03ff019ef59eeaaed;
    decBuf[4555] = 256'h8bede1ed2fee77eeb7eef2ee6fef22f0c8f060f19bf189f158f149f13cf148f1;
    decBuf[4556] = 256'h69f15ff156f17ff1b4f1fff131f216f2ccf15ef1bbf024f073ef9eeed4ed52ed;
    decBuf[4557] = 256'h99edddee38f178f383f5c7f50ef515f339f180f028f1f3f21ff595f6e9f7abf7;
    decBuf[4558] = 256'h73f7daf6abf6d5f649f7f7f7d4f864f97ef9d8f8bff765f6daf55cf5cff5c3f6;
    decBuf[4559] = 256'ha1f730f87ff8f5f836f9c0f9f5f9e5f925f906f8adf6c5f59bf5a7f66df898fa;
    decBuf[4560] = 256'h0efcdafc9cfcf4fb8ffaa7f9d1f92bfbccfcc5fe91ffcfff97fffefe2cffaaff;
    decBuf[4561] = 256'hb7006501070104003efe8efc56fceffcedfec90079022203ef02aa01d8001800;
    decBuf[4562] = 256'hafff0e0064007e009600550069009e003101e1018802f402e00287027602c002;
    decBuf[4563] = 256'h8903ff0464064b0776079c07bf071e08ad089909f709db09f00894074f067c05;
    decBuf[4564] = 256'ha305970671085d0b4f0d130f660f850e210ce209d6070a074807d108020b0d0d;
    decBuf[4565] = 256'hd90d9b0d630dca0c9c0c720c980c010d9f0d2f0e4e0f0e10771096104010bd0f;
    decBuf[4566] = 256'h0510c710b211901273125411ad0f250e8c0dba0d350f0011b012c9136214ed14;
    decBuf[4567] = 256'h17153e151b153a15e41496141f14b3139f138d137d13c7130a1416140b149d13;
    decBuf[4568] = 256'hdd12261280116a11f4110013a6142f162e175c17321772163815661459131f12;
    decBuf[4569] = 256'ha1112e1151112e126a138e159917fd19981be31b9f1bef19d6187117e6161017;
    decBuf[4570] = 256'h37175917fb16311612155214e91348144b153f169e1648165d1501141913ef12;
    decBuf[4571] = 256'haf132e15f9162e18661833184b1779160616e31502165916a7161e178a171318;
    decBuf[4572] = 256'hd8185a194319ab18fb17251708178b176118f018a2186d17f2158d14a513cf13;
    decBuf[4573] = 256'h8f14c915f01663178617661710175916831581148d132e134a13011436150916;
    decBuf[4574] = 256'hc91631171217f516db16c31682164716a6150f15fb1478154c168817af18d518;
    decBuf[4575] = 256'hf8185a189117da1634167115ba1414147c139013e9135b14e014f214a1141c14;
    decBuf[4576] = 256'h9f138e13f613be1488150a162216e115cd1598154715fd146a1492130213e812;
    decBuf[4577] = 256'h5f134d142a1580156615c014d21334138a13751410169917fe18e61968190e18;
    decBuf[4578] = 256'h1016ac131112311175112e12b7131c15a7157d15bd143d133e12b311dd115012;
    decBuf[4579] = 256'hb912181335131b13a4128e12a212fb12ce135e1444149e135912b8102f0f960e;
    decBuf[4580] = 256'h680e8f0fe8108912a213a1142c15561530150d15ae145814a113cb123c12b911;
    decBuf[4581] = 256'ha111e2111d125312c0119a10cb0e9f0c290b5d0a9b0ab30be40d5a0fae106711;
    decBuf[4582] = 256'ha01107117b10a90f9c0eee0d100d810c9b0ce20c4e0d260eb60e380f800fc10f;
    decBuf[4583] = 256'had0f9b0f090fe20d670c020bbe09e809a80a270cf20dac0e730e740d760b9a09;
    decBuf[4584] = 256'he108a9084209cd094b0a720ac3092509cf08b508cd0839094c09f308ff07c506;
    decBuf[4585] = 256'h4a054b041d044405ea067308d809630a9009370896060d05740445046f049604;
    decBuf[4586] = 256'h73049603cc0215022d02f0020f046905f405ca050a058a03bf018a0052001f00;
    decBuf[4587] = 256'haa0029019c01bf01de01c201dc01f3010902a7019b0041ffa0fda7fbdbfa9dfa;
    decBuf[4588] = 256'hb6fb1bfd5ffe86ffadffb9fe9cfd8ffce1fbc1fb51fc08fddefda7fef5feaefe;
    decBuf[4589] = 256'h17fe18fd23fc07fb47fadef9bff9dbf9c1f909fa75fa4dfb16fccdfce4fc22fc;
    decBuf[4590] = 256'hcefad0f8f4f6bff587f554f5dff55ef6d1f639f759f73cf7eef677f636f64af6;
    decBuf[4591] = 256'ha3f615f79af7acf77bf7d9f66df659f6d6f6caf7bef8def887f868f7c2f539f4;
    decBuf[4592] = 256'h3af3aff2d9f24cf3b5f3d4f3b8f335f330f23cf15ef0ceef1df064f0fbf036f1;
    decBuf[4593] = 256'h24f1f4f0c7f0d5f02af1cff175f2e1f21cf32ef33ef34df33ff3baf2f5f1d6f0;
    decBuf[4594] = 256'hc9efa7ef05f042f1bdf2bcf38df3bbf215f18cef27ee3fed18eca5ebf7ead7ea;
    decBuf[4595] = 256'h67ebefece8ee4cf1e7f232f366f2b5f0bceee0ec30eb17eae4e9ccea47ec12ee;
    decBuf[4596] = 256'hc3ef4cf1e5f159f187f0c7ef5eefffee56ef3cef95eed3edb3ecf3eb16ecb4ec;
    decBuf[4597] = 256'hb7edabee49eff3ee08ee2eec52ea1de975e8a8e88fe9b6ea10ecb1ed59eef2ee;
    decBuf[4598] = 256'h21efa2ee96eda2ec07eb7ee97fe8f4e7c9e7d6e810eadfeb90ed18efb1efe0ef;
    decBuf[4599] = 256'h0def01ee0ced6eec18ecfeeb28ebece971e80ce781e653e7f9e863eb47ee72ef;
    decBuf[4600] = 256'h17ef20ee80eb06e90fe82fe7fbe730e948ea47eb2fec56ed63ee11eff2ee28ee;
    decBuf[4601] = 256'ha0eca7eacbe812e84ae849e9ebeae4ec38ee75ee3dee3eed9deb14ea15e9e7e8;
    decBuf[4602] = 256'h0eea00ecdced8def35f036ef95ed0ceca7ea1cea46ea9febe4ec0bee7eee5bee;
    decBuf[4603] = 256'hbdedf4eca5ecbdec80ed6bee48efd8eff2ef7befe4ee33ee8ded9fec82eb29ea;
    decBuf[4604] = 256'h41e9c3e8cfe995ebc1edccef20f15ef1b5f050ef0cee39ed13ed7bed59ee95ef;
    decBuf[4605] = 256'h67f074f1ddf1bdf12df142f026efb2eed5ee34efc4ef47f0ffef68ef69ee75ed;
    decBuf[4606] = 256'h55edabed96eeb3ef73f0dcf07df0b3efc8eeebedceede8edbeeec1efb5f053f1;
    decBuf[4607] = 256'he3f131f219f2d9f176f1f9f0a8f05ef086f03cf127f244f351f4b9f4d9f483f4;
    decBuf[4608] = 256'h98f37bf26ef1c0f022f03ff059f0cff03cf1c5f142f2b4f2fef25bf3b0f3bbf3;
    decBuf[4609] = 256'h61f3abf28cf17ff0d1efb1efb4f034f2fff333f54cf67ff651f626f6b3f54bf5;
    decBuf[4610] = 256'hecf496f4b0f4f7f463f514f6baf6fbf6e7f66af6b7f541f500f5ecf4fef4eef4;
    decBuf[4611] = 256'hdff407f5bdf5a8f6c5f7d1f8f4f895f8ccf7adf6edf584f525f542f590f537f6;
    decBuf[4612] = 256'hf9f619f872f95afa81fba7fbcafb6bfbdbfa25faaef96df9a8f901fa73fa9ffa;
    decBuf[4613] = 256'hadfaa0faabfa05fb8bfb2cfc6dfc32fc91fb25fb11fbd6fbf5fc4efedafeaffe;
    decBuf[4614] = 256'ha3fdf4fc96fcecfcd7fdf4feb3ffd6fff9febdfd96fc23fc46fc62fdbcfe0000;
    decBuf[4615] = 256'h2701e7015002ee027d03cc03b4031d03f6017b007cfff1fe1bffdbffcf00ec01;
    decBuf[4616] = 256'hf802a70345040e059105d80597050e052504090396027302d2029b0386042405;
    decBuf[4617] = 256'hed057006b706f8060c07d60685061e06a50575058305c60533069b06dd061a07;
    decBuf[4618] = 256'h5107ab073008d1083d09a0098e093c09d508270881071507da061007e3071f09;
    decBuf[4619] = 256'h9a0aff0b440d6e0dae0c740bf9099408660890085009fe095d0a400a260a9d0a;
    decBuf[4620] = 256'h8b0ba70cb40d1d0e7f0d420c1b0ba80a110bee0bb80c3a0d220d8b0cb30b5d0b;
    decBuf[4621] = 256'h770bee0b850c5d0d260edd0e540f950f5a0fb90ecb0dee0c980cb20cf90c900d;
    decBuf[4622] = 256'hcb0d250e550ebd0e350fa70fb50f8d0f080f430ec10d790d640dc60d670efe0e;
    decBuf[4623] = 256'haf0ff60f0c10d10f540fe20eb60ec30e180f910fe20ff10fe40fa70f860fa40f;
    decBuf[4624] = 256'hd20ffb0f11100a10f80f1f106210b41001111f11f11096102910a50f4b0f1a0f;
    decBuf[4625] = 256'h0c0f340f700fa70fc50faa0f700f3c0f350f6d0fde0f9010071148115c116e11;
    decBuf[4626] = 256'h9e11e811101235121412a6113e11fb10d710f81052118f11f2111a123e124912;
    decBuf[4627] = 256'h2b12d91176111811c410a310c110ee1028113e112a113d1137113c1153114f11;
    decBuf[4628] = 256'h24110811e410e0101f11a811a7125613f4134a143014e9137d13421354138413;
    decBuf[4629] = 256'hce1311141d14d0134e138a12d3115c11f010dc10121184112612e8126b13e213;
    decBuf[4630] = 256'hf7139513f41232127b110411c310b01009117b110012a01263134e14ec147c15;
    decBuf[4631] = 256'h6215eb142914091349129b11fd10e010fa1012117e112f1204130714b6141415;
    decBuf[4632] = 256'hbe14d313771233116010ed0f5510331136126f13ee13c71319133c1239118b10;
    decBuf[4633] = 256'h6b108810a210ba10a4109010ea109c11d112f813b8144f1433134011ec0f330f;
    decBuf[4634] = 256'hfa0e930f7b104e115b12c312e3128d12d6117110720f8b0e0c0ecc0ec00fdd10;
    decBuf[4635] = 256'he9115212f3119d111a1174103310f80f7b0f090f4a0ec70d800d6a0dcc0d6d0e;
    decBuf[4636] = 256'h300fe70f5d107310ea0f250f3a0e5d0dcd0cb30cfa0c910df30d050ef50dc90d;
    decBuf[4637] = 256'ha10dad0db80dc20ddd0dd50dbe0db80d8c0d370d820ccb0b240b8d0a790aaf0a;
    decBuf[4638] = 256'h210bc30b2f0c430c0d0c9b0bf90a620ab1093a09fa080d098a093d0ae30a7b0b;
    decBuf[4639] = 256'hb60b5c0b680a2f090808fb06d80637073a082e09cc09220a080a6209cb084108;
    decBuf[4640] = 256'hc40793078507ad07e90720082a082108c6075907d5067b062a061b060e060206;
    decBuf[4641] = 256'h0d062b0646064e060b068205d1042b0415049f0463051a06910625064d051104;
    decBuf[4642] = 256'h3e037e02a102000390034704bd04fe0412050005af042a0465037a02dc018601;
    decBuf[4643] = 256'h38014f019001cb01010231025e0286027a0259022702f901bf018b0131017c00;
    decBuf[4644] = 256'h90ff35fe4dfdcefc41fd7bfef6ff5b01e70168010f0011febdfc88fb50fbe9fb;
    decBuf[4645] = 256'hd1fca3fd63fe12ffb0ff7900c700df001c00c9fe27fd9ffba0fa71faf0fa63fb;
    decBuf[4646] = 256'h11fc70fc53fc05fc5ffb9cfa19fad2f9bcf9d0f929fa5afaa4fab1fabdfac8fa;
    decBuf[4647] = 256'haafa58fac9f9f1f8eff740f7e1f6c5f67cf751f81bf9d1f919fad8f94ef966f8;
    decBuf[4648] = 256'hc8f7fff6b0f699f6aef6c2f6d4f604f731f759f77df75cf716f78df6b5f5b3f4;
    decBuf[4649] = 256'hbff3e1f251f237f220f260f2c3f263f3fbf384f4def4adf446f498f3c2f26cf2;
    decBuf[4650] = 256'h52f299f230f36bf37df3ebf2ecf1f7f01af0fdef80f085f179f217f334f37df2;
    decBuf[4651] = 256'h49f122f015efaceecceee9ee37ef7eefbfefd3ef2cf05df06cf05ef0f1ef32ef;
    decBuf[4652] = 256'h7bee75edc7eca7ec8bec0ded13ee4cef1ff0dff076f05aef00ee5fec46eb13eb;
    decBuf[4653] = 256'h9eebc5ec6bee14ef47ef18ef46ee39ed8bec2cecd6ebf0ebd8ebeeeb01ecefeb;
    decBuf[4654] = 256'hdfebeeebc6ebbaebc5ebbbebb2eba9eb93eb8cebabebc7eb0aec6eec96ecbbec;
    decBuf[4655] = 256'hc6ec6cece6eb22eb37ea59e9cae87be893e82ae9dbe981eaedeadaea80eaeee9;
    decBuf[4656] = 256'h3de9f6e8e1e81be999e92beab4ea31eb83eb91eb69ebfcea3cea51e9b3e823e8;
    decBuf[4657] = 256'h09e8afe872e991ea51eb74eb55ebfeea13ea36e9a6e858e86fe807e9b7e95eea;
    decBuf[4658] = 256'hcaeaddeaa8ea57ead2e955e924e9bde895e8b9e806e974e916ea82eabdea17eb;
    decBuf[4659] = 256'h27eb71ebceebf3ebe8eba2eb19eb8fea5aea49ea76eaeeea1feb69ebfcebacec;
    decBuf[4660] = 256'h53ed15ee2feeb9edcbec6feb87ea09eae2e905ea64ea81eacfea16ebaeeb37ec;
    decBuf[4661] = 256'hfcec7eed96edaced71ed3bedeaeca0ec93ec9fecc0ec2eedb3ed0cee3dee4cee;
    decBuf[4662] = 256'h3eee63eeb0eeceeed7ee9dee2cee39edd0ecb0ec40ed2bee09ef98efe7efcfef;
    decBuf[4663] = 256'h63efdaee39ee76ed28edb1ecf2eca2eda8ee9cef3af057f0d4ef2eef40eee1ed;
    decBuf[4664] = 256'h37eeeeee23f09ef19df2cbf2a1f2e1f1a8f0d5ef62ef3fefddef6df0bbf0d3f0;
    decBuf[4665] = 256'hbdf0d1f04ef121f224f318f438f4e2f3c2f269f1c7ef1fefecee77eff2f0bdf2;
    decBuf[4666] = 256'hf2f30bf53ef556f4dbf210f156f01ef01df11bf3f7f4a8f650f71df735f663f5;
    decBuf[4667] = 256'h56f462f342f325f374f3bbf327f489f406f578f5c2f5cff5dbf5a4f586f5a2f5;
    decBuf[4668] = 256'hfdf59af632f7bbf7cdf77cf7bcf69cf5ddf4e8f3c9f31ff4d6f4dbf515f73cf8;
    decBuf[4669] = 256'h49f9f7f956fa73faf0f91af9def7b7f6f7f51af6f7f66df838fa6dfb15fc48fc;
    decBuf[4670] = 256'h60fb8efa34f94df8cef7f5f75df8fbf8fef938fb0bfccafcedfccefc77fcf5fb;
    decBuf[4671] = 256'hddfbc7fbdbfbedfbfdfbeefb31fccffc92fd7dfe5affb0ff96ff7eff3eff2aff;
    decBuf[4672] = 256'h60ff70ff7fff56ffe9fe65fe2ffe60fe02fff0ff0c01cc017b029a024402f601;
    decBuf[4673] = 256'h7f013e017901f601a9024f03e6037004a504d604c7049f0463040004bd03b103;
    decBuf[4674] = 256'he8036a04e704790502065c06ce067007dc073e085008de075907b9064c063906;
    decBuf[4675] = 256'h4b069c0603074607b30755081809cf09750ae10a1c0be70a950a4c0a090afd09;
    decBuf[4676] = 256'h1e0a780a150bad0b840c4e0d9c0db40d730dea0c6c0c1b0c0c0c4f0ced0c840d;
    decBuf[4677] = 256'h350eac0ec10eae0e780e270efb0d080e450ea80eea0ede0ee90ecb0ec20e1d0f;
    decBuf[4678] = 256'hbb0fa81086118912f1121113bb1238129211fa104a1032109e104f1154124813;
    decBuf[4679] = 256'he6133c14ee1348130713f3124d13ff137614b7145514b413c6122812d2112012;
    decBuf[4680] = 256'h25131a143615a9158615e8141f143413d512f21274131b140915e615af163217;
    decBuf[4681] = 256'h79178f17a2174917f816cb16a31667163016d6155015d314611418145b14e014;
    decBuf[4682] = 256'ha5155b1602176e1781174c17da1690164d161116321650167d16b716ec160017;
    decBuf[4683] = 256'h52179f17e517491871181c188d17dd160716b115ff1576168f174f18fd185c19;
    decBuf[4684] = 256'h06194f18d8174117df16f0166217c9170c18001887171517ae168616f3167817;
    decBuf[4685] = 256'hf5172618fa17b717c317e4173e18ab189c1809185817b2167116d316bc179918;
    decBuf[4686] = 256'h6219e5199e1906192f186517ae163816f7150a161c162d169416f1162e177b17;
    decBuf[4687] = 256'h99174717e4165116c715b61507168c165017d317eb17aa1720177f163f162b16;
    decBuf[4688] = 256'h3d166e165f16011694152d15b414a41478146b1477149814de146715f0154916;
    decBuf[4689] = 256'h7a1630169d15ed1417148713391321130b136d13c71318147f14a71483142014;
    decBuf[4690] = 256'h7213cc128b127712ad12fe12481370137c1387137d13ab1392133113b8120612;
    decBuf[4691] = 256'h5f111e1132118b11fd110c12ae11f8104210cb0fe00f6a10e71059114a11d210;
    decBuf[4692] = 256'h1f10490fb90ed30eeb0e570fb90fa80f770f4b0f080fe30e040f360f2d0f140f;
    decBuf[4693] = 256'ha40ed10d070d1c0c7e0b9b0b1e0cc40c5b0dbd0d880dd50cd00b960ac3095009;
    decBuf[4694] = 256'hb909960a5f0bae0bc50b030b4c0a7609e60864084c083608fc07ea07b907c807;
    decBuf[4695] = 256'hd507f907ee07e407c907c107c807dd07ca078c0711074c0695051e05dd041805;
    decBuf[4696] = 256'h4e057f055205f5045704c00385039703c803f403cc038f0300037702d6019501;
    decBuf[4697] = 256'ha901de017002fa0253034303dc02130210016200c4ffe1ff97009d019102f002;
    decBuf[4698] = 256'h99027a012100dcfe09fee3fd4cfeeafe40ff26ff80febdfd6ffd27fd68fda3fd;
    decBuf[4699] = 256'hb5fd84fd3bfdddfcd1fc08fd26fd41fd18fdb6fc59fc04fce3fbd9fbbefb63fb;
    decBuf[4700] = 256'hc5fa03fa4cf904f945f9f6f9ccfa95fbaffb68fb4ffa42f94ef8b0f7cdf71bf8;
    decBuf[4701] = 256'hc1f802f9eef871f8bff7e9f659f60bf6f3f534f647f636f605f6bbf578f584f5;
    decBuf[4702] = 256'he7f595f66bf7fbf749f802f814f7f7f5ebf43cf4ddf3faf349f490f4a5f492f4;
    decBuf[4703] = 256'h80f44ff405f4ddf370f309f3abf26ff27af2fcf279f3ebf3f9f39cf3e6f22ff2;
    decBuf[4704] = 256'h89f173f1fcf19df235f397f361f3cff21ef278f137f172f1a8f1f9f108f2c5f1;
    decBuf[4705] = 256'h58f10ef1e6f00af157f175f16cf143f1e1f084f078f057f075f07ef054f0f3ef;
    decBuf[4706] = 256'h7bef09efa2ee94eed1ee34efacefddefceef8befeeee82ee6eee80ee12efeaef;
    decBuf[4707] = 256'h40f05af013f050ef9aee23ee0dee6fee10ef7cef90ef5aefa8eed2ed09ed52ec;
    decBuf[4708] = 256'h0aecf5eb08ec62ecd4ec3bedb3ed45ee80eeb6eee7eebaee78ee3beec2ed50ed;
    decBuf[4709] = 256'h06eda9ec6cec77ec81ecafecf9ec3fed7fedb9eda2ed72ed3aede7ecc6ecf8ec;
    decBuf[4710] = 256'h38ed93ed00ee0feee7ed7aedd7ec40ecb7eb81eb91eb16ec6fecc1ec0aedc7ec;
    decBuf[4711] = 256'h8bec6aec4cec9eec17ed89edd2ede0ed8bed28edb0ec5eec15ec3dec61ecaeec;
    decBuf[4712] = 256'hf4ec22ed5bed81ed7aed67ed4bedfeecc7eca9ec7cec84ec8bec77ec3fecfbeb;
    decBuf[4713] = 256'ha9eb88ebe2eb80ec6ded4beea1eebbee15eefcecefeb41eb21ebeaeb0aed16ee;
    decBuf[4714] = 256'h0bef2aef0def8bee44eed7ed9dedaeed5ded4eed26ed02ed23ed55ed95edf0ed;
    decBuf[4715] = 256'h5deea6eee9ee26ef05efbfee7fee45ee4deea6eefbee48ef66ef14ef9bee29ee;
    decBuf[4716] = 256'hdfed22eed8eec3efe0f0edf155f236f2dff128f182f0ebef61ef2cef5defc4ef;
    decBuf[4717] = 256'h72f018f1aff1eaf1d8f167f1fff0bcf098f0e5f07bf13ef2c0f237f34df3ebf2;
    decBuf[4718] = 256'h91f2fff1c4f1d6f127f28ef222f35cf34bf31af3b3f28af2aff212f3daf3ddf4;
    decBuf[4719] = 256'h8cf52af60df6bff518f581f41ff4e9f3d9f3e8f3f5f332f469f4c3f430f57af5;
    decBuf[4720] = 256'h87f57bf55af578f5eef5c2f68bf742f85af8edf73df767f6d7f5bdf504f6c7f6;
    decBuf[4721] = 256'h7ef754f8e3f866f94ef9e2f880f8dff79ef7d9f756f809f9aff947fa82fa93fa;
    decBuf[4722] = 256'h83fa74fa67fa2afa09fafff9e4f90dfa42fa80facafae8fa03fb2dfb70fbd4fb;
    decBuf[4723] = 256'h4dfcdffc41fd53fd63fd37fd0ffdd2fcb1fc93fc9cfcb5fcf9fc39fd62fd96fd;
    decBuf[4724] = 256'hc6fd24fed2fea8ff7100f400ac0093ff3afef5fc23fcfcfbabfc07fe4bff7200;
    decBuf[4725] = 256'h320155013501df005c0045002f006a009f00f10058018001a401af0191017601;
    decBuf[4726] = 256'h5d01470140015f01650155011001a2005800800036018a028804dc059506cd06;
    decBuf[4727] = 256'h68052404a902aa017b01fa016d021b037a039703b103f80339049b0418058a05;
    decBuf[4728] = 256'hf105340640064b062d06db0578050005af04a004c8041d05ac053506d6066d07;
    decBuf[4729] = 256'hd00705081508cc073907af06560646068f063d07e307a608290940090009c508;
    decBuf[4730] = 256'h4808f607ad078407a907e0074e08d3085009c1090b0a330af709c00966094109;
    decBuf[4731] = 256'h4c097e09d0091d0a4f0a460a0d0aba0957092f096c09fb09d20ad50b3e0c9d0c;
    decBuf[4732] = 256'h460c900be90a7d0a420a780aa90ad50afd0af10ad00ada0ae30afc0a5d0bbb0b;
    decBuf[4733] = 256'h100c730cb60cc20ca10c5b0cf60b990b740b690bc30b490cc60c170d260de30c;
    decBuf[4734] = 256'h760c0f0cb10ba50bdc0b360cbb0c380daa0d110e1f0efa0d970d040d540cdd0b;
    decBuf[4735] = 256'hc70bdb0b7c0c130d9d0dd20de20db60d8e0d820db90d130e680e890e6b0e060e;
    decBuf[4736] = 256'h730dea0cb40ca40cee0c4b0db90d200e7d0ea20ead0eb70e9b0e830e6c0e2e0e;
    decBuf[4737] = 256'hf50da20d550d4b0d660da00df30d2a0e200e170e0e0ef80d0c0e130ee00d940d;
    decBuf[4738] = 256'h260dbf0ccd0c3a0df90d190fd90f41102210920f730eb30d040da50c890cd70c;
    decBuf[4739] = 256'h4e0dba0df50d070e170e080ee00dec0de10dff0d1b0e230e0c0ece0d630dde0c;
    decBuf[4740] = 256'h850c540c630cc10c460de70d530eb50ea30e520eeb0d3d0dc60cb10cc40cfa0c;
    decBuf[4741] = 256'h4b0d5a0d670d5b0d500d6e0d9c0dc50dbd0d720df00c960c450c360c790cff0c;
    decBuf[4742] = 256'h7c0dcd0df90db60d310d6c0cb60b3f0bfe0aea0a440bb50b3a0cdb0c470d5b0d;
    decBuf[4743] = 256'h490d180db10c530c2f0c500c960cfa0c220dfe0c9b0ced0b760b0a0bf70a2c0b;
    decBuf[4744] = 256'h5d0ba70bea0b0e0c190c0f0ce10b870b1a0bb20a550a610a820ac80a080b200b;
    decBuf[4745] = 256'hec0abc0a840a7c0a9e0ad70afc0a030bd70a8e0a700a670a800ab40ae40af70a;
    decBuf[4746] = 256'hf20ac30a7f0a2d0aca096c092f090e09040920093809400955094e093d092e09;
    decBuf[4747] = 256'h2009240947097109770953090d09770889072b070e0790073708ce087f09c609;
    decBuf[4748] = 256'hb0094e09f508a4083c081408f007fb07190822080908a8072f07be0674068106;
    decBuf[4749] = 256'hbe06210749075507080786062d061c062b06a40636079807aa079a073207ba06;
    decBuf[4750] = 256'h4806e1059e0561052a050c0503053d05ae054006a206d806a7062206a5053305;
    decBuf[4751] = 256'he904f7040305f804da047604fd03ac038003c30330049704f5040105ca047004;
    decBuf[4752] = 256'h0304b903910385037a039803d703110437043004f80396031e03cc0283029002;
    decBuf[4753] = 256'hb402010347038703b103b803a3036b03fb0289020402ab017a016b019301d001;
    decBuf[4754] = 256'h070225021c02e201ae017e015e015901540161016e019101d60130029e02ca02;
    decBuf[4755] = 256'h8702d101e600090079ff93ff3900270104022102d3012d013f00a1ff4aff64ff;
    decBuf[4756] = 256'hacffedff0000eeffdeffb2ff6fff32ffe5feb3feaafec3fe24ffb8ff1a002c00;
    decBuf[4757] = 256'hdaff38ff75fef3fdacfdc1fd4bfeebfe58ffbaffa8ff57ffd2fe31fe9afd10fd;
    decBuf[4758] = 256'hdbfcaafcb9fcabfc9ffc94fc8afc93fcbcfc00fd64fda7fdccfd95fd27fd67fc;
    decBuf[4759] = 256'h7cfbdefa4efa34faaafa42fbf2fbc8fc58fd72fd5afdeefc3efc68fb9ffa1cfa;
    decBuf[4760] = 256'hd5f9eaf925fa7ffaaffabefacbfad8faf9fa03fbf9faaffa41fa9ff9dcf85af8;
    decBuf[4761] = 256'h12f8fdf75ff800f997f921fa56fa46fa1afaa1f90ff986f82cf8dbf7ccf7f4f7;
    decBuf[4762] = 256'h31f87ef888f86df833f8e0f7bff7ddf71df857f86ef822f88cf7c9f612f69cf5;
    decBuf[4763] = 256'hb1f513f691f602f74cf759f74df716f7bcf667f6eef55cf5d3f479f469f4d0f4;
    decBuf[4764] = 256'h49f5dbf564f653f622f6d8f57af56ef579f56ff542f5c6f401f44af303f3eef2;
    decBuf[4765] = 256'h77f35ff43df5ccf51bf6a4f50df535f46cf3b5f26df258f26bf2c5f237f39ef3;
    decBuf[4766] = 256'h16f426f418f4baf31cf385f24af238f269f2eef247f398f3c5f39df378f341f3;
    decBuf[4767] = 256'h0ff3cff296f252f224f20cf213f236f26ef293f2a8f2aef287f263f24cf226f2;
    decBuf[4768] = 256'h0cf2fef1e9f1ddf1f6f112f23cf26ff276f263f23cf203f2def1e5f1dff1e4f1;
    decBuf[4769] = 256'he9f1c9f1a3f19ef1abf1ebf174f2d6f20cf3dbf274f2c6f14ff1e3f0cff029f1;
    decBuf[4770] = 256'h7af1a6f1e9f10ef219f25ff268f270f24af2e3f17cf139f12df164f1bef113f2;
    decBuf[4771] = 256'h34f23ef210f208f21ff241f279f2bdf2c6f29df24af2bbf132f1fcf02df1b2f1;
    decBuf[4772] = 256'h9af277f307f455f43ef47bf390f2b3f123f109f120f1b8f141f2bef251f3b3f3;
    decBuf[4773] = 256'h0cf41cf40ef4b0f343f3dcf299f28df2daf234f3b9f312f423f414f406f4e2f3;
    decBuf[4774] = 256'hedf31ff43af453f45bf438f419f41ff42ef46af4c5f402f539f557f54df524f5;
    decBuf[4775] = 256'h0ef5ebf4ccf4d2f4cdf4e4f41bf54ff59bf5f5f519f624f62ef638f640f656f6;
    decBuf[4776] = 256'h5df657f63bf60df6e1f5e7f50af650f6d2f64ff7c1f728f835f829f808f8aef7;
    decBuf[4777] = 256'h72f751f747f762f7acf7f2f720f85af861f876f87cf88df8a6f8d9f8fcf80ef9;
    decBuf[4778] = 256'h09f9dbf8a2f88cf893f8d8f84ef9e0f943fac0faf0fa1dfb2afb06fbe5fa9ffa;
    decBuf[4779] = 256'h5ffa25fa0ffa31fa8ffa22fbabfb28fc59fc68fc25fcd0fb83fb65fb6efbb8fb;
    decBuf[4780] = 256'h26fc8efcd1fcf5fc00fdcefcc5fcbdfce2fc20fd6afd88fd91fd79fd44fd2ffd;
    decBuf[4781] = 256'h4ffda3fd10feb2fe1fff81ffb6ffa6ff7aff37ffe2feabfe8dfea8fee2fe35ff;
    decBuf[4782] = 256'h98ffdbff17003800420039001000eaffbaffa7ffcfff1c007f0012017401aa01;
    decBuf[4783] = 256'h99016d012a010601110143019501f8013b025f0254024a024102490260029002;
    decBuf[4784] = 256'hc802fd021f033e03390334031c030703fc02ff02150340036c039e03dc031604;
    decBuf[4785] = 256'h4b047b048d0488046e0445044a047804d6044e05a005cc05a4053705cf048d04;
    decBuf[4786] = 256'h8004b7042505aa052706ba06f40606071707ea068d0650061906fb0504063e06;
    decBuf[4787] = 256'h8106d4060b0729073207290713070c071207180727072c0717071b0725075407;
    decBuf[4788] = 256'hbb074008e1084d0960092b09b9081708ab0770078207b2073708910802094c09;
    decBuf[4789] = 256'h74098009a10997097c0953090f09bd08700852085b08a508ff083c0989099309;
    decBuf[4790] = 256'h8a099209b809da09060a220a130afb09e609db090f0a530a920abc0ab40a840a;
    decBuf[4791] = 256'h580a3c0a2d0a3b0a470a3c0a310a2e0a3d0a640ab80a560bc20bfd0beb0b9a0b;
    decBuf[4792] = 256'h330bba0a890a7b0a880aac0ae30a010b1d0b250b0f0b230b360b690bc20b170c;
    decBuf[4793] = 256'h380c560c3a0c010cea0be30b030c400c7a0c640c260cbb0b360bdc0aed0a190b;
    decBuf[4794] = 256'hac0b350c6b0c9c0c8d0c4a0c3e0c330c3d0c580c710c4c0c370c180cfc0b2a0c;
    decBuf[4795] = 256'h620c970cb90c9a0c450cd80b8e0b810ba50b080c660cd30cff0cf20ce60caf0c;
    decBuf[4796] = 256'h690c3b0c120cfc0bf50bfb0bf50bf00be20bcd0be00b0e0c460c990cd00c020d;
    decBuf[4797] = 256'hf90ccf0c6e0c100ca30b3c0b2e0b3b0b5c0ba20be10bfa0b110cfc0bdd0be20b;
    decBuf[4798] = 256'he80bff0b1c0c300c250c160cf60bc70bb50baf0b950b910b7b0b510b290b060b;
    decBuf[4799] = 256'hd30abe0a9f0a830a920aa00abe0af80a630bad0b0a0c2f0c0e0cc80b3f0b8e0a;
    decBuf[4800] = 256'he8097c0968099e09ef09560ab40ac00a9f0a590a190af009f8090c0a2b0a480a;
    decBuf[4801] = 256'h4d0a360a200afd09cb098d094209fc08e108d908ef081f093f092309ea089808;
    decBuf[4802] = 256'h610857088408df084c09960989094c09bd083408da07a9077d07a507e2070308;
    decBuf[4803] = 256'h21082a0822080b08e907b1079a078607730784079d07a20795076307fc069406;
    decBuf[4804] = 256'h52061506360654068206bb06d206d906eb06f106e206c10682061d06da05b605;
    decBuf[4805] = 256'hed0547069c06a7067506ec053b05950454046804e5047705d905eb05ba057105;
    decBuf[4806] = 256'h1305ef04fa04180533052b050505c7046d0430040f04f103e803cf03c803cf03;
    decBuf[4807] = 256'he103fd0317042e042a041e04ff03e103d503bd039b0371033303f902c502b002;
    decBuf[4808] = 256'hb602d302e202d402ae026b023e0235025b029902d202e902c70275021202b501;
    decBuf[4809] = 256'h78016d0177018001570131010f01fc0018015b019b01d501dc01ba0169011c01;
    decBuf[4810] = 256'hd600a8008f00880081007b00750070006b0067004400ffffa5ff38ff0bfffefe;
    decBuf[4811] = 256'h53ffccff3e00a500cd00a9005c00020094ff4bffd2fe81fe37fe0ffe34fe6bfe;
    decBuf[4812] = 256'hc5fe19ff66ff70ff55ff0bffb1fe44fedcfd7ffd5afd65fd97fd0efe80fee7fe;
    decBuf[4813] = 256'hf4feb8fe3ffe8cfde6fc7afc3ffc51fc81fcaefcf1fc2dfd4efd6cfd75fd6dfd;
    decBuf[4814] = 256'h48fdfcfca2fc35fcebfb8dfb81fba2fbe8fb28fc41fc2afcfafbc2fb8efb94fb;
    decBuf[4815] = 256'hb4fbc5fbcafb8efb22fbbbfa43fa12fa3efa81fad6fa23fb2dfbfffaa5fa37fa;
    decBuf[4816] = 256'heef9c6f9d2f909fa4ffa6afa72fa5cfa39fa0efafdf9e3f9b0f965f90bf99ef8;
    decBuf[4817] = 256'h54f82cf838f89bf8f8f866f9aff9d7f9b3f966f9f8f891f84ef82af81ff83df8;
    decBuf[4818] = 256'h58f871f896f882f849f8f7f794f751f745f766f798f7eaf70bf801f8e6f7acf7;
    decBuf[4819] = 256'h86f79bf7baf7e2f7e7f7a1f733f7ccf66ef64af66bf6b1f603f73af744f729f7;
    decBuf[4820] = 256'hdff699f66bf652f63cf635f62ff61ef62df64df66bf68ef6a5f687f64df614f6;
    decBuf[4821] = 256'hc1f5a0f596f58df5a6f5daf5eff502f612f6f9f5cff59df551f50bf5ddf4c5f4;
    decBuf[4822] = 256'hccf40af544f587f5c7f5cff5aaf55ef5f0f4a6f499f48df4c4f40af538f550f5;
    decBuf[4823] = 256'h58f528f5fcf4d5f4bbf4b6f4d4f4d8f4cdf4b8f48cf43bf41af438f48af419f5;
    decBuf[4824] = 256'h7bf5b1f5a1f53af5a6f444f4ebf3dbf307f42ff46cf48df497f4a0f4b9f4def4;
    decBuf[4825] = 256'h0ef53af51ef5dbf489f426f4fef33bf488f4f6f45df56af546f5f9f49ff44af4;
    decBuf[4826] = 256'h3ff435f463f48cf4b1f4c6f4e5f4ebf4faf411f51ef52af53bf525f500f5d2f4;
    decBuf[4827] = 256'h8df44df445f45bf4a7f415f55ff5bcf5c9f5a8f576f548f50ef507f51bf52ef5;
    decBuf[4828] = 256'h4af564f55ff55bf567f56af57af594f597f58ef58bf578f57bf59bf5cef50bf6;
    decBuf[4829] = 256'h35f63cf635f62ff613f618f62ff633f637f63bf61ff60bf616f632f66cf6d7f6;
    decBuf[4830] = 256'h3ff781f7bef7b3f76df71bf7a2f651f642f66af6d7f65cf7d9f74bf877f84ff8;
    decBuf[4831] = 256'h12f8aff76cf748f769f7aff713f88cf8bdf8e9f811f9edf8ccf89af86cf843f8;
    decBuf[4832] = 256'h4af86df8b1f816f959f97df988f96af94ff957f97cf9c8f922fa5ffa80fa76fa;
    decBuf[4833] = 256'h36fafcf9e5f9dff9fef947fa79fa94fa9dfa86fa71fa84faa0fad9fa1cfb4afb;
    decBuf[4834] = 256'h73fb99fb9ffbbffbdbfbeafbeffbebfbc0fb8dfb6bfb65fb97fbfefb66fcdefc;
    decBuf[4835] = 256'h2ffd3efd31fddcfc79fc36fc12fc33fc8dfc12fdb3fd1ffe81fe6ffe3efed7fd;
    decBuf[4836] = 256'h5ffd0efde1fc09fd5efdc1fd3afe6afe97fea4feb0fed1fe03ff55ffa2ffc0ff;
    decBuf[4837] = 256'h93ff38ffcbfe64fe3bfe60fed9fe8cff3200c90004011601e5009b0059003400;
    decBuf[4838] = 256'h1300f5ffdaffd2fff7ff3500a00007018001b101dd01b501780141010f010601;
    decBuf[4839] = 256'h1f016201d9014b02b202da02e602af027d023d0214020c022102400251026102;
    decBuf[4840] = 256'h78029e02eb024e03ab0300040b04c50373031003e8020c036f03e8035a048604;
    decBuf[4841] = 256'h5e042104ea03cc03d503ee031304440463047f04b7040a0557058905a4057b05;
    decBuf[4842] = 256'h2805f104d30401053b057e05ac0593055f052f0541058a050c068a06db06af06;
    decBuf[4843] = 256'h5106cc0572056205c90577061d0789079d076707f60671063b060b0637067a06;
    decBuf[4844] = 256'hb606ed060b0739078307dd07320869085f080d0894072207d806cb0620078307;
    decBuf[4845] = 256'h1608510863083208e807a5079907ba0714088108e908f608ea089d082f08e507;
    decBuf[4846] = 256'hd807fc0749088f08bd08c508a0086f0869087a08b20805093c0946092b091209;
    decBuf[4847] = 256'hec0801092d09540978096a092a09ea08c108ab08db08130948096a0957093009;
    decBuf[4848] = 256'h160908090d0947099109c309030a0b0af509d2099a0956093b0912090a092d09;
    decBuf[4849] = 256'h7109c409270a690a760a550afb098d09440951097509d809360a730a680a0e0a;
    decBuf[4850] = 256'h88092f091f092d09a609180a440a510a150a9c094a093c096409d109560aaf0a;
    decBuf[4851] = 256'he00ab30a560ae9099f095c093809430925092e0936094d099809f209470a7e0a;
    decBuf[4852] = 256'h880a480aed09800919090c09000921096709a609bf09c709c009880962092409;
    decBuf[4853] = 256'hea08e308dc08e208fe080e091c09420966098f09cd09f709e009a2093709b208;
    decBuf[4854] = 256'h3508e407d50718086d08d0082d0982098d09830956091c09d808860839081b08;
    decBuf[4855] = 256'h24083d088108c108d908d208af085e082708090812082b084208480836081a08;
    decBuf[4856] = 256'h0a0818083e0877089c08a30877082308ce076b0743074f077007b607e407ec07;
    decBuf[4857] = 256'h0208ee07db07ca07bb079a078e076b07380723070407f3060d071b0727073307;
    decBuf[4858] = 256'h2207f906d206a30684068a06ae06ce06fd061c070b07fc06c906a70694068e06;
    decBuf[4859] = 256'h890684065e061106c4057e0563057c05bf0511065e0668064d061306c1057405;
    decBuf[4860] = 256'h6a0573057b05a105a705950584056a05530557054c0533051705e504b504a204;
    decBuf[4861] = 256'ha704cb040705310556054f0530050905db04af048704640443041d040304f503;
    decBuf[4862] = 256'h0204250445045b046e047204620459044c0437041d04e803b403840365035f03;
    decBuf[4863] = 256'h8d03d203ff0318040204a8035303f002ae02a102d8021e037103a8039e035e03;
    decBuf[4864] = 256'h1303b9027d025c0266029302ac02b402ad0281024e021e02f301d601d101d601;
    decBuf[4865] = 256'hda01ee01f101fa01fd01f501e501c501920162012a010401e200e800ee00f300;
    decBuf[4866] = 256'h01010d010a01ff00e900cf00b7009b00780057002900fdffd6ffc6ffc2ffd7ff;
    decBuf[4867] = 256'hfaff110015000200d4ffa8ff76ff53ff41ff19fff5fed5fec0fecbfef9fe3eff;
    decBuf[4868] = 256'h7eff96ff71ff17ff92fef1fdb0fd9dfdd2fd24fe8bfeb3fea7fe5afe00fec3fd;
    decBuf[4869] = 256'ha2fdacfdc8fdd0fdc8fd8afd40fde6fcc2fca1fcabfcd8fc02fd18fd1ffd0cfd;
    decBuf[4870] = 256'hf0fcd7fcadfc86fc62fc2ffc0cfcedfbe8fbf7fb17fc35fc39fc2efc00fcb4fb;
    decBuf[4871] = 256'h6efb1cfbe5fac7fad0faf9fa1ffb41fb47fb36fbfefabbfa7bfa41fa2afa31fa;
    decBuf[4872] = 256'h44fa55fa6ffa73fa5efa43fa0efadaf99cf962f93df928f92ef93ff96df999f9;
    decBuf[4873] = 256'hb5f9baf9a3f963f911f9c4f86af846f825f82ff85df875f89bf8bdf8c3f8b3f8;
    decBuf[4874] = 256'h99f85df813f8cdf77af759f74ff759f761f786f7a9f7c8f7e4f7f3f7f8f7e3f7;
    decBuf[4875] = 256'ha9f74ef7f9f696f653f65ff680f6b2f604f725f72ff714f7ebf6a7f67af650f6;
    decBuf[4876] = 256'h3af633f62df61cf621f60af6fdf509f60cf616f61ef607f6def5b7f589f576f5;
    decBuf[4877] = 256'h70f56bf566f562f54ff53df53af532f53ff559f56af574f577f54ff51df5ecf4;
    decBuf[4878] = 256'h9bf464f45af451f46af480f495f4a8f4b9f4bef4b9f4b5f49af473f44ff41cf4;
    decBuf[4879] = 256'hfaf3f4f3e3f3e8f308f40df418f42af41af40cf404f4eff3e0f3d8f3c3f3baf3;
    decBuf[4880] = 256'hc7f3caf3d9f3eff3e0f3cef3b4f386f367f36df37cf393f3c2f3c8f3c3f3a9f3;
    decBuf[4881] = 256'h64f31ef302f3e9f20ff34df387f3bbf3ddf3cbf3aff395f359f330f319f304f3;
    decBuf[4882] = 256'hfef204f313f32af351f36af38bf3a8f3a4f3a1f398f36cf34df331f303f3f0f2;
    decBuf[4883] = 256'hebf2dbf2e0f206f32af35df39bf3b3f3acf397f35ff32bf308f3f5f2fbf21ff3;
    decBuf[4884] = 256'h3ff36ef39af3abf3baf3bff3a1f386f36df34bf33df341f345f35ef38df3aff3;
    decBuf[4885] = 256'hcef3eaf3eff3fdf30af406f411f41af411f40af411f402f404f40df40bf40ff4;
    decBuf[4886] = 256'h21f428f448f47bf49ef4c9f407f520f527f52ef528f517f512f504f508f51cf5;
    decBuf[4887] = 256'h34f55df590f5b2f5d1f5f9f5fef50cf618f61cf62ef64af655f667f689f6a0f6;
    decBuf[4888] = 256'hcff607f72df74ff762f75cf74df752f75ef781f7b4f7d7f7f6f712f821f838f8;
    decBuf[4889] = 256'h67f893f8c6f8f6f808f90ef913f90ff924f94ef981f9b1f9ddf9e3f9f2f900fa;
    decBuf[4890] = 256'h0dfa37fa80fac6fa06fb2ffb46fb3ffb2cfb10fb01fb18fb3efb81fbd3fb36fc;
    decBuf[4891] = 256'h79fcb5fcd6fce0fceafce1fcdafce1fce7fc0efd3cfd75fdc7fd14fe5afe9afe;
    decBuf[4892] = 256'hb3febafec1feaefea9feb8fecffefefe36ff6bffa9ffe2ff26006600a000c500;
    decBuf[4893] = 256'he700ee00f300ee00fc0011013c017a01b401e80118022b023c0255026d029302;
    decBuf[4894] = 256'hcb02000330036803ac03d90302040a0411040b040504140435047404b4040f05;
    decBuf[4895] = 256'h4c056d058b0594058c0593059a05b905e10519064d069906cb060b0724073a07;
    decBuf[4896] = 256'h4f0749072c072707350742076d07b607e8073a087108a308be08c608b008b708;
    decBuf[4897] = 256'hbd08c308f10829095e099b09b409ad09c109c809d809070a3f0a640a940a9b0a;
    decBuf[4898] = 256'h950a900a950a990abc0aef0a110b490b6f0b830baf0bcb0bd00be70bec0be80b;
    decBuf[4899] = 256'hf20b020c100c380c6a0c8d0cb80cc90cce0ce60cfb0c060d2d0d510d5f0d7c0d;
    decBuf[4900] = 256'h900d930d9d0da00d920da30dbf0dda0d0e0e520e6d0e960e8f0e6d0e660e550e;
    decBuf[4901] = 256'h460e700e970ebb0eee0e100f160f270f370f320f470f530f480f580f5b0f5e0f;
    decBuf[4902] = 256'h810fa50fbc0fe20ff20fe40fe80fe40fda0ff00ffe0ffb0f1a10271023103c10;
    decBuf[4903] = 256'h521054106c107510671074107b1079109710b510b910d110c810ae10b210ae10;
    decBuf[4904] = 256'h9a10b210c210bf10dc10ef10f91022113e11431164115f11441133111011e710;
    decBuf[4905] = 256'hec10fc100a11411175118a11a911a4118a11731155112b1125112a1125114c11;
    decBuf[4906] = 256'h7011741192119e119311a311a6118e11911183115b114a113b112d1153117711;
    decBuf[4907] = 256'h8e11b511b0117d115a113b1108111d1130114111651172115511511131110311;
    decBuf[4908] = 256'hfc10eb10d210d610ca10b610c810cb10bd10ca10be109e108710691037102210;
    decBuf[4909] = 256'h1c1016103a105a105f106a1052102310ca0f750f3e0f340f2b0f330f670f7c0f;
    decBuf[4910] = 256'h820f7d0f590f130fe10eb40e7a0e630e4f0e300e400e460e380e3c0e210ef30d;
    decBuf[4911] = 256'he10db90d950d870d720d570d540d310d080deb0cd20c9f0c8a0c6b0c440c3f0c;
    decBuf[4912] = 256'h310c1b0c1f0c0e0ce50bc90b910b4d0b200bf60ad10aca0ac40aa80a980a780a;
    decBuf[4913] = 256'h490a2a0a190aff09040ae609bc097e093309d9089d087c0872088d08a608ad08;
    decBuf[4914] = 256'ha70887083e08f807940751071407dd06d306ca06c206ba06b406940662063206;
    decBuf[4915] = 256'hed05ad0573053f050f05fc04e004d004cc04ae047c044b040704c7038d036803;
    decBuf[4916] = 256'h530340032f030b03eb02bc02840250021202e801c301a1018101650141012a01;
    decBuf[4917] = 256'h0c01ea00c0008d004f001600e1ffa3ff6aff44ff14ff01fff0feebfef0feecfe;
    decBuf[4918] = 256'hd0fe9cfe49fee6fda4fd4ffd2efd10fd19fd21fd1afd13fdf3fcccfc9efc66fc;
    decBuf[4919] = 256'h31fcf3fbbafb76fb48fb1ffb18fb11fb17fb1dfb03fbd0fa92fa48fa02fad4f9;
    decBuf[4920] = 256'habf995f980f96df951f942f918f9f1f8d7f8aef891f878f84ef827f803f8d9f7;
    decBuf[4921] = 256'hbdf7aef797f78af76ff741f709f7d5f6a4f66cf656f641f63bf640f631f611f6;
    decBuf[4922] = 256'hf3f5b9f56ff551f523f5faf401f5edf4daf4d4f4bbf49af485f462f438f411f4;
    decBuf[4923] = 256'hd9f3a4f382f363f352f357f352f356f35af334f306f3e6f2a9f26ff258f244f2;
    decBuf[4924] = 256'h31f22bf21cf217f213f2f0f1d0f1b2f178f14ff138f124f12af146f137f129f1;
    decBuf[4925] = 256'h1cf1e2f0a8f074f043f024f02af025f033f050f04cf049f04cf021f0f5efd9ef;
    decBuf[4926] = 256'h96ef69ef50ef2bef24ef43ef54ef59ef67ef49ef26ef06efcfeea9eea2ee83ee;
    decBuf[4927] = 256'h7dee8dee7fee72ee7eee65ee5cee70ee5eee52ee50ee32eef2edd6ed9ded86ed;
    decBuf[4928] = 256'ha9edbbedd7ed06eef3edd7edb3ed77ed4ded55ed5ced7bedaeeda7ed94ed78ed;
    decBuf[4929] = 256'h40ed0bed12edffec1bed3fed3bed36ed3aed14ed04ed12ed05ed09ed22ed0ced;
    decBuf[4930] = 256'hfeec00edebecf3ec16ed1aed2fed43ed31ed22ed19edf7ece9ecf6eceaecf5ec;
    decBuf[4931] = 256'h11ed15ed26ed42ed46ed58ed74ed60ed4fed4ced26ed17ed25ed29ed4ced7fed;
    decBuf[4932] = 256'h86ed99edb5eda5eda1edaded9aed9eedb3edb6edc9edecede7edf5ed0aeeffed;
    decBuf[4933] = 256'h09ee2cee30ee45ee68ee6dee7aee95ee8aee94eea2ee9aeea1eec1eec6eedbee;
    decBuf[4934] = 256'h0def22ef41ef5def58ef5def59ef45ef50ef78ef89efadefe0efe7ef06f022f0;
    decBuf[4935] = 256'h32f052f078f088f096f0abf09ff09cf0b2f0b4f0d1f004f126f15ef193f1a7f1;
    decBuf[4936] = 256'hbaf1d6f1d1f1dff1f4f100f218f247f25cf288f2baf2cff2e2f2fef203f31af3;
    decBuf[4937] = 256'h49f35cf38ef3bef3def3faf313f418f436f451f462f48bf4bef4e0f4fff432f5;
    decBuf[4938] = 256'h46f572f59af5a9f5d3f5faf509f620f647f656f66df693f6adf6e0f61ef747f7;
    decBuf[4939] = 256'h7cf7acf7bef7dbf7eaf7eff7fbf716f82ff858f895f8cff804f942f96bf990f9;
    decBuf[4940] = 256'ha5f9abf9b1f9c0f9cef9f4f92dfa61fa91facafaeffa11fb31fb4dfb71fba4fb;
    decBuf[4941] = 256'hc6fbe5fbf6fbfbfb09fc27fc42fc76fcbafcfafc34fd59fd6efd80fd86fd95fd;
    decBuf[4942] = 256'hbffdf2fd30fe59fe7efe85fe8bfe91feb5fef1fe4cffa1ffeeff0c0027001f00;
    decBuf[4943] = 256'h0800010014003c007400b700e5001f01440174019401c601e901080224022902;
    decBuf[4944] = 256'h37024c0267029c02d002010339035e0381039303bb03d403f503240443046a04;
    decBuf[4945] = 256'h84049b04b904dc04fc0422055b058005a205c205d305ec050d0622064c067f06;
    decBuf[4946] = 256'ha106cd06e906f906fd060a0716073c077507a907f507270842085b0853083f08;
    decBuf[4947] = 256'h450856086f08a208e00809094d097b099309aa09b109aa09bb09cb09cf09f609;
    decBuf[4948] = 256'h190a310a5f0a8b0a9c0ac00ae00af50a180b390b3d0b500b620b650b790b910b;
    decBuf[4949] = 256'h9a0bbf0bd90bf00b160c3a0c510c800c930c990ca80ca30c9f0cb20ccb0ce70c;
    decBuf[4950] = 256'h190d4a0d500d6c0d710d630d780d940da50dd40df60d090e1a0e150efe0d020e;
    decBuf[4951] = 256'h060e020e310e540e730ea50ec80ec20ed20ecd0eb60ec30ecf0ecb0eed0efb0e;
    decBuf[4952] = 256'h000f220f300f3d0f580f6a0f6d0f7b0f790f680f6e0f740f6f0f870fa00fa30f;
    decBuf[4953] = 256'hbd0fc70fbe0fd20fda0fd30fea0ff40fe50ff20ff00fdd0fe50fe70fd80fee0f;
    decBuf[4954] = 256'hf70ffa0f14102510221030102910131010100810f30f01100410f80f07101110;
    decBuf[4955] = 256'h05101d10281025103310301011100510f10fd90fdc0fd90fcc0fe10fe40fd70f;
    decBuf[4956] = 256'he30fe50fdb0feb0fed0fd30fcf0fb30f890f780f680f5b0f700f7b0f780f8e0f;
    decBuf[4957] = 256'h850f6e0f5e0f440f250f200f1c0f0b0f140f0c0fea0edc0ecf0eac0eb10eac0e;
    decBuf[4958] = 256'h990ea40e940e740e700e550e350e3a0e2e0e160e120e040ee20dd40dbf0da40d;
    decBuf[4959] = 256'ha00d910d710d6d0d520d390d300d210d0f0d080df50ccd0cbc0ca30c820c7e0c;
    decBuf[4960] = 256'h7a0c690c660c520c2f0c180cea0bbe0ba20b920b720b6e0b6a0b580b550b470b;
    decBuf[4961] = 256'h2a0b170bf70ac80aa90a8d0a690a5b0a4e0a3b0a2a0a140af409df09c4099d09;
    decBuf[4962] = 256'h8e0980096b095f09470924090409de08af0890087f0866086a08660853084108;
    decBuf[4963] = 256'h1f08ec07ca079e077607670750073b0727071607fa06e606ce06b806a4068c06;
    decBuf[4964] = 256'h640647061906ee05d105b805a1059405810568055205330515050105e904c704;
    decBuf[4965] = 256'haf04920467044b0431041a040504f203d903bd039a0370035403300319030403;
    decBuf[4966] = 256'hf102d802c202ae0291027e02650243022c020e02f301d401b6019b017b015d01;
    decBuf[4967] = 256'h420131011b010d01fa00e000c100a30080006900540040002f001f000b00eeff;
    decBuf[4968] = 256'hcbffabff85ff6bff54ff47ff34ff29ff1aff05ffeefed2feaffe8efe79fe66fe;
    decBuf[4969] = 256'h54fe3efe2afe13fefdfde3fdcafdbbfda7fd9afd89fd76fd5efd48fd2efd16fd;
    decBuf[4970] = 256'h00fdf2fcdffccffcbcfca9fc94fc7afc68fc5ffc4bfc39fc23fc0ffcf2fbd7fb;
    decBuf[4971] = 256'hbffbaffba6fb9efb97fb8dfb7ffb6bfb54fb38fb1dfb12fb02fbfafaf7faebfa;
    decBuf[4972] = 256'hd8fac6faa7fa89fa7efa73fa70fa73fa70fa64fa55fa37fa1afa0efafdf9f9f9;
    decBuf[4973] = 256'h02fafaf9eef9e4f9cef9baf9acf99cf991f993f98af97ff978f96bf960f95bf9;
    decBuf[4974] = 256'h52f94bf94df942f93af936f926f91ff925f924f91ff920f911f9fff8f3f8e0f8;
    decBuf[4975] = 256'hd8f8dbf8ddf8e7f8f3f8eef8e4f8daf8c7f8baf8bcf8bff8c5f8d4f8cef8c4f8;
    decBuf[4976] = 256'hbbf8a9f8a2f8adf8aff8bbf8caf8c8f8bff8b7f8a3f89bf899f897f8a1f8b4f8;
    decBuf[4977] = 256'hb7f8b9f8c4f8bef8c0f8c8f8c0f8bcf8bbf8acf8a2f8a7f8a6f8b0f8c5f8cef8;
    decBuf[4978] = 256'hd5f8ddf8d2f8c8f8caf8c2f8c0f8caf8cdf8d5f8e0f8dcf8ddf8e3f8e0f8e3f8;
    decBuf[4979] = 256'heef8f3f8fbf804f9fef8fdf802f9faf8fef80bf90cf914f922f91df91ef929f9;
    decBuf[4980] = 256'h25f92bf93af93cf93df945f93bf93cf945f944f94bf958f95af95cf961f95ff9;
    decBuf[4981] = 256'h66f976f97df98bf99af99df997f991f97ff978f983f989f9a0f9bcf9c7f9d2f9;
    decBuf[4982] = 256'hdbf9cdf9c0f9c2f9c0f9c6f9d6f9dcf9e6f9f6f9f4f9f6f9fff9faf9f8f9fff9;
    decBuf[4983] = 256'hf9f9faf905fa06fa10fa23fa30fa37fa3dfa33fa2bfa2cfa28fa2ffa41fa54fa;
    decBuf[4984] = 256'h64fa73fa71fa6cfa67fa57fa50fa52fa51fa5ffa79fa84fa8dfa9bfa99fa96fa;
    decBuf[4985] = 256'h94fa8efa90fa9bfaa0faa7fab2faaefaa9faadfaaafaadfabafac0fad0fadffa;
    decBuf[4986] = 256'hddfadefae3fadffadbfae1fae4faebfaf8fa06fb13fb24fb22fb20fb1efb12fb;
    decBuf[4987] = 256'h0afb0efb12fb22fb36fb43fb53fb5afb54fb4efb50fb49fb4afb58fb64fb76fb;
    decBuf[4988] = 256'h8bfb9afba7fba9fb9afb88fb81fb7bfb85fb9ffbbafbdafbeffbf3fbe8fbd9fb;
    decBuf[4989] = 256'hd0fbcdfbdefbedfb03fc17fc1ffc1cfc1ffc1dfc1efc2dfc3bfc47fc56fc58fc;
    decBuf[4990] = 256'h5afc5bfc54fc58fc66fc72fc84fc99fca2fcaafcacfcaefcb0fcb9fcbefcc2fc;
    decBuf[4991] = 256'hc9fccffcd7fce6fcf1fcfbfc0efd1bfd1efd24fd22fd24fd25fd2dfd3cfd52fd;
    decBuf[4992] = 256'h60fd6dfd70fd69fd5ffd5afd59fd63fd78fd92fdb1fdc6fdd2fdcefdd2fdc9fd;
    decBuf[4993] = 256'hc1fdc8fdcffdddfdecfdf7fd05fe15fe1bfe21fe2afe2bfe2afe2bfe32fe3efe;
    decBuf[4994] = 256'h53fe67fe74fe85fe87fe89fe87fe86fe8afe97fea5feb7fec3fec9fecbfecafe;
    decBuf[4995] = 256'hcbfed0fed9feeafef9fe07ff13ff18ff1fff21ff27ff31ff3bff48ff58ff5eff;
    decBuf[4996] = 256'h64ff6dff75ff7aff83ff87ff88ff8bff90ff96ffa3ffb9ffcdffdfffebffe9ff;
    decBuf[4997] = 256'hdfffdaffd8ffe3fff5ff0f0027003d0046004300370028002200280036004c00;
    decBuf[4998] = 256'h66007800870096009800960098009a00a300ab00b200bc00c500c800cf00db00;
    decBuf[4999] = 256'he300e700f400fc0006011001190123012c01330138014101450148014f015401;
    decBuf[5000] = 256'h5a0163016d01780183018a018b018e0191019701a501b301c201d501e301e501;
    decBuf[5001] = 256'he701e501e301e801f001fc010b02150221022c022b022702280229022e023b02;
    decBuf[5002] = 256'h4d025e0275028502880285027e0278027a0282029102a302af02b902bf02c102;
    decBuf[5003] = 256'hbc02c102c502cb02dc02e802f30201030d030e0316031a031b03230324032a03;
    decBuf[5004] = 256'h34033b0341034d03560357035b035f035e0367036d037703890395039b03a503;
    decBuf[5005] = 256'hab03a203a703a803aa03b603c503cf03de03e503e303dd03d903d103dd03ec03;
    decBuf[5006] = 256'hfe0318042a043304300428041804110413041c0431043a04420449044b044904;
    decBuf[5007] = 256'h4e04530458045e04650468046f047304780485048f048d04950494048d048904;
    decBuf[5008] = 256'h8604830490049e04a304b204b804b304b104ac04a804b104bd04c604d604dc04;
    decBuf[5009] = 256'hda04d504cd04c004c104c004c104ce04d204d104d804dc04d804df04e204df04;
    decBuf[5010] = 256'he504e304db04de04df04dd04e304e404e404eb04e804e204e404e404df04e404;
    decBuf[5011] = 256'he404dd04d904d604d204d804d904d804e204e604dd04de04d704ca04c804c304;
    decBuf[5012] = 256'hbb04bc04c004bf04c904ca04c704ca04c104ae04a604a4049e04a804b004af04;
    decBuf[5013] = 256'hb304aa0497048a04830478047e0483048204860485047a0475046e0463046104;
    decBuf[5014] = 256'h6004570454044f0449044b0449044104400439042c04260416040b0409040b04;
    decBuf[5015] = 256'h09040e0412040c040604f903e903e303dd03db03e003e203d803cf03be03a403;
    decBuf[5016] = 256'h9a0390038e039503a1039f03a103950380036c035f0357035e03640366036a03;
    decBuf[5017] = 256'h630354034603330320031e031c0316031b0319030f030b030203f602f402ef02;
    decBuf[5018] = 256'he602e502dd02d002ca02c602c102c202c102b902b202a5029302870281027f02;
    decBuf[5019] = 256'h8b029302950291027e026602500242023f024b025a02600265025d0247023102;
    decBuf[5020] = 256'h1d02150217021e02240229022702200213020502fb01f601f701f601f701f301;
    decBuf[5021] = 256'hee01eb01e301d401ce01cc01c801cc01cb01c401c101b801b401b501b401b501;
    decBuf[5022] = 256'hb801b501ad01a8019f0199019501940195019901950188017a016e0166016701;
    decBuf[5023] = 256'h6e017e019101990197018801720158014e0144014d015a016b01750173016a01;
    decBuf[5024] = 256'h59014801390133013c014a0154015a0158014e01410136013101380143014b01;
    decBuf[5025] = 256'h4c014b013c012a011f0118011a0123012e0133013101290123011c011d012101;
    decBuf[5026] = 256'h2601280126011c010d0103010101000107010e011901180111010601fb00f400;
    decBuf[5027] = 256'hf300fb000601100112010601f900e600d300cc00d300dd00ec00f700f900ed00;
    decBuf[5028] = 256'hd800c300bc00b900bb00c900d600de00d900d200c500b800b000af00b000af00;
    decBuf[5029] = 256'hb200b100ab00a00094008d0089008a0092009700940092008b0085007f007e00;
    decBuf[5030] = 256'h7d007d00780076006e00610059005200500054005a005b0056004e0042003300;
    decBuf[5031] = 256'h2d00280030003b003f00400036002a001e0011000c000d000f00130014000e00;
    decBuf[5032] = 256'h0100f5ffe7ffe1ffdfffe4ffe8ffeffff0ffedffe6ffd9ffc7ffbbffb0ffaaff;
    decBuf[5033] = 256'hb0ffb4ffb6ffb5ffacffa2ff9bff95ff93ff98ff99ff97ff8fff87ff7aff6eff;
    decBuf[5034] = 256'h69ff67ff66ff65ff61ff58ff4dff46ff41ff40ff41ff46ff49ff45ff3dff2eff;
    decBuf[5035] = 256'h20ff17ff0fff0eff12ff13ff12ff11ff0bfffefef0fee3fedbfeddfedefee2fe;
    decBuf[5036] = 256'he3fedefed4fec8feb9feb3feb5febdfec5fec9fec5febbfeacfe96fe88fe80fe;
    decBuf[5037] = 256'h7dfe7bfe85fe87fe89fe81fe77fe6ffe67fe60fe5dfe5cfe56fe54fe53fe4bfe;
    decBuf[5038] = 256'h45fe40fe3cfe37fe35fe2ffe29fe26fe20fe18fe15fe10fe09fe09fe06fe00fe;
    decBuf[5039] = 256'hf8fdf0fde9fde8fde6fde5fde7fde5fdddfdd5fdc6fdb3fdabfda4fda6fdacfd;
    decBuf[5040] = 256'hb1fdb0fdaefda7fd97fd8cfd82fd7afd7bfd7afd7bfd7afd70fd63fd58fd47fd;
    decBuf[5041] = 256'h41fd3ffd41fd46fd50fd4ffd46fd3efd2ffd1cfd14fd0dfd0ffd15fd13fd0ffd;
    decBuf[5042] = 256'h0afdfefceffce9fce0fcdbfcddfcd6fcd2fccffcc4fcbffcbefcbdfcbcfcbdfc;
    decBuf[5043] = 256'hb5fcabfca1fc91fc8afc8cfc8bfc8cfc94fc8dfc7ffc73fc61fc50fc4efc50fc;
    decBuf[5044] = 256'h56fc5efc5cfc58fc52fc43fc35fc30fc28fc23fc27fc24fc20fc1dfc12fc07fc;
    decBuf[5045] = 256'hfffbf8fbf4fbfafbf5fbf4fbf7fbedfbe1fbd5fbc8fbc3fbc4fbc0fbc1fbc7fb;
    decBuf[5046] = 256'hc4fbbdfbbefbb1fba3fb9efb92fb8efb8cfb86fb87fb88fb82fb7efb7ffb77fb;
    decBuf[5047] = 256'h71fb6cfb61fb55fb4efb47fb46fb4bfb48fb49fb4afb3dfb2ffb2afb1efb17fb;
    decBuf[5048] = 256'h1bfb1cfb24fb2ffb2bfb21fb16fbfffaf0faedfaeafaecfaf7faf9faf7faf6fa;
    decBuf[5049] = 256'he5fadbfad5faccfacdfad8fad9fad3fad2fac7fabffabefab3fab4fac1fabffa;
    decBuf[5050] = 256'hbbfab9faaefaa6faa2fa9afa98fa9ffa9ffaa1faa7faa3faa0faa3fa9bfa98fa;
    decBuf[5051] = 256'h9ffa99fa92fa95fa8dfa8cfa91fa8efa8ffa95fa95fa94fa93fa87fa83fa87fa;
    decBuf[5052] = 256'h86fa8cfa9bfa9dfaa2faa3fa96fa8afa8bfa84fa85fa93fa9cfaa1faaefaacfa;
    decBuf[5053] = 256'habfaa9faa2faa1faabfaadfab0fabafab9fabafac0fabffac2facdfacffad0fa;
    decBuf[5054] = 256'hd7fad6fad2fad7fad6fadefaedfaeffaf8fa00fbfefa00fb06fb07fb12fb20fb;
    decBuf[5055] = 256'h21fb23fb2afb26fb2afb32fb35fb3ffb4bfb50fb57fb5efb5dfb63fb70fb75fb;
    decBuf[5056] = 256'h7afb8afb91fb97fba3fba4fba6fbadfbacfbadfbb6fbc1fbcefbe2fbeafbf1fb;
    decBuf[5057] = 256'hfbfbf9fbfbfbfdfbfefb08fc18fc27fc35fc45fc4bfc4dfc56fc57fc5cfc66fc;
    decBuf[5058] = 256'h6cfc76fc80fc83fc8dfc9afca5fcb3fcc2fcc9fccffcd8fcd9fce1fceafceefc;
    decBuf[5059] = 256'hf8fc07fd0dfd13fd1bfd1ffd26fd36fd45fd53fd63fd69fd6ffd78fd7afd81fd;
    decBuf[5060] = 256'h8bfd91fd9bfdaafdb0fdb9fdc4fdc9fdd5fde1fde5fdeffdfdfd05fe0dfe18fe;
    decBuf[5061] = 256'h22fe2dfe3afe43fe48fe4ffe54fe5afe64fe6efe79fe89fe94fe9afe9cfea1fe;
    decBuf[5062] = 256'ha5feb1febafec7fed7fee6fef0fefcfefefefffe06ff11ff1cff28ff33ff38ff;
    decBuf[5063] = 256'h3fff45ff4dff54ff5eff6aff72ff7aff80ff89ff91ff9affa8ffb1ffb9ffc3ff;
    decBuf[5064] = 256'hc7ffc9ffceffd5ffddffe7fff4ffffff09000e00110017001e0026002b003800;
    decBuf[5065] = 256'h4500500058005e00620066006b006b00770085008f009c00a400a500a400a500;
    decBuf[5066] = 256'ha900b200ba00c700d500e300ec00f100f500f100f500fb00000106010e011301;
    decBuf[5067] = 256'h1a0120012c013a0144014a014b01500154015801620169017101770182018a01;
    decBuf[5068] = 256'h8b018c01920193019501a101ac01b401c301c901cb01c901ca01cc01d501df01;
    decBuf[5069] = 256'he801f60102020402080207020302090210021a022602310236023a023b023a02;
    decBuf[5070] = 256'h3d0241024902580266026f02770278027402780279027802800288028b029402;
    decBuf[5071] = 256'h9e029f02a702aa02ad02b102bb02bf02c502c602c902cf02d002d602e202ea02;
    decBuf[5072] = 256'hee02f002ef02eb02ec02ef02f50202030c0315031a031b031203100311031203;
    decBuf[5073] = 256'h1e0329033403400342033703360332032c032f033b0343035003560351034f03;
    decBuf[5074] = 256'h4b034a03500359035f0369036d036903680363035f0365036b036e0372037303;
    decBuf[5075] = 256'h6d036e036f036f0377037d037e03820381037a0376037503730377037f038003;
    decBuf[5076] = 256'h8703860382037f037b03750377037c03800388038b0382037e03790370036f03;
    decBuf[5077] = 256'h720375037f038503840381037a036d036703650367036b037203760377037203;
    decBuf[5078] = 256'h65035f035d035f0363036703630362035d0352034a034503440348034b034e03;
    decBuf[5079] = 256'h52035003460342033c033403350336033303360333032b032603230320032603;
    decBuf[5080] = 256'h2703240324031a030e030503fb02fa02020308030d0313030f030203fc02f302;
    decBuf[5081] = 256'he702ec02f002f102f502f402ec02e402d902ce02d002d102d202d902de02d702;
    decBuf[5082] = 256'hd102cb02c302c202c302c202c702c802c102bf02b502ae02ab02ac02ad02b302;
    decBuf[5083] = 256'hb702b602b402ac029d029b02990298029c029e029c029e029902920290028d02;
    decBuf[5084] = 256'h8e02940292028d028e028b0282027e027a027b02840288028702860280027402;
    decBuf[5085] = 256'h6f026b026c027202760277027b0277026d02690263025f02640269026d027202;
    decBuf[5086] = 256'h6f026502610256024e025002540255025a025c025a02570253024d024c024d02;
    decBuf[5087] = 256'h4c024b024a02470245023f0238023d023f024002430246023f023b0231022d02;
    decBuf[5088] = 256'h2c022b022a022d022d02290225021f02170218021d0223022602260224021f02;
    decBuf[5089] = 256'h12020402ff01fd01ff0109020f0210020b020002f701f001e901ea01f401fb01;
    decBuf[5090] = 256'hfa01f701ee01e201d501cc01cb01d201d901dd01de01d901cd01c201b801b601;
    decBuf[5091] = 256'hb501b601b301b401ae01a201a1019c0198019c019d019e019b01920185017d01;
    decBuf[5092] = 256'h73016f0170017101740175016d0163015c0151014c014e014c01490148014001;
    decBuf[5093] = 256'h3601320129011f011b011a011b011c011b0115010d010101f500ee00e700e600;
    decBuf[5094] = 256'he700e600e000d900d200ca00c500bd00b900ba00b600ae00a6009b0091008700;
    decBuf[5095] = 256'h7e007d007e007d007d0078006f00620057004f004b004700440043003b002f00;
    decBuf[5096] = 256'h230019000f000e00110010000e0009000000f3ffe8ffdeffd9ffdbffd5ffd2ff;
    decBuf[5097] = 256'hceffc2ffb7ffacffa6ffa2ffa3ffa2ff9fff9dff95ff88ff7dff73ff69ff60ff;
    decBuf[5098] = 256'h61ff60ff5eff5bff57ff4fff42ff3aff33ff2cff2dff2aff25ff20ff19ff0cff;
    decBuf[5099] = 256'h04fffdfefefefffefefefffefcfeeffee1fed9fecdfec9fecafec6fec5fec4fe;
    decBuf[5100] = 256'hbcfeb4feb1feaafea6fea9fea7fea4fea3fe99fe8dfe88fe7efe77fe76fe77fe;
    decBuf[5101] = 256'h78fe79fe74fe6efe6afe62fe5afe59fe5afe57fe56fe50fe48fe40fe37fe31fe;
    decBuf[5102] = 256'h35fe38fe3afe3ffe3efe36fe2cfe22fe17fe15fe11fe10fe16fe17fe12fe10fe;
    decBuf[5103] = 256'h08fe02fe01fe00fe03fe07fe06fe00fefafdf2fdeafde3fddffde3fde9fdecfd;
    decBuf[5104] = 256'hebfdeafde4fde0fddafdd2fdd3fdd8fdd5fdd4fdd5fdcdfdc6fdc3fdc2fdc3fd;
    decBuf[5105] = 256'hc9fdcdfdd0fdcffdc9fdc1fdbbfdb6fdb7fdbafdb9fdbbfdbefdbafdb5fdb8fd;
    decBuf[5106] = 256'hb5fdb8fdbbfdbdfdbefdbffdb5fdaefdabfda7fda8fdb0fdb6fdb9fdbdfdbefd;
    decBuf[5107] = 256'hbdfdbbfdb8fdb5fdb8fdb7fdbafdbcfdb6fdb4fdb4fdb4fdb4fdb9fdbdfdc7fd;
    decBuf[5108] = 256'hd0fdcffdd0fdcffdc9fdc5fdc7fdc8fdcdfdd5fddafdddfde0fdddfddcfddbfd;
    decBuf[5109] = 256'hdcfde6fdedfdeefdf4fdf9fdf4fdf2fdf3fdf3fdf8fd03fe0bfe13fe17fe16fe;
    decBuf[5110] = 256'h17fe1afe1bfe1ffe25fe2afe30fe31fe30fe32fe37fe39fe43fe4dfe55fe5ffe;
    decBuf[5111] = 256'h66fe63fe64fe65fe64fe66fe70fe7afe85fe8ffe91fe92fe93fe96fe9bfea6fe;
    decBuf[5112] = 256'haefeb6febcfebefebdfec0fec2fec7fed2feddfeebfef4fef8fefdfe01ff02ff;
    decBuf[5113] = 256'h03ff0aff12ff1aff25ff2dff2eff34ff38ff3dff45ff51ff60ff6aff76ff7bff;
    decBuf[5114] = 256'h7cff7eff7cff80ff85ff8eff9bffa6ffaeffb2ffb8ffc2ffc9ffd2ffe0ffeaff;
    decBuf[5115] = 256'hf3fff8fff9fff8fff9fffdff0600130020002e0038003e004200440048004e00;
    decBuf[5116] = 256'h560061006c00730079007c007f0085008f009b00a700b400b900c200c000bf00;
    decBuf[5117] = 256'hc200c800cf00d900e200eb00f500fc00000105010c0114011e012b0130013401;
    decBuf[5118] = 256'h36013901380139013f014b0156015e016701700173017401770178017a018201;
    decBuf[5119] = 256'h8f019401980199019b019e01a301a701b501bf01c401c901c701c601c701c801;
    decBuf[5120] = 256'hc701cf01d901e001e601ea01eb01ed01f201f801fc01fd01000202020102ff01;
    decBuf[5121] = 256'hfc01fb01fc0102020c0213021c021d021e021f021e021b021c021d021f022002;
    decBuf[5122] = 256'h23022402250220021e021d022102290231023402310230022c02280227022802;
    decBuf[5123] = 256'h2a022f0230022f022e022b0227022802290228022902260222021d0219021602;
    decBuf[5124] = 256'h1902180217021d0220021d021c021b02150213020d020c02090205020002ff01;
    decBuf[5125] = 256'hf901f501f401f501f801f801f401f101f101e901df01dd01d701d401d501d201;
    decBuf[5126] = 256'hce01cd01c801bf01b801b701b301b001af01ab01a701a0019a0192018d018601;
    decBuf[5127] = 256'h8101810180017f017e017b01730169016001590154014d014a01480140013801;
    decBuf[5128] = 256'h35012f012e012f012e01290122011a01110108010001f700ee00e900e600e100;
    decBuf[5129] = 256'he000e000d900d500d200ce00ca00c400ba00b300ad00a500a0009a0094008c00;
    decBuf[5130] = 256'h8b00880083007d0075006d00640061005d005a00590057005100490041003c00;
    decBuf[5131] = 256'h3800370032002c00280022001a0012000d000500fffffafff8fff5fff3fff2ff;
    decBuf[5132] = 256'hefffebffeaffe7ffe1ffd7ffd1ffc8ffc4ffbfffb9ffb7ffb4ffb0ffadffaaff;
    decBuf[5133] = 256'ha6ffa2ffa1ff9bff96ff94ff8fff89ff87ff82ff7cff78ff77ff74ff72ff6dff;
    decBuf[5134] = 256'h6bff66ff64ff5cff58ff53ff51ff4eff4aff44ff3fff3dff3aff3bff3cff3bff;
    decBuf[5135] = 256'h38ff30ff26ff22ff21ff20ff1dff1aff19ff17ff0fff0bff0aff08ff09ff0bff;
    decBuf[5136] = 256'h0cff09ff07ff01fffcfef6feeefeebfeecfeeffeeffeeffeecfee9fee7fee6fe;
    decBuf[5137] = 256'he5fee2fedefedffee0fedffedcfed8fed3fed3fed5fed6fed7fed8fed5fed4fe;
    decBuf[5138] = 256'hd2fecdfecbfeccfeccfeccfecbfec8fec7fecafecbfecafecbfecdfed0fecffe;
    decBuf[5139] = 256'hcefecdfecbfec5fec5fec8fec5fec6fecbfeccfecbfeccfecbfecafec9fec8fe;
    decBuf[5140] = 256'hd0fed6fed5fed4fed5fecefeccfec9fec8fecdfed5fed6fed9fedafed7fed4fe;
    decBuf[5141] = 256'hd3fed1fed2fed4fed7fedafedcfedbfedafedafed5fed6fedefee1fee2fee1fe;
    decBuf[5142] = 256'hdffedcfedbfed7fed6fedafee1fee7fee9fee7fee2fee3fee2fee3fee4fee7fe;
    decBuf[5143] = 256'he9feecfee6fee1fee2fee0feddfee1fee6fee7fee9fee8fee9fee7fee2fee1fe;
    decBuf[5144] = 256'he4fee3fee6feecfee9fee8fee8fee1fee1fee3fee6fee7fee9feeafee9fee3fe;
    decBuf[5145] = 256'hdffedefedffedefee2fee8fee9fee8fee8fee3fee1fee3fee2fee3fee2fee5fe;
    decBuf[5146] = 256'he6fee3fedffedefedffee0fee1fee3fee4fee3fee2fee3fee2fee1fedffee3fe;
    decBuf[5147] = 256'he8fee8fee9fee8fee6fee1fedffee0fee4fee8feebfeeefeedfee8fee9feecfe;
    decBuf[5148] = 256'hebfeeafeedfeeefef0feeffeeffef1feeffeeafeedfeeffef0fef5fefbfef8fe;
    decBuf[5149] = 256'hf9fef8fef6fef3fef6fefafe00ff06ff05ff06ff05fffffefbfefcfefefe04ff;
    decBuf[5150] = 256'h09ff0aff09ff08ff05ff06ff05ff0aff10ff16ff13ff12ff13ff14ff13ff12ff;
    decBuf[5151] = 256'h13ff14ff17ff18ff19ff18ff15ff16ff13ff12ff17ff1fff22ff23ff24ff20ff;
    decBuf[5152] = 256'h1dff1eff1dff20ff22ff27ff2dff2cff26ff21ff20ff20ff22ff28ff2bff2eff;
    decBuf[5153] = 256'h2eff2cff29ff2aff2bff2aff2eff31ff34ff36ff37ff35ff34ff35ff34ff35ff;
    decBuf[5154] = 256'h35ff36ff3bff3dff3bff3aff39ff3aff3cff41ff47ff48ff4aff4bff45ff41ff;
    decBuf[5155] = 256'h42ff44ff49ff4dff53ff52ff51ff51ff51ff52ff55ff58ff5cff5fff65ff64ff;
    decBuf[5156] = 256'h63ff66ff68ff66ff66ff6dff6fff70ff73ff74ff73ff74ff76ff77ff7aff7eff;
    decBuf[5157] = 256'h82ff8aff8eff8dff8cff8dff8cff90ff98ff9bff9eff9fffa2ff9fff9dff9eff;
    decBuf[5158] = 256'ha4ffa8ffacffb1ffb3ffb4ffb7ffb8ffbcffc2ffc7ffc9ffceffcfffcfffcfff;
    decBuf[5159] = 256'hd1ffd4ffd8ffddffe1ffe4ffe8ffebffebffebffedfff0fff2fff9ff00000600;
    decBuf[5160] = 256'h09000a0009000a000d00130019001d002200280029002600290028002a003000;
    decBuf[5161] = 256'h38003e00430047004a004b004d005000540059005f0063006800690069006e00;
    decBuf[5162] = 256'h7000730076007c00840089008e009300970098009b009d009e00a200aa00ae00;
    decBuf[5163] = 256'hb100b200b400b900bf00c100c700ce00d200d500db00dc00dc00e100e900f100;
    decBuf[5164] = 256'hf600fa00fe0001010201060109010b011201160119011f012101240128012d01;
    decBuf[5165] = 256'h33013b0143014a014e0151015101540151015201570159015f0167016d017201;
    decBuf[5166] = 256'h7801790176017c0184018c018f019201940199019a019b01a101a301a801ae01;
    decBuf[5167] = 256'hb201b501b701bc01bd01c101c501c801cc01d101d201d601d901da01de01e201;
    decBuf[5168] = 256'he501eb01ef01ef01f301f401f101f601f801f901fd01020206020b020a020b02;
    decBuf[5169] = 256'h0f021002120219021d021a021d021e021d0220021f021e022002230227022c02;
    decBuf[5170] = 256'h2b022c02300231022e022e023002330235023802390238023702350235023602;
    decBuf[5171] = 256'h3b023d023e023c023c023c0237023602370238023c0241023c023d023e023d02;
    decBuf[5172] = 256'h3c023a0237023c023b02350232022f022d022c022b022c023002310232023302;
    decBuf[5173] = 256'h2d022702260225022202250222022102240220021602120211020f020e020e02;
    decBuf[5174] = 256'h0d020e0207020102ff01fe01fb01fa01f901f701f601f201ed01e901e301de01;
    decBuf[5175] = 256'hdd01db01d801d701d101cf01ce01c801c301c101c001bd01be01bb01b501b101;
    decBuf[5176] = 256'hab01a501a0019a019601970192018c01880182017a017b017c0179017a017601;
    decBuf[5177] = 256'h70016b0160015401560152014c014801450141013c0133012c012d0128012501;
    decBuf[5178] = 256'h25012101190116010f0105010101fd00fc00f900f500ef00e900e200db00d300;
    decBuf[5179] = 256'hce00c900c700c100bc00b800b200a800a100a0009f009e00990095008d008500;
    decBuf[5180] = 256'h80007a00740070006b0063005e0057004b00470042003e003a00390034003000;
    decBuf[5181] = 256'h2a0023001d0017000f000c000b0007000200fafff2ffebffe5ffdcffd5ffd1ff;
    decBuf[5182] = 256'hceffcdffc8ffc2ffbeffb9ffb0ffa9ffa8ffa2ff9dff9aff94ff8eff88ff80ff;
    decBuf[5183] = 256'h7bff76ff6fff6bff67ff5fff59ff56ff52ff4fff4dff46ff42ff38ff32ff2eff;
    decBuf[5184] = 256'h28ff21ff1dff18ff12ff11ff0fff0aff04fffefefafef7feeffeeafee9fee3fe;
    decBuf[5185] = 256'hdcfed6fed2fecffec9fec1febefebdfeb7feb2feb2feabfea7fea3fe9bfe95fe;
    decBuf[5186] = 256'h96fe94fe8dfe8bfe86fe80fe7efe78fe73fe72fe70fe6afe69fe63fe5cfe5afe;
    decBuf[5187] = 256'h57fe4ffe4cfe49fe48fe45fe43fe42fe43fe3efe38fe36fe31fe2dfe2afe26fe;
    decBuf[5188] = 256'h23fe22fe20fe1bfe1bfe16fe12fe13fe0efe0cfe0dfe06fe04fe05fe06fe06fe;
    decBuf[5189] = 256'h06fefffdfdfdfafdf6fdf3fdf4fdf1fdf1fdf0fdeafde9fdeafde3fde4fde7fd;
    decBuf[5190] = 256'he1fddefde4fde3fde1fde2fde3fde2fde3fde2fdddfddefdddfddcfdddfddbfd;
    decBuf[5191] = 256'hd8fdd7fdd6fdd5fdd6fdd5fddafddcfddafddbfdddfddbfdd6fddbfddcfdd9fd;
    decBuf[5192] = 256'hdafdd9fddafddefdddfddcfdddfddcfdddfde2fde1fde2fde6fde5fde6fdeafd;
    decBuf[5193] = 256'he8fde9fdeffdeefdf1fdf7fdf2fdf3fdf9fdf8fdf8fdfefdfdfdfcfd00fe01fe;
    decBuf[5194] = 256'h04fe0afe0bfe0dfe12fe14fe17fe1afe19fe1afe1cfe1ffe22fe26fe25fe26fe;
    decBuf[5195] = 256'h2afe2ffe35fe3dfe40fe41fe45fe48fe4bfe51fe53fe5afe5efe5ffe65fe69fe;
    decBuf[5196] = 256'h68fe68fe6cfe6ffe76fe7efe7ffe84fe8afe89fe8dfe99fe9efea2fea9feaafe;
    decBuf[5197] = 256'haefeb9febafebbfec2fec5feccfed4fed5fedcfee0fee0fee4feeffef1fef5fe;
    decBuf[5198] = 256'hfffe05ff09ff12ff15ff1bff22ff25ff2bff31ff35ff3aff3eff41ff42ff49ff;
    decBuf[5199] = 256'h4fff56ff5cff62ff68ff6fff73ff7bff7eff83ff8bff91ff96ff98ff9dffa3ff;
    decBuf[5200] = 256'ha9ffadffb3ffbaffbcffc1ffc8ffceffd1ffd4ffd8ffdbffe1ffe7ffebfff5ff;
    decBuf[5201] = 256'hfcfffdff03000a000b000f0017001a001d002300220025002b00300036003a00;
    decBuf[5202] = 256'h3d0043004b005000530058005a0060006300620065006b006e00700076007c00;
    decBuf[5203] = 256'h7f00800084008a008f00930098009a009b009c009f00a300a700aa00ad00b300;
    decBuf[5204] = 256'hb500ba00bc00bf00c200c600c900cb00cc00cf00d100d600da00de00df00e400;
    decBuf[5205] = 256'he600e900ec00f000f100f200f300f300f400f700fb0000010101050109010c01;
    decBuf[5206] = 256'h0b010e0110011101140118011b011c0120012301240124012401240129012a01;
    decBuf[5207] = 256'h29012d0130012d01320136013701360139013b013c013d014001400143014601;
    decBuf[5208] = 256'h48014601450147014a0147014801470148014d014f014e014f0152014f015201;
    decBuf[5209] = 256'h5301500155015501550155015601540153015201530155015601550155015001;
    decBuf[5210] = 256'h4f0150014f014e014f0152015101540151014d014a014b014a01490147014601;
    decBuf[5211] = 256'h4701470145014201430140013e013b013a01390139013401320131012e012d01;
    decBuf[5212] = 256'h2c012a012901280124011f011e011c011b011c01190116011601110110010e01;
    decBuf[5213] = 256'h090108010901050102010001fb00fa00fa00f500f600f300ef00ec00ec00e700;
    decBuf[5214] = 256'he600e400df00de00da00d600d500d600d100d000ce00cb00ca00c800c500c200;
    decBuf[5215] = 256'hc000bb00bc00b600b200b100b200af00b000af00ad00aa00a600a1009f009a00;
    decBuf[5216] = 256'h99009a0099009700960093008f008c008b008700840082007f00800081007b00;
    decBuf[5217] = 256'h780077007500740075006e006e006d006800660061005b005e005f005a005800;
    decBuf[5218] = 256'h5700540053004d004b004b004b004600450043003e003d003900360036003300;
    decBuf[5219] = 256'h32002f002f002e002d002a002b0028002400210021001e001b00150013001500;
    decBuf[5220] = 256'h14001000110010000d000c000a000700030002000100feffffff0000fffffdff;
    decBuf[5221] = 256'hfcfff7fff7fff6fff7fff7fff5fff4fff5fff0ffeaffebffecffe9ffe7ffe6ff;
    decBuf[5222] = 256'he9ffedffeaffebffeeffebffe9ffe8ffe9ffe9ffe9ffe8ffe7ffe4ffe2ffe1ff;
    decBuf[5223] = 256'he0ffe1ffe3ffe6ffe3ffe6ffe5ffe1ffe2ffe6ffe7ffe9ffeaffedffeeffebff;
    decBuf[5224] = 256'he7ffe6ffeaffebffe9ffe9ffeeffefffeeffeffff0ffeffff1fff4fff3fff4ff;
    decBuf[5225] = 256'hf5fff2fff5fff7fffafff7fff7fff7fffafffdfffefffefffefffeffffff0200;
    decBuf[5226] = 256'h0500050006000500050005000a000c000c000b000d0013001300120013001200;
    decBuf[5227] = 256'h0f00120013001200140019001a0019001b001e001f0020001f00200022002500;
    decBuf[5228] = 256'h2200230022002500220025002800280029002e0030002c002b002c002d002e00;
    decBuf[5229] = 256'h3200330034003600340033003400310034003800390036003700380037003600;
    decBuf[5230] = 256'h37003a003b003c003e003d003d003d003e003d003e00430042003f0040003f00;
    decBuf[5231] = 256'h400041003e004100440046004700480047004a004b0048004500460045004a00;
    decBuf[5232] = 256'h4900440044004400440044004b004d004c004b004b004b004c004f004c004b00;
    decBuf[5233] = 256'h4c004b004c004d004e004d004b004b004c004b004c004a0049004a004c004b00;
    decBuf[5234] = 256'h4c004b0049004a004b004b004b004a0049004600440044004500460047004a00;
    decBuf[5235] = 256'h4900460045004400420041004200410042003f0040004100420041003e003c00;
    decBuf[5236] = 256'h3d003c003b003a00370038003700360036003600360033003200350032002e00;
    decBuf[5237] = 256'h2d002f002f002a002b0028002800280029002800280025002200250026002100;
    decBuf[5238] = 256'h1f00200021002000210020001a00170018001500140013001300120013001300;
    decBuf[5239] = 256'h140012000f0010000d0010000f000c000c000c000800050005000000fefffeff;
    decBuf[5240] = 256'hfafff7fffcfff9fff7fff7fff7fff7fff7fff2fff3fff6fff1ffefffeeffedff;
    decBuf[5241] = 256'hecffe9ffe3ffe2ffe3ffe1ffdeffdbffd9ffd6ffd5ffd4ffd2ffcdffd0ffd3ff;
    decBuf[5242] = 256'hd2ffcfffcdffcaffc7ffc6ffc4ffc1ffc0ffbaffb6ffb7ffb6ffb0ffadffaeff;
    decBuf[5243] = 256'hadffaaffaaffa5ffa4ffa5ffa4ffa2ffa1ffa2ff9fff9eff9aff94ff91ff90ff;
    decBuf[5244] = 256'h91ff92ff8fff8dff8aff87ff87ff82ff81ff80ff80ff7dff7cff7dff7aff79ff;
    decBuf[5245] = 256'h79ff79ff7aff76ff73ff74ff72ff6fff70ff6bff69ff6bff6bff6aff6bff68ff;
    decBuf[5246] = 256'h65ff64ff64ff64ff67ff6aff69ff64ff65ff64ff64ff5fff5dff5cff5dff5cff;
    decBuf[5247] = 256'h5bff5aff5dff5dff5dff5cff5dff5dff5eff61ff62ff5fff5eff5fff5eff5dff;
    decBuf[5248] = 256'h60ff5dff57ff58ff5dff5dff5eff5cff5bff5cff5eff5dff5dff5fff5eff5fff;
    decBuf[5249] = 256'h62ff61ff60ff61ff62ff5fff5eff5dff5dff5dff5eff5fff62ff61ff60ff61ff;
    decBuf[5250] = 256'h60ff63ff65ff63ff60ff63ff64ff64ff65ff66ff65ff63ff62ff64ff67ff64ff;
    decBuf[5251] = 256'h65ff68ff6cff6fff6eff6dff6eff6dff6cff71ff72ff6fff70ff74ff73ff76ff;
    decBuf[5252] = 256'h77ff74ff77ff7dff7eff7bff7cff7fff80ff82ff83ff86ff8aff8bff8aff8eff;
    decBuf[5253] = 256'h91ff8eff8fff94ff95ff94ff95ff95ff98ff9cffa1ffa3ffa8ffa9ffaaffaeff;
    decBuf[5254] = 256'hafffb0ffb1ffb5ffb9ffbaffbbffbcffbdffbeffc0ffc5ffc7ffcaffceffd3ff;
    decBuf[5255] = 256'hd5ffdaffdbffdbffdeffe1ffe2ffe6ffe7ffe4ffe9ffedffeeffeffff5fff7ff;
    decBuf[5256] = 256'hfafffdfffefffeffffff0400050007000a000e00110013001300150018001a00;
    decBuf[5257] = 256'h1b001c001d001e001f001e001f00210026002a002b002a002b002f0030003300;
    decBuf[5258] = 256'h36003600360035003400310036003a003700350037003d003e003d003d003d00;
    decBuf[5259] = 256'h400041003e003d003e003c003d00410044004300440044004500440044004300;
    decBuf[5260] = 256'h3e00410044003f003e0041003e0041004400430045004a004b00460045004300;
    decBuf[5261] = 256'h420041003e003d003e00410042003f003e003d003d003d004200440045004300;
    decBuf[5262] = 256'h40003f003e004100420043004400440045004800470044004500460044004300;
    decBuf[5263] = 256'h440041004000410040004400470048004b004d004e0051004e004a004c004f00;
    decBuf[5264] = 256'h4c004d004c004d00500051005000510052005100520052005300540057005400;
    decBuf[5265] = 256'h5300540055005600570058005700580057005400530052005200560055005200;
    decBuf[5266] = 256'h530052005300560057005900590058005700580053004f004c004b004c005100;
    decBuf[5267] = 256'h4e004f004e004a0049004a00470044004400430044003f003b0038003b003a00;
    decBuf[5268] = 256'h3b00380036003a0039003600340031002f002f002d002700240021001d001a00;
    decBuf[5269] = 256'h1a0019001a001a001b001a001a00150011000c00060005000800050003000400;
    decBuf[5270] = 256'h03000000fffffdfffcfffdfffcfffdfffcfff7fff5fff0ffecffedffecffebff;
    decBuf[5271] = 256'heaffe9ffe7ffe4ffe5ffe8ffeaffebffe9ffe9ffe7ffe2ffe2ffddffd5ffd6ff;
    decBuf[5272] = 256'hd7ffdaffddffdfffddffdcffdeffdeffddffdcffd7ffd8ffdbffd8ffd6ffd5ff;
    decBuf[5273] = 256'hd2ffd1ffd7ffdcffd9ffd7ffd6ffd5ffd4ffd5ffd4ffd5ffd6ffd5ffd6ffd3ff;
    decBuf[5274] = 256'hcfffceffd0ffd3ffd4ffd3ffd4ffd7ffd6ffd3ffd2ffd3ffd0ffd0ffd0ffceff;
    decBuf[5275] = 256'hcfffceffcfffd0ffcfffccffcdffceffcdffcaffc9ffc7ffc6ffc7ffc4ffc2ff;
    decBuf[5276] = 256'hc2ffc3ffc6ffc7ffc8ffc7ffc8ffc5ffc2ffc2ffc2ffc2ffc2ffc2ffc2ffc0ff;
    decBuf[5277] = 256'hbbffb9ffb4ffb2ffafffb2ffafffb2ffb4ffb5ffb8ffb5ffb4ffb5ffb4ffb4ff;
    decBuf[5278] = 256'hb4ffb4ffb1ffb0ffb1ffb0ffb1ffb2ffafffabffaaffa9ffa6ffa6ffa6ffa7ff;
    decBuf[5279] = 256'haaffabffaaffadffacffabffaaffabffa8ffabffacffabffaaffabffacffadff;
    decBuf[5280] = 256'hacffb0ffb3ffb2ffb1ffb4ffb3ffb4ffb3ffb2ffb3ffb2ffafffb2ffb1ffaeff;
    decBuf[5281] = 256'hb1ffb4ffb3ffb4ffb6ffb9ffbaffbcffbfffc0ffc2ffc2ffc2ffc3ffc2ffc3ff;
    decBuf[5282] = 256'hc9ffccffcbffcaffcdffccffc9ffc9ffc8ffc9ffc9ffceffd4ffd7ffd6ffd8ff;
    decBuf[5283] = 256'hdbffdcffddffdcffdbffdcffd9ffdaffdeffdeffdeffe5ffe7ffe8ffecffedff;
    decBuf[5284] = 256'he9ffeaffebffe8ffe9ffeaffebffedfff0ffeffff0fff1fff2fff3fff3fff4ff;
    decBuf[5285] = 256'hf3fff3fff3fff4fff5fff8fff9fff8fffafffdfffcfffbfffcfffdfffafffbff;
    decBuf[5286] = 256'hfefffffffcfffbfffcffffff0000fdff00000200070008000800080007000600;
    decBuf[5287] = 256'h0300020005000600080008000700080007000100000001000100060007000800;
    decBuf[5288] = 256'h0c0010001300160011001000130010000f000f000c000d000f00100015001b00;
    decBuf[5289] = 256'h1c001b001d001e001d0020001d001b001c001d001c001d001d001e001f002000;
    decBuf[5290] = 256'h23002200240029002b00300032003200340039003b003a003b003e003f003e00;
    decBuf[5291] = 256'h3b003a003d0040003f003e00420043004000410042004300470048004d005300;
    decBuf[5292] = 256'h5500560059005a005b005c005c005d0060005d005b005d006000630063006300;
    decBuf[5293] = 256'h630068006a006a006700660065006400650068006900680069006b006e007100;
    decBuf[5294] = 256'h710078007a007800770078007300720071006f00700071007100740077007600;
    decBuf[5295] = 256'h7700780077007600770074007300740075007400730072007500740071007100;
    decBuf[5296] = 256'h7300740071007100730072007500740071007100700071007000710070006d00;
    decBuf[5297] = 256'h6c006b006a006b006a006a0069006a0069006a006c006f006c006d0070007100;
    decBuf[5298] = 256'h70006d006900680069006600670064005e005d00600061006200630063006600;
    decBuf[5299] = 256'h67006600670066006700640065006600670068006a006a006900680065006300;
    decBuf[5300] = 256'h62005f005c005d006000610060005f005c005c005c005f0060005f005e005f00;
    decBuf[5301] = 256'h6300640060005f0060005d005c005d0060006100620064006700660065006400;
    decBuf[5302] = 256'h63005d005b00560054004f004d004e004e004f00520056005b005c005e006100;
    decBuf[5303] = 256'h62005f005c005c005900550050004e004d004c0049004a0049004a004d004c00;
    decBuf[5304] = 256'h4d004f005400510050004e004900470042004000400040003f003c003d003e00;
    decBuf[5305] = 256'h3900390038003300340039003800370039003900320030002d0029002a002900;
    decBuf[5306] = 256'h2a002b002d002e002f002c00260022001d001d001c00170018001b001a001b00;
    decBuf[5307] = 256'h1a001700150010000c0008000700040003000600070006000300060007000800;
    decBuf[5308] = 256'h07000600070004000100fffffafffafffafff8fff5fff6fff3fff1fff2ffefff;
    decBuf[5309] = 256'he9ffe6ffe5ffe5ffe5ffe8ffe9ffecffecffecffecffecffe9ffe6ffe0ffdfff;
    decBuf[5310] = 256'hdeffdcffd9ffdaffd7ffd8ffdbffd8ffd9ffdcffddffdcffddffd8ffd4ffd1ff;
    decBuf[5311] = 256'hcdffcaffc9ffcaffcdffceffcfffd1ffd4ffd3ffd0ffd0ffcbffc9ffc8ffc7ff;
    decBuf[5312] = 256'hc8ffc7ffc8ffc5ffc6ffc3ffc1ffc0ffc1ffc0ffc1ffc3ffc4ffc3ffc1ffc0ff;
    decBuf[5313] = 256'hbbffb9ffb6ffb5ffb4ffb7ffb8ffb9ffbbffc0ffbbffbbffbbffb9ffb6ffb5ff;
    decBuf[5314] = 256'hb3ffaeffadffadffaaffa7ffa8ffabffacffaeffb3ffb4ffb3ffb4ffb3ffaeff;
    decBuf[5315] = 256'hb1ffadffaaffabffacffa9ffaaffabffa6ffa4ffa1ffa0ff9eff9dff9aff99ff;
    decBuf[5316] = 256'h98ff99ff98ff99ff9effa0ffa3ffa6ffa6ffa7ffa6ffa4ffa1ffa0ff9eff99ff;
    decBuf[5317] = 256'h98ff99ff9aff9bff9eff9fff9eff98ff95ff92ff91ff8fff8eff8fff91ff94ff;
    decBuf[5318] = 256'h97ff98ff95ff96ff93ff92ff97ff98ff98ff9fffa1ffa0ffa1ffa0ff9eff9bff;
    decBuf[5319] = 256'h9aff98ff97ff99ff9eff9fff9eff9fff9eff9bff98ff96ff93ff94ff95ff92ff;
    decBuf[5320] = 256'h97ff9bff9effa4ffaaffaeffb4ffb9ffbbffbeffbfffbcffb6ffaeffabffa6ff;
    decBuf[5321] = 256'ha3ffa2ffa5ffabffb0ffb6ffbeffc3ffc6ffc9ffcaffc9ffc6ffc2ffbfffc0ff;
    decBuf[5322] = 256'hc1ffc2ffc4ffcbffcfffd3ffd9ffdeffdfffe0ffdfffdcffd6ffd2ffcdffcbff;
    decBuf[5323] = 256'hc6ffc9ffcfffd7ffdfffe4ffe6ffecfff1fff2fff3fff2fff1ffeeffefffecff;
    decBuf[5324] = 256'heaffe7ffe6ffe5ffe8ffecfff1fff7fffafffcfffbfff9fff3ffebffe5ffe0ff;
    decBuf[5325] = 256'hddffdeffe4ffecfff6ff000006000c00110012000d0007000100f9fff6fff3ff;
    decBuf[5326] = 256'hf2fff3fff6fffaff020005000600070006000200fcfff7fff3fff0ffeffff2ff;
    decBuf[5327] = 256'hf5fffdff020009000f00150018001b001d001c00180014000f00090007000200;
    decBuf[5328] = 256'hfefffbfffeff000007000e00190022002b002e002f002d0025001d0014000e00;
    decBuf[5329] = 256'h08000b000e0014001c0024002b003100350036003500320030002f002e002f00;
    decBuf[5330] = 256'h33003900410047004a004b0046003f0037002e0025001d001a001e0025003000;
    decBuf[5331] = 256'h3f00510061006c007200740072006d00640059004b0042003a00360034003600;
    decBuf[5332] = 256'h39003c0044004e00550060006b0071007a0080007f007e007b00720068005d00;
    decBuf[5333] = 256'h55004e004b0047004a00520058005d0061006400650064005f005f005f006400;
    decBuf[5334] = 256'h6a0072007c0088009000920093008d0083007400660053004000390033003900;
    decBuf[5335] = 256'h480057006d00810094009b009d00930083007400620057005400520054005c00;
    decBuf[5336] = 256'h61006a00730074007500730070006d006d006a006d006f007200730072006d00;
    decBuf[5337] = 256'h6900610059005200510054005c0064006d0076007900780074006d0067005f00;
    decBuf[5338] = 256'h580055005400550055005c006200660069006a0065005d0055004c0046004700;
    decBuf[5339] = 256'h4e005b006900790084008a0085007600600040002b0018000600090012002400;
    decBuf[5340] = 256'h3e005e0073008e0099009c0093008600710051003c00210016000d000a000d00;
    decBuf[5341] = 256'h14001e0028003100390041004a00510059005c005c0058004e00420037002c00;
    decBuf[5342] = 256'h2000180016001500110010000f000b0006000200fcfff4ffeeffebfff1fffbff;
    decBuf[5343] = 256'h0a002400440059006c007000600046002000f2ffb9ff94ff71ff6bff71ff80ff;
    decBuf[5344] = 256'ha1ffc7ffebff0b0020002c002f0020000c00f9ffdfffceffbeffbbffb9ffc0ff;
    decBuf[5345] = 256'hc2ffc0ffbbffafffa2ff92ff83ff7dff7fff87ff94ffa8ffb5ffc5ffd0ffd2ff;
    decBuf[5346] = 256'hcdffc5ffbaffabff9dff8dff83ff7dff74ff6fff6eff6cff66ff65ff62ff61ff;
    decBuf[5347] = 256'h65ff71ff83ff93ffabffbaffc3ffc0ffb0ff94ff71ff47ff2bff12ff0dff11ff;
    decBuf[5348] = 256'h1dff3cff5aff7dff94ffa1ffa5ff9aff84ff65ff3fff25ff0eff0aff0dff1fff;
    decBuf[5349] = 256'h3bff5eff75ff82ff86ff74ff65ff4bff32ff1cff0eff0bff0eff14ff1eff2aff;
    decBuf[5350] = 256'h36ff3dff3cff38ff30ff29ff27ff26ff2aff34ff3dff46ff4eff4bff40ff31ff;
    decBuf[5351] = 256'h1bff07fff4fee4feddfedffee8fef4fe04ff0fff19ff1eff20ff1eff1dff1bff;
    decBuf[5352] = 256'h1dff22ff2fff39ff45ff50ff52ff4bff38ff1bfff8fecffeb3fe99fe94fe99fe;
    decBuf[5353] = 256'hacfed3fef6fe20ff3cff4cff50ff4cff48ff37ff2dff30ff33ff3fff49ff4fff;
    decBuf[5354] = 256'h4dff3cff18fff4fec1fe91fe72fe6cfe71fe9bfecefe19ff5fff9fffc8ffdfff;
    decBuf[5355] = 256'hd8ffb9ff91ff63ff2bff05ffe3fed0fecbfed0fed4fed9fee4fef6fe05ff14ff;
    decBuf[5356] = 256'h2bff41ff5bff7bff90ffa3ffaeffb1ff9dff85ff63ff39ff12fff8feeafeeffe;
    decBuf[5357] = 256'hfafe13ff35ff4cff6aff76ff80ff7dff6fff67ff64ff62ff6cff7fff97ffadff;
    decBuf[5358] = 256'hbbffc3ffc1ffaeff91ff6eff4eff30ff1cff12ff15ff2fff4eff75ff99ffc2ff;
    decBuf[5359] = 256'hdefff8ff06000a00feffedffd7ffb7ffa2ff8fff7dff7aff7dff8aff9bffaeff;
    decBuf[5360] = 256'hc0ffd1ffdcffe2ffe0ffdeffd7ffd0ffcaffc4ffc3ffc6ffccffd9ffebff0000;
    decBuf[5361] = 256'h20003e00590071007b007d006b0047001900e1ffbcff8bff79ff73ff8dffc0ff;
    decBuf[5362] = 256'hfdff37006c009c00bb00b500a6007c0055003b002400200033005a008800c000;
    decBuf[5363] = 256'he600ed00e600ca0088004800feffb8ff9cff94ffaaffdbff2c008f00ec002901;
    decBuf[5364] = 256'h760194018b0183015d011f01e600b100810055002e001400fdff010005001e00;
    decBuf[5365] = 256'h40007300b100fb0041018101aa01d001d701c401910153010901af0072003b00;
    decBuf[5366] = 256'h1d0014002d0053008300bb00ef0020013f015001550150014c0150015a016401;
    decBuf[5367] = 256'h72018401870180016a0145011701df00aa0088006900630072009300c100fa00;
    decBuf[5368] = 256'h3d016b019401ba01ce01e101db01d601bf01aa018701670138010c01d900a900;
    decBuf[5369] = 256'h8a0079007e009f00cd0012015201ad01e9010a0228021f020702d20194015a01;
    decBuf[5370] = 256'h2601f600d700d100d600e400f90014012d0149015c0175018b019901ab01b701;
    decBuf[5371] = 256'hc201c001b701a5018601690146012501100105010801180132014a0160016e01;
    decBuf[5372] = 256'h7b01790173016501550146013c0133012e013601400150016301750186019501;
    decBuf[5373] = 256'h9f01a1019c01910182016c0152013a011e010201e300ce00c200bf00c200ca00;
    decBuf[5374] = 256'hdd00f200060123013e015e017b019701af01bf01c701bf01aa0190016a013c01;
    decBuf[5375] = 256'h1001dd00ad0081004f002c000d0007000d0024004a008200d50022017c01d101;
    decBuf[5376] = 256'h08023a0231021802d4017001f80086001f00dcff9fff7eff88ffb6ff00004600;
    decBuf[5377] = 256'h9800cf0001012f0137012f0129010901ed00c900b20094007900610051003d00;
    decBuf[5378] = 256'h2b001f0014000a000c0014002800440067009100b800dc00f30000010401f200;
    decBuf[5379] = 256'hd600ac006e002400deff8bff3efff8feddfed5feebfe29ff84fff1ff7600f300;
    decBuf[5380] = 256'h4401ab01d401e001a9016301ec007a00d8ff6cff0affb0fe80fe8efeb7fedbfe;
    decBuf[5381] = 256'h28ff6effaefff8ff160031004a0043002e00280017001c002a003f005a006c00;
    decBuf[5382] = 256'h75006d0050001d00dfff95ff4fff0fffd6febffec6fed9fe0bff3bff74ffa8ff;
    decBuf[5383] = 256'hcbffddffd8ffbeffa7ff81ff67ff50ff54ff6fff96ffceff120052006a008100;
    decBuf[5384] = 256'h7a004e000500abff56fff3fe96fe41fe0afe00fe09fe32fe85fed2fe2cff80ff;
    decBuf[5385] = 256'hcdffffff1b0023001c000700e8ffc0ff9cff85ff70ff64ff61ff6aff73ff76ff;
    decBuf[5386] = 256'h73ff60ff43ff11ffe1fea8fe74fe52fe4bfe51fe75fe9efedcfe27ff6dffacff;
    decBuf[5387] = 256'he6ff0c0020000e00e6ffaeff6aff2aff01ffebfee4fe03ff36ff74ffbefff0ff;
    decBuf[5388] = 256'h0b001300eeffb0ff45ffc0fe43fed1fd6afd42fd36fd6dfdc7fd64fefcfed4ff;
    decBuf[5389] = 256'h63001a016101a2018f015901e7006300c2fffffe7cfe06fec5fdb1fdc3fdf4fd;
    decBuf[5390] = 256'h3efe9bfef0fe3dff6fff78ff80ff6aff48ff28ff17ff08ff03ff10ff24ff51ff;
    decBuf[5391] = 256'h89ffbeffeeff26003d0044003d002100f3ffbbff77ff37fffefed8fea8fe89fe;
    decBuf[5392] = 256'h78fe73fe77fe84fe98feb0fec6fed4fee7fefcfe10ff2dff50ff7affb7fff1ff;
    decBuf[5393] = 256'h260064009d00c300e500eb00db00ac005b00f8ff65ffdcfe3bfea3fd41fdc4fc;
    decBuf[5394] = 256'h93fc85fcc8fc1cfdc1fd68fe56ff3300fc00b30159029a02ae027802e6013501;
    decBuf[5395] = 256'h600096ffdffe0afe7afd60fd48fd5efd99fd16fe87feeffe4cff89ffaaffa0ff;
    decBuf[5396] = 256'h72ff39ff13fff1fef7fe2aff83fff0ff750016018201e401f601c50140019f00;
    decBuf[5397] = 256'hddfff2fe14fe85fd02fdbbfcfcfc36fdd7fd9afe51fff7ff6300c500d700a600;
    decBuf[5398] = 256'h5d00ffff92ff48ff05fff9fe1aff60ffd7ff6900cb0048019a018b016301f600;
    decBuf[5399] = 256'h7100acfff5fe4ffeb8fd56fd44fd74fdbefd51fedbfe7cff13007500ab00bb00;
    decBuf[5400] = 256'hac00840047001000deffd5ffdefff4ff32006c00af00ef0018012f011a01e200;
    decBuf[5401] = 256'h8f001600a5ff20ff7ffe13feb1fd57fd47fd56fd7efdebfd70fe11ffd3ffbf00;
    decBuf[5402] = 256'h5d012602a9021f033503fa02a1020e0237016d0082ffe4fe1bfeccfd85fd9bfd;
    decBuf[5403] = 256'haefd08fe7afee1fe59ffaafff4ff02000e000300e5ffdcffe4ff09005500c300;
    decBuf[5404] = 256'h4801c5011602600288024b02d20120014a0047ff53fe76fdacfc5efc46fcb2fc;
    decBuf[5405] = 256'h3cfd24fe41ff4d004101e0016f02be02760236028501df001c0065ffeefed9fe;
    decBuf[5406] = 256'hecfe46ffb8ff5a00f1005301ad019c015301a500cfffccfed8fd3afdaafc5cfc;
    decBuf[5407] = 256'h74fc0bfd0afe44ff6b00c401ac027f03f203cf037003a702bc019f0093ff9efe;
    decBuf[5408] = 256'h00feaafdc4fd0bfea3fe2cffcdff6400c700d800c8006100ceff1dff77fe0bfe;
    decBuf[5409] = 256'ha9fdbbfd0cfeaefe71ff5c00780138022c038b03a8035a03b302c601a9009cff;
    decBuf[5410] = 256'h62fe90fd1dfdfafc19fda9fd60fe65ff5900f8004e019c015501e900380092ff;
    decBuf[5411] = 256'hcffe4dfe35fe4bfeadfe4eff1000fb00d9016802eb020303ed026402c3010001;
    decBuf[5412] = 256'h150038ffa8fef1fdaafd69fd7dfdd6fd48feeafe81ff3200a900150150016201;
    decBuf[5413] = 256'h3101e700a4004f000200e4ffdbff050048009a00fd0040017d0188015601f100;
    decBuf[5414] = 256'h7900c6ff20ff89fefffda6fdb6fde2fd40fedefe75ff2600cc006301ed014602;
    decBuf[5415] = 256'h7702a302960259020c028a01e900260070ffc9fe07fe84fd3dfd27fd62fd03fe;
    decBuf[5416] = 256'hc6fe7cff8200760114026a0250023802a10118015300d0ff89ff73ff87ff0400;
    decBuf[5417] = 256'hb7005d01f5012f024102f0014e01600043ffeafd02fd2ffc09fc2cfccafc06fe;
    decBuf[5418] = 256'h81ffe6008802a0039f04ce04a404e403aa022f01caff28fe10fd77fc48fcc7fc;
    decBuf[5419] = 256'h87fdc1fe3c00a101e502b8032b040804a903a7026d01f2ff8dfe48fd75fc02fc;
    decBuf[5420] = 256'h25fcc3fcfffd7bffe00081029a03cd03fb037d0370023601bbffbcfed4fd56fd;
    decBuf[5421] = 256'h7cfde5fd01ff5b009f011a031904a504cf040f04d5025a018fffdffde5fb19fb;
    decBuf[5422] = 256'h60fa98fa31fb76fc45fef6ffef01cb03ff04a8057505ea041704be021c0193ff;
    decBuf[5423] = 256'h2efe47fdc8fca2fc50fdeefd2bff51005e015202f002d402850280018c0030ff;
    decBuf[5424] = 256'h48fe75fd02fd6bfd09fe0cff4600c101c002a803d2035f03f602d90180003bff;
    decBuf[5425] = 256'h69fe5cfdf4fcd4fc2afdadfdb2fea6ffc300cf017e02dd023303190301039502;
    decBuf[5426] = 256'he4013e01a700f6ff50ffb8fe2ffef9fdc9fdd7fd00fe6dfef1fe6fff21009800;
    decBuf[5427] = 256'h04016601780168013c011401bf009e00800077008f00a600d600f50011010c01;
    decBuf[5428] = 256'hec00ac005a00f7ff7fff0dffa6fe63fe3efe49fe7bfecdfe46fff9ff9f006201;
    decBuf[5429] = 256'he5015b02c802b4027e02ec0114014b002cff6cfe78fdd9fc83fc9dfc44fd06fe;
    decBuf[5430] = 256'h5aff9e001a027f036604e504be0456043903e0013e00b6feb7fdcffc50fc2afc;
    decBuf[5431] = 256'hd8fcb6fdb8feadffc9008901f201d2017c01c5001f0087fffefec8feb8fe1fff;
    decBuf[5432] = 256'h98ff4a002001b0016702ae02c40289022f027d01d600e9ff0bff7bfec5fd7dfd;
    decBuf[5433] = 256'h68fd7bfdf8fd8bfe3bff1100da005d01d401e901d6015901c60016009fff08ff;
    decBuf[5434] = 256'hcdfebbfeecfe70ffedffa00017018301970185015401ed005a00f8ff7aff4aff;
    decBuf[5435] = 256'h1dff2bff80ffcdff3b00a200e500f100d0008a002600adff1bffb9fe83fe52fe;
    decBuf[5436] = 256'h61fe89fedefe2bff85fff2ff5a00d2004401ab0109024502660270024302f801;
    decBuf[5437] = 256'h7601d50013005cffb6fe1efe95fd5ffd70fd9cfd14fea6fe30ffd1ff6800f100;
    decBuf[5438] = 256'h4b017c018a017d0159010c01c60061001e00c9ff7cff4aff1dff25ff3cff6cff;
    decBuf[5439] = 256'hbdff0a006400a100d800f600ec00c30080004000f6ffb0ff82ff7aff90ffb3ff;
    decBuf[5440] = 256'hebff1f00420048002c00f3ffb0ff5eff11ffdffec3febbfed2fef4fe2cff7fff;
    decBuf[5441] = 256'he2ff3f00c50042019301dd01ea01de01a7014d01e00079001b00c6ff79ff33ff;
    decBuf[5442] = 256'h06ffdcfec6fecdfee0fe12ff42ff6eff95ffafffb4ff9eff7cff49ff26ff07ff;
    decBuf[5443] = 256'h0dff45ff98ff2700d7007d014002c30239032403e902240239011d0010ff1cfe;
    decBuf[5444] = 256'h3efde8fccefc45fd07fef3fe0f001c01ca01680285026b02c501d700f9fff7fe;
    decBuf[5445] = 256'h03fea4fd4dfd68fddefd76fe26fffcff8c004301e9015502b702ed02dd02b002;
    decBuf[5446] = 256'h53029d01e600100047ff90fe49fe08fe1cfe51fec3fe0dff6affa7ffdeffe8ff;
    decBuf[5447] = 256'hdfffc6ffb0ff7fff6dff72ffa0fff2ff6b00fd00860103025502810259020402;
    decBuf[5448] = 256'h5f018900c0ffd5fef7fd68fd4efd65fdfdfdd5fed7ff1101e401a40252033203;
    decBuf[5449] = 256'hdc02250250014d0013ff40fe80fdd2fcb2fc96fce4fc8afd4dfe38ff55006101;
    decBuf[5450] = 256'h550233038903a3035c03f0023f0269016700b8ffdbfe85fe36fe1ffe5ffec2fe;
    decBuf[5451] = 256'h62fffaffaa00210137012301ca00380087ffe1fe49fee7fdb2fdc2fd0cfeb9fe;
    decBuf[5452] = 256'h8fff9200860163022d037b03630322034b024801540037ff2afe7cfd1dfd00fd;
    decBuf[5453] = 256'h83fd29fe17ff340040017a02f9026c034903ab026f01f3ff8efe4afd23fc63fb;
    decBuf[5454] = 256'h86fbe5fbaefc02fea3ff2c01910279034b042504bc03df02a3017c0023ff3bfe;
    decBuf[5455] = 256'h68fd42fdaafd88fe8aff7f005c01250274022c029501bd0081ff5afe4dfd59fc;
    decBuf[5456] = 256'hfafbdefb2cfc31fd6bfee6ff4b01ed0205049e047004f1033203f8017d0018ff;
    decBuf[5457] = 256'h76fd5efcc5fb96fbc0fbcdfc07fe82ff4d0182029a033304050487037a024001;
    decBuf[5458] = 256'hc5ffc6fe81fd03fdddfcfffc5efdeefdd9fe77ff070055006d002c00f1ff74ff;
    decBuf[5459] = 256'h23fff7fee9fe3effb7ff6a00400109028c02020343033003d60224021e012a00;
    decBuf[5460] = 256'h0effb4fdccfcfafb87fb64fb83fb13fccafccffd09ff30003d013102cf025f03;
    decBuf[5461] = 256'had036603fa022202e500bfffb2fe78fdfafc87fceffc4efd17fe37ff43003701;
    decBuf[5462] = 256'hd6016502b4026c02000228015f0040ff80fed2fd73fd1cfd37fd7efdeafd4cfe;
    decBuf[5463] = 256'ha5fef7fe5effd6ff28008f00ec0029014a0168015f013601f200a0002700b5ff;
    decBuf[5464] = 256'h4efff0feb4fe93feb1fef1fe3bff81ffc1ffdaffd2ffb0ff77ff34ff06fffefe;
    decBuf[5465] = 256'h06ff36ff93fff1ff46007d0087006c0011008bffebfe7efef5fdbffdaffdf9fd;
    decBuf[5466] = 256'h71fe24ff29001d01fb018b02d902c10255027d017a0041ff1afe5afdf1fcd2fc;
    decBuf[5467] = 256'heefca5fd7bfe44ff2f000d019c01b7019f01330182007dff43fe70fd64fcfbfb;
    decBuf[5468] = 256'h1bfc71fc5cfd79fed2ff73018c02f1037c04a60433043f0322027c00f3fef4fd;
    decBuf[5469] = 256'hb0fc86fc5ffcc8fc27fdf0fda7fe1eff8affc5ffb3ff82ff56ff2eff09ff14ff;
    decBuf[5470] = 256'h46ffabff3e00c7006801ff013a022802d70152018e00a3ffc5fe36feb3fdcbfd;
    decBuf[5471] = 256'h0cfe95fe36fff8ff7b00f2000701f4009a002900a4ff03ff6cfe0afed4fdc4fd;
    decBuf[5472] = 256'hf0fd83fe34ffdaff9d005301ca010b021f02e9017701f30052008fff0cff66fe;
    decBuf[5473] = 256'h25fe12fe47fe99fe1dff77ffe8ff15003d0061006c0076007f00880080006b00;
    decBuf[5474] = 256'h40002400f5ffe3ffc7ffc1ffaaff84ff56ff11ffd1fe98fe72fe87febffe2fff;
    decBuf[5475] = 256'hc2ff72004801d80126023e022802ed014d01b5002c008bff1fffe4fed2fec2fe;
    decBuf[5476] = 256'hd1fef9fe1dff54ff86ffb4ffedff220060008900af00c300c900b90095005900;
    decBuf[5477] = 256'h0e00b4ff78ff2bff21ff2aff64ffb6ff2f00a10008018001b101dd01d001c401;
    decBuf[5478] = 256'h77011d01b0002b00d2ff60ff16ffeefecafea9fe8bfe82fe79fe81feb1fe02ff;
    decBuf[5479] = 256'h7bff2e00d4006c011c029302d402c0028b02f8016f01ce003700adff54ff44ff;
    decBuf[5480] = 256'h52ff7bffcfff0600380042002900f4ffa9ff4fff12fff1fe0fff4fffcbff6c00;
    decBuf[5481] = 256'h2e01e5015c029d02890230029d01ed00170087ffd0fe89fe74feaefe2cffdeff;
    decBuf[5482] = 256'h85004701ca011102fb01c10120018800ffff82ff51ff60ffa3ff10007700ef00;
    decBuf[5483] = 256'h41016d017a0156011f01c5004000c2ff71ff27fffffe0bff42ffb0ff18009000;
    decBuf[5484] = 256'h22018401de012f023e024b022702da016c01ca003200a9ff4fffdefeb1fea4fe;
    decBuf[5485] = 256'he1fe2eff9cff3e00d5005f01dc012d021e02db015601b5001e0094ff3bff0aff;
    decBuf[5486] = 256'h19ff77fffcff9d0034019601f001e001b301560101019e005b0037001600f8ff;
    decBuf[5487] = 256'hdcffc3ff9eff97ff9dffb9ffe8ff2c006c00a600cb00e000e600e100d100c300;
    decBuf[5488] = 256'hae00a3009f00a800bd00d900f500f800e200b7005900c6ff3dffc0fe6efe60fe;
    decBuf[5489] = 256'ha3fe10ffb2ff750060013d02cd024f03670326037602a0019d0063ff91fed1fd;
    decBuf[5490] = 256'h68fd49fd65fdb4fd5afef1fea2ff4800b4003e017301c501f10119023d024802;
    decBuf[5491] = 256'h3e02fe01b4013201b500230099ff40ff0fffc6fe9dfe79fe58fe4efe45fe5efe;
    decBuf[5492] = 256'ha1fef3fe6cffdeff6300e0005201b901170253025e0254021402a90107014400;
    decBuf[5493] = 256'h8dffe7fe50fe15fedffd10fe5afeb7fe3dffbaff2c009300d600fa00ef00e500;
    decBuf[5494] = 256'hca00b100b800b200b800a7006f000d007afff1fe50fee4fda9fdbbfd2cfeecfe;
    decBuf[5495] = 256'hd7ffb5007e0135027c0292025702da0127018100beff3bffc5fe84fe49fe5bfe;
    decBuf[5496] = 256'h6bfe97febffefcfe33ff51ff48ff2fff19ff1fff58ffb9ff4c00fd00a3013b02;
    decBuf[5497] = 256'h7502640212027001ad00c2ffe5fe1cfe99fd22fd0dfd20fd7afdebfd70feedfe;
    decBuf[5498] = 256'h80ffe2ff5f00d10038019501ea010b02ed018901f60045006fffa6fe24fedcfd;
    decBuf[5499] = 256'hc7fd02fe37fe88fef0fe18ff3cff47ff3dff34ff0bfff4feedfe00ff33ff9aff;
    decBuf[5500] = 256'h3c00ff00ea0188025103a003b7032003fa017f00b4fe03fd7afb15fa8af9b4f9;
    decBuf[5501] = 256'h74fa68fb04fd8cfef1ff36015d021d038503a503c2037303fd023a024f017200;
    decBuf[5502] = 256'ha8ffbdfe1ffe8ffd0dfdc5fcdbfc16fd6ffd02fe8bfe08ff7affe1ff24006100;
    decBuf[5503] = 256'h9800ca00d300ca00a50067000c00b7ff6aff4cff56ff7fffc2fff0fff8ffe2ff;
    decBuf[5504] = 256'hb2ff60ff13ffe1feeafe14ff57ffbcff19006e0079005b001b00b0ff49ffebfe;
    decBuf[5505] = 256'haefea3fe99feb5fedefe13ff50ffabff18009d001a018c01d601c8018c011301;
    decBuf[5506] = 256'h3f0076ff8bfeaefde4fc96fcaefc1afdcbfdd0fe0a00dc00e901520271025402;
    decBuf[5507] = 256'hd2012c01bf005d000400d3ffc4ff82ff45ffe2fe6afef8fd91fd68fd5cfd7dfd;
    decBuf[5508] = 256'hd7fd5dfefefeebffc90092017d02dc023203e4023e025001330027ff32fe13fe;
    decBuf[5509] = 256'hf6fdadfe53ff4100df006f015501de001b00fcfeeffd41fda3fcc0fc0efde4fd;
    decBuf[5510] = 256'he7fe200047015402bd02dc02bf023d0267019e00b3ff15ff85fe6bfe53fe94fe;
    decBuf[5511] = 256'h1dff9aff4d002301b3016902b1027002e601da0081ffe0fdc7fcc8fb3dfb67fb;
    decBuf[5512] = 256'h27fc1bfd77fe1800310196027e03fc036f0492047204e303f8029c01570030ff;
    decBuf[5513] = 256'h24fe75fdd7fcbafcd4fc1cfd88fd11feb2fe1effa8ff25007600dd0020017501;
    decBuf[5514] = 256'hc2011c027102a802c602cf029502250272019c00d3ff1cff46feb7fd68fd50fd;
    decBuf[5515] = 256'h3bfd76fdf3fd85fe36ff0b00d5008c01020243023002fa01a901410119013e01;
    decBuf[5516] = 256'h7501cf012402450213028a01b200afffbbfe1dfe8dfd3ffd56fd6cfda7fd00fe;
    decBuf[5517] = 256'h72fef7fe74ff2700fc00c6014802ef025b039603a70397034d03f00252029001;
    decBuf[5518] = 256'ha40088ffc8fed4fd75fd1ffd39fd51fdbdfd1ffe9cfe4ffff5ff8c0016019301;
    decBuf[5519] = 256'h050231022302ff01c801820154011b01f500c5009900670037000b00effff4ff;
    decBuf[5520] = 256'h1d005b00a600d800f300b9005800c5ff3bff9afe59fe1ffe30fe82fecbfe29ff;
    decBuf[5521] = 256'h96fffdff91004101e701aa026103d803ed03b20312034f02640147003bff8cfe;
    decBuf[5522] = 256'haffd59fd0afd22fd63fdecfd8dfe50ff0700ad00ee000101ef00df00b300c000;
    decBuf[5523] = 256'he5001c016201b401eb011d023802510249022702c90136015e005cff22fe4ffd;
    decBuf[5524] = 256'h42fcdafbf9fb50fc07fddcfda6fec5ffd20080015d022703a903200461044d04;
    decBuf[5525] = 256'hf40362038a02c001d500f8fff5fe47fe69fda0fc1efcd6fbc1fbfcfb9cfcb6fd;
    decBuf[5526] = 256'h0fff54007a01d4025f03dd030404e1038203f20207022a01270033ff95fe05fe;
    decBuf[5527] = 256'hb7fdcefd3afe9dfe3dffd5ff5e00b8000901350142011e01d1004f00aeff17ff;
    decBuf[5528] = 256'h66fe1ffe35fe6ffe10ffd3ff8a0001016d01cf0104021502410234022702f001;
    decBuf[5529] = 256'h6e01ce00e0ff02ff39fe82fd0bfdf6fc09fd3ffdd1fd5bfe1fffd6ff7c003f01;
    decBuf[5530] = 256'hf6016d02d90214030203d1024c028801d100fbff32ff7bfed5fd69fd06fdf5fc;
    decBuf[5531] = 256'h25fdaafd6ffe5aff37003a01e801470264024a02d3013c018b00e5ff22ff6bfe;
    decBuf[5532] = 256'hf5fdb4fdc7fd44fe18ff1a000f01ec01b5020403bc025002a001ca00010015ff;
    decBuf[5533] = 256'h38fe6ffdecfc75fc35fc6ffc10fdfefd1bff74005c018302f6025f033f03e902;
    decBuf[5534] = 256'h6602c0012901780001006aff08ff8bfe39fe0dfecafdbefdb3fdd1fdfffd6afe;
    decBuf[5535] = 256'heffe90ff5200d5007b01bc01d0019a012801c100630027000600100019002100;
    decBuf[5536] = 256'h0b00bfff65fff8fe91fe68fe75fec2fe30ffb4ff3100a300cf00c2009e003b00;
    decBuf[5537] = 256'hddff70ff09ffabfe6efe79febffe48fff9ffcf005e01e101f9018d0103016200;
    decBuf[5538] = 256'ha0ffe9fea2fe61fe74fecefe1fff69ffc6ffebfff6ffd8ffaaff70ff3cff27ff;
    decBuf[5539] = 256'h47ff9bff2000c1002d018f01c5017401ef002a003fffa1fe11fef7fd0ffe50fe;
    decBuf[5540] = 256'hb2fe2fffa1ff26007f00b000fa000701fb00c4006a00fdff5affeefe65fe2ffe;
    decBuf[5541] = 256'h1ffe86fe19ffcaffa0006901b701ff0193010901450059ff7cfeecfd9efdb6fd;
    decBuf[5542] = 256'hf7fda7fe4dff3b00d9006901b80170012f017f00d9ff6cff0affd5fee5fef4fe;
    decBuf[5543] = 256'h37ff8bffc2ffe0fffcff0400fdffdaffc7ffb7ffb1ffdbff19007400c9000001;
    decBuf[5544] = 256'h0a01b7003e008cffb6fe26fed8fdc0fd01fe8afe4fff3a001701a701f6010d02;
    decBuf[5545] = 256'hcc014301a200e0ff5dffb7fe76fe3bfe4dfe7efeaafeedfe42ffa5ff02005700;
    decBuf[5546] = 256'ha400ea0005010e01f700d5009d0059001900f0ffbbff8bff6cff50ff36ff0dff;
    decBuf[5547] = 256'hf1fecdfeb6feb1fed4fe1aff88ff2a00c1007201e90129021602bc012a017a00;
    decBuf[5548] = 256'ha4ffdbfe58fee1fda0fdb4fd0dfe7ffe04ffc8ff4b00f1005d01c001d101e201;
    decBuf[5549] = 256'hb501730105018100e0ff48ffbffe42fe11fe02fe10fe4cfeaffe28ffbaff4300;
    decBuf[5550] = 256'h9d000f0176019e01c201a1016f011d01a4003200aeff31ffbffe75fe4dfe41fe;
    decBuf[5551] = 256'h4cfe92fef6fe89ff1300b4004b01d4010a021a020b02ae012801640079ff9bfe;
    decBuf[5552] = 256'hd2fd4ffd08fd1efd80fd45fe30ff4c0059014d02ac020203e8027102da012901;
    decBuf[5553] = 256'h8300c0ff3effc7fe5bfe20fe32fe42fe8cfecffe3cff86ffe3ff08003f007100;
    decBuf[5554] = 256'h8c00c600090149019301b101a8016f010d017a00c9ff23ff8cfe2afe18fe48fe;
    decBuf[5555] = 256'hb0fe5eff0400c60049019001a6016b01ca003300a9ff09ffc8feb4feeafe3bff;
    decBuf[5556] = 256'ha2ffe5ff3a008700b900e7001001440167016d0151010401a100290096ff34ff;
    decBuf[5557] = 256'hdbfeaafe9bfe8efeb2fee9fe2fff81ffe4ff4200af0016017401b101d201c801;
    decBuf[5558] = 256'hbf0195015201ed007500e3ff59ffb9fe4cfe12fe00fe51feb8fe4bfffcffa200;
    decBuf[5559] = 256'h3a019c01ae019d013601be004c00c7ff6eff3dff4cff8ffffcff9e003501bf01;
    decBuf[5560] = 256'hd101c0015901c600eeff25ffa2fe5bfe45fe59fed6fe48ffafff0d0062008300;
    decBuf[5561] = 256'h8d009600af00c500da00e000f100ec00de00c900b5009d008700670049003600;
    decBuf[5562] = 256'h1e000800eeffceffa0ff5bff09ffbcfe8afe6efe98feeafe8fff3500f800af01;
    decBuf[5563] = 256'h5502960282024d02ba0131019000f9ff97ff1affe9febdfecafed6fe0dff67ff;
    decBuf[5564] = 256'hbcff1f007d00ea0016013e014a012901f700a5004200e4ff5fffe2fe70fe44fe;
    decBuf[5565] = 256'h37fe8bfe1affcbffd0007f015c02ec023a032203b6022d028c019e00c1ffbefe;
    decBuf[5566] = 256'hcafd2cfdd6fcbbfc03fd9afd4bfe50ff4400e200ab012e0275028b0277021e02;
    decBuf[5567] = 256'hac010a017300e9ff90ff5fff6eff96ffebff220040003700ecff92ff3effdbfe;
    decBuf[5568] = 256'hb2febffef6fe64ffcbff4300b500ff00270133012801f600c8007e0038000a00;
    decBuf[5569] = 256'h0200fbff0f0022003e004e0049003c00290010000100feff00000300f8ffdaff;
    decBuf[5570] = 256'h9aff24ffb2fe68fe5bfe7ffee2fe90ff66002f01e6018c02240337034903f802;
    decBuf[5571] = 256'h7302af01c300a7ff9afe60fd8efccefbabfb8bfb1bfcd2fc07fe82ffe7008802;
    decBuf[5572] = 256'h110410059b05c505520518049d02d20022ff99fd34fca9fb2bfb9efb06fc23fd;
    decBuf[5573] = 256'h30fe69ff90009d014b02e9020603ec02a50239028801e2001f009dfff6fe8afe;
    decBuf[5574] = 256'h4ffe1afe2afe39fe7cfed0fe49ffdcff6500e20054018001a8019c0165011f01;
    decBuf[5575] = 256'hcd006a000c00b8ff55ff12ffbdfe70fe52fe5bfe74fec6fe29ffa2ff34009600;
    decBuf[5576] = 256'hef0041016d015f013b010401be007e0044001f000a0011000b00fcffc9ff7dff;
    decBuf[5577] = 256'h0fffa8fe2ffefffd0dfe50feeefe85ff5d00ed007001b701cc0192011401a300;
    decBuf[5578] = 256'h3b00deff89ff52ff48ff51ff7affbefffeff27004c0061004e002700e4ff92ff;
    decBuf[5579] = 256'h45fffffed2feb9fec0fee3fe34ff97ff0f00810006015f0190019f015c010701;
    decBuf[5580] = 256'h8e001c0097ff3effedfedefeb6fec2fecdfed7fef2fe1cff5fff9fffe9ff4300;
    decBuf[5581] = 256'h9800cf0001011d0135013d012801f0008e00160063ffbdfefafdacfd65fd7afd;
    decBuf[5582] = 256'hddfd7dfe40ff2b000901d201200267025202f0019601e4003d00a6ff1dff9ffe;
    decBuf[5583] = 256'h4efe3ffe32fe56fe8dfebffefffe39ff7dffbcfff6ff2b005b007a009600b000;
    decBuf[5584] = 256'hd000ff0037016c018e0194016201fb003b0050ff72fea9fd26fddffcf5fc57fd;
    decBuf[5585] = 256'hd4fda7fe71ff2700fd005301d601ee010302f001de018d014301cb003800afff;
    decBuf[5586] = 256'h0eff77fe15febbfdabfdbafdfdfd51fee0fe91ff3700cf0031018a019a018c01;
    decBuf[5587] = 256'h49010c01bf0079002700daff94ff42fff5feaffe81fe69fe70fea0fee5fe37ff;
    decBuf[5588] = 256'h9aff12008400eb0049018601a7019d015d01e1006400d2ff48ffeffe9efe8ffe;
    decBuf[5589] = 256'h82fea6feddfe23ff51ff9bffcdff1f006c00b20004013b0145013c010201a100;
    decBuf[5590] = 256'h4300beff41ffeffec3feb6fedafe27ff81ffd6ff3900610085007a005c004100;
    decBuf[5591] = 256'h1800010008001b0037005b00720076005b002e00e9ffa9ff80ff5aff46ff3fff;
    decBuf[5592] = 256'h45ff5fff76ff94ffc6ff04004e009400e6003301510148010e01ad003400a2ff;
    decBuf[5593] = 256'h40ffc3fe92fe83fe91fee6fe5ffff1ffa20018018401bf01ad017d01f8005700;
    decBuf[5594] = 256'hc0ff36ffb9fe88fe7afea2fef7fe5affb7ff0c0059009f00bb00e400eb00f200;
    decBuf[5595] = 256'hec00e600d700c000ab00880055000900afff42fff8feb5fe91feb2fef8fe6fff;
    decBuf[5596] = 256'he0ff4800a500e20003010d010401eb00b70086004e001a00f7ffccffa4ff95ff;
    decBuf[5597] = 256'h90ffa5ffd8ff16004f008400a600a0008f006b0038000800d0ff9cff79ff66ff;
    decBuf[5598] = 256'h77ff9bffceff0c0046006b0080007a00520024000500e9ffeeff17006100a700;
    decBuf[5599] = 256'hf9001a0124010801cf007c002f00c1ff5aff17ffc2fe8bfe81fe9cfef7fe7dff;
    decBuf[5600] = 256'hfaff8c0015016f019f01ae01bc01970160010601b1003800c7ff5fffe7feb6fe;
    decBuf[5601] = 256'h8afeb2fed6fe23ff7dffd2ff35009300e80035017b01a801b1018b014d01f300;
    decBuf[5602] = 256'h8500010084ff32ffe9fec0feb4fed5fe1bff5bffa5ffebff3e008b00d1001001;
    decBuf[5603] = 256'h3a015f01660153012c01f400b00070002600e0ff8eff41fffbfecdfec5fedbfe;
    decBuf[5604] = 256'h19ff74ffe1ff48008b00e0001701490165015c013701f9009e003100caff6cff;
    decBuf[5605] = 256'h30fff9fe03ff1eff47ff9affe7ff41009600cd00ff002c0145014c0138010001;
    decBuf[5606] = 256'hbc006a000700a9ff54ff1dffebfed0feb7fecefee2fe1bff5effc3ff3b00ad00;
    decBuf[5607] = 256'h4f01bb011d0253024302f9019b01fe006600ddff60ff0effc5feb7fec3fee4fe;
    decBuf[5608] = 256'h16ff56ff80ffa5ffbaffccffddff010034008000c6002a016d01910186016801;
    decBuf[5609] = 256'h1601b30056000100b4ff6eff40ff27ff11ff18ff37ff6affa7fff2ff4c008800;
    decBuf[5610] = 256'hbf00f100e800e000ba008a006b004f00400028000b00e0ffadff7dff5eff42ff;
    decBuf[5611] = 256'h47ff55ff7bffb4ffe8ff26006000b200ff0045018501ae01b60178011d019800;
    decBuf[5612] = 256'h1b0088fffffe82fe31fe04fef7fd34fe97fe2aff020091004801bf010002ec01;
    decBuf[5613] = 256'hda0189015d01ff00c30060001d00b0ff66ffeefe9cfe53fe2afe37fe84fe06ff;
    decBuf[5614] = 256'ha6ff69002001c601070242023002ff017b01fd004b00a4ff38ffaffe79fe69fe;
    decBuf[5615] = 256'h78fea0fef5fe42ff9cfff1ff3e008400c400ed001201270121011001ec00c200;
    decBuf[5616] = 256'h9b0077004d0031000d00edffbeff86ff52ff21ff02ff08ff2cff68ffa2ffd6ff;
    decBuf[5617] = 256'h060019002a004e008100a300c200bd0099005d0033000e0007000d001e003800;
    decBuf[5618] = 256'h460063006f006b004f001500cbff85ff45ff3dff44ff67ff86ffb9ffe9ff1400;
    decBuf[5619] = 256'h310040003b0026000b00f2ffe9fff2ff04001e003e005b007e0095009a007f00;
    decBuf[5620] = 256'h51001900e4ffd0ffd6ffe7fff6fff2ffd4ffa9ff8dff88ff8dffaaffb6ffb9ff;
    decBuf[5621] = 256'haaffa1ffa4ffb4ffd4fffeff2500490073009a00b400c200b5009a006c004100;
    decBuf[5622] = 256'h0e00ecffc0ff8dff5dff31ff15ff06ff14ff3aff5eff91ffc1fff9ff2e005e00;
    decBuf[5623] = 256'h89009a008b00740056002b00f9ffd6ffb7ffa6ffa1ffb8ffd6fff1fff5ffe5ff;
    decBuf[5624] = 256'hcbffa5ff8bff74ff70ff74ff8cffa8ffcbffebff010005000800ffff02000400;
    decBuf[5625] = 256'h07000400f2ffd8ffc0ffb6ffbfffd7ffedfff5ffe3ffbfff91ff65ff49ff3aff;
    decBuf[5626] = 256'h2cff30ff3cff69ffaeff00004d007f009b0092007c0059003a001300e5ffb9ff;
    decBuf[5627] = 256'h86ff64ff38ff27ff22ff1eff19ff25ff3dff53ff6dff7fff95ffa9ffc0ffdcff;
    decBuf[5628] = 256'hf8ff100019002200340058009000b600cb00920031009eff14ffbbfe8afe7bfe;
    decBuf[5629] = 256'h89feadfee4fe16ff56ffa0ffd2ff000008001000fbffe8ffd7ffc8ffbaffadff;
    decBuf[5630] = 256'hb1ffbcffcbffe0ffe2ffe0ffd1ffbbffa1ff89ff73ff59ff47ff3eff4cff69ff;
    decBuf[5631] = 256'h8cffacffb9ffb5ffabff9bff87ff6fff5aff40ff27ff1eff2cff49ff74ff90ff;
    decBuf[5632] = 256'hb4ffc2ffd7fff2ff18003c005d0072005f00380000009eff41ffecfe89fe61fe;
    decBuf[5633] = 256'h54fe75fea7fefafe47ff79ff94ffbdfff2ff300059006f0068003d00ffffc5ff;
    decBuf[5634] = 256'h82ff42ff08ffd3fe96fe7dfe93fed1fe3cffa4ff37009900f20023013201ef00;
    decBuf[5635] = 256'h8200e0ff48ff98fef1fd85fd4afd5cfd8dfdf4fd87fe38ffdeff7600d8003101;
    decBuf[5636] = 256'h620171014801f4007b00e8ff5fff06ffd5fea9fe80fe5cfe25fe1bfe36fe91fe;
    decBuf[5637] = 256'h17ffb7ff2400ad00e300f300c7009e003100caff52ffe0fe96fe6efe62fe6dfe;
    decBuf[5638] = 256'h8bfecbfe26ff7affddff3b005f0080007600800077004300f7ff9dff18ffbefe;
    decBuf[5639] = 256'h8efe7ffea7fee4fe1bff61ffb3ff00005a007e0073001900acff45ff02ff0eff;
    decBuf[5640] = 256'h2fff61ff7cffa6ffbcffecff180034002500dfff85ff31ffe4fec6fecffee7fe;
    decBuf[5641] = 256'h1cff68ffd6ff7800e40046013401e3005e00bdff51ffc8fe92fe61fe18fe0afe;
    decBuf[5642] = 256'h2ffe92fe25ffaeff2b007d00a900d100f5000001f600db0091003700caff80ff;
    decBuf[5643] = 256'h58ff4cff41ff23ff19ff22ff29ff3eff44ff4aff45ff40ff44ff5fff86ffbeff;
    decBuf[5644] = 256'hf3ff31006a009f00c100c700a00068002400f7ffeeff05000c00f9ffbbff71ff;
    decBuf[5645] = 256'h2bffebfef3fe0aff2cff4bff5cff80ffbcff17008400eb0049016d0178014601;
    decBuf[5646] = 256'hf4007b00e9ff60ff06ffb5fe89fe96febafe07ff61ffcfff36009300d000db00;
    decBuf[5647] = 256'hbd00a200780062004d00470041003c004a0068008b0099007b004100e6ffa9ff;
    decBuf[5648] = 256'h9effa8ffc4ffccffa7ff84ff71ff8effc6ff180065009700c500ff0015012a01;
    decBuf[5649] = 256'h2401f100a50073005800500066007b005c002900ebffc2ffabffb2ffc5ffbfff;
    decBuf[5650] = 256'hb0ffa2ffb7ffeaff35008f00e4001b014d0156015f01570143012301fc00ce00;
    decBuf[5651] = 256'ha2007b0042000e00d0ffb7ffb0ffd2ff0a003f006f009b00c200e60010012c01;
    decBuf[5652] = 256'h450141012b011801f200c3008b002a00ccff77ff40ff4aff9cff15008700ee00;
    decBuf[5653] = 256'h4c018901d6011c025b0285027d023f02c4014601b4002b00aeff3cff10ff1dff;
    decBuf[5654] = 256'h41ff8effe8ff5600bd005001b2010b025d024e020b029e011901c0008f006300;
    decBuf[5655] = 256'h3b0016000b0029008e0006019801fa0130022002d60193013e01db004800bfff;
    decBuf[5656] = 256'h42ff31ff5efff1ffa1004801df011a02500280028f029c026002fd019f011a01;
    decBuf[5657] = 256'hc0006f002500e3ffbeffc9ff0f008600f8005f01a201c601d101ef010a020202;
    decBuf[5658] = 256'hce016701ff00a2007d009e00d00010014a0160018301a201a80198016f012601;
    decBuf[5659] = 256'he000b2009900b000e0000c0149018301d601230255024c021202bf0172014001;
    decBuf[5660] = 256'h25012d01350120010d01080117012e013b012001eb008a0062008600d3002d01;
    decBuf[5661] = 256'h82018d016f0166016e01a301ee0120024e0246022f0228021502f901ac014901;
    decBuf[5662] = 256'hd1005f0016000800fcff1d006300c7005b010b02b102f2020603ad021a029101;
    decBuf[5663] = 256'h1401c300960039001400f3ff110088001a01a401fd010d02fe01d601e201ed01;
    decBuf[5664] = 256'hf701dc01b3017e015c0156015b014201fc008e002700c9ffeeff3b00d1003d01;
    decBuf[5665] = 256'h9f01d501e501f40101020d020202e401a4015a0128010d01e300be009c007c00;
    decBuf[5666] = 256'h6b0071009100b700e500110144017401a001c701cc01ac0174012201bf006100;
    decBuf[5667] = 256'h0c00ebffe1fffdff37007a00cc002f01a80119029e02d4020403bb024202b001;
    decBuf[5668] = 256'hff005900c2ff60ff06ffd6fec7feeffe44ffbdff4f00d8005601c7012f028c02;
    decBuf[5669] = 256'hb102a6026002fb016801df006200cfff6dff38ff07ff33ff76ffb3ff00003200;
    decBuf[5670] = 256'h7100bc0002016601a901cd01d801a60179014f0139010901b8005500c1ff38ff;
    decBuf[5671] = 256'h02fff2fe1eff7cffd1ff1e006400a4000f017601b901c5017801f60032007bff;
    decBuf[5672] = 256'h04ff98fe84fe96fee7fe6cff0d00d0008701ce01e301a9014f01bd003400daff;
    decBuf[5673] = 256'h89ff3fff17ff0bff2cff4aff65ff7eff95ffa9ffc8fff0ff1e00310036003b00;
    decBuf[5674] = 256'h40005e0081009800940059000f00c9ff89ff60ff3bfffdfeb2fe6cfe3ffe37fe;
    decBuf[5675] = 256'h6bfeb7fe11ff66ffc9ff26007b009c00a6008b0040000e00cfffa5ff71ff25ff;
    decBuf[5676] = 256'hb7fe6dfe45fe6afeb7fe39ff92ffa2ff94ff86ff62ff41ff0fffcffe85fe7bfe;
    decBuf[5677] = 256'h96fe01ff86ff030034004300e5ff90ff17ffa5fe21fea4fd52fd26fd33fd88fd;
    decBuf[5678] = 256'h01fe94fef6fe2bff7dffe4ff4100660071003f00daff62ff11ffc7fe69fefcfd;
    decBuf[5679] = 256'h95fd1dfdecfc18fd76fdfbfd55fe85fe94fea1feaefee5fe17ff44ff2bfff7fe;
    decBuf[5680] = 256'hb9fe90fe79fe72fe6cfe5bfe37fe20fe1cfe28fe39fe23fef8fdb3fd86fd6dfd;
    decBuf[5681] = 256'h93fddefd24fe64fe7dfe75fe7cfe69fe59fe2afefffdd7fdd2fdfcfd50fea5fe;
    decBuf[5682] = 256'hdcfee6fecbfeb2fe9bfe79fe34fed0fd72fd05fdd9fcccfcd8fcf9fc03fd0cfd;
    decBuf[5683] = 256'h14fd3afd93fd00fe67fec5fe02ff39ff57ff60ff36ffe4fe6bfef9fd92fd34fd;
    decBuf[5684] = 256'hdffc7cfc1ffccafb93fbb1fb28fcdafc81fd43fec6fe6cffadff0f002100f0ff;
    decBuf[5685] = 256'ha6fff9fe52fe90fd0dfd67fc26fc12fc00fcf0fb1cfc5ffcb4fc17fd90fde1fd;
    decBuf[5686] = 256'h2bfe38fe2cfe21fe2bfe46fe3efe45fe3ffe45fe56fe6ffe7dfe5ffe25feaafd;
    decBuf[5687] = 256'h2cfddbfcaffc87fc62fc57fc61fcb4fc17fdaafd0cfe1efe2efe3dfe80fed4fe;
    decBuf[5688] = 256'h0bff15ffd6fe5afeb9fd4dfd39fd4bfd5bfd4dfd0afde5fcf0fc0efd4efd67fd;
    decBuf[5689] = 256'h50fd20fdf5fc05fd52fde1fd92fe09ff1eff32fffcfeccfe9ffe42feedfd8afd;
    decBuf[5690] = 256'h11fde1fcb4fcddfc19fd50fd96fdb2fdcafde1fd03fe2ffe56fe7afe91fea7fe;
    decBuf[5691] = 256'hb2fec4fec7feb8fe91fe48fe02feb0fd79fd47fd2bfd02fdddfcbafcc1fc0afd;
    decBuf[5692] = 256'h8cfd2dfeeffe3eff85ff9aff60ff4eff3dff11ffb4fe46fec2fd68fd38fd46fd;
    decBuf[5693] = 256'h89fdc6fdfdfd1bfe48fe72feb5fef5fe2fff36ff22fff6fecffeabfe8afe53fe;
    decBuf[5694] = 256'h10fed0fdc7fdedfd39fe93fecffedafed0fed9fef2fe09ff02ffc9fe77fe2afe;
    decBuf[5695] = 256'h0cfe3afea5fe0cff4fff5bff50ff5aff75ff8eff96ff58ffdcfe5ffeedfdfcfd;
    decBuf[5696] = 256'h5afedffe5cffadffbcffafffa3ff98ff7aff4cfff1fe9cfe65fe6ffeaffe1aff;
    decBuf[5697] = 256'h82ffc5ff01000c001600e9ff9eff44ff08ffd1fedbfef6fe0fff25ff3aff66ff;
    decBuf[5698] = 256'hbaff2700ac00e200d100a50047000b00eaffb8ff41ff8efee8fda7fd09fecefe;
    decBuf[5699] = 256'hb9ff9700ed003b01b201f3012e02f80166013f0019ff59fe36fe55fee5fefffe;
    decBuf[5700] = 256'h47ff87ff11001d01dd014502e701e400aaffd7feb1fed4fe72ffc8ffe2ff5900;
    decBuf[5701] = 256'hf000f001e4024303b302fc01c700f5ff81ff5fff3fffe9fe03ff1bffb2ff8a00;
    decBuf[5702] = 256'h5301d6011d02dc01c801b701c701d60193010d016c00d5ff9affacfffdff6500;
    decBuf[5703] = 256'ha700cc00030149019b01fe012602e9018601f30091007f00b000fa0022011601;
    decBuf[5704] = 256'hf50013016501de01700284024e02bc013301d900c90013013b012f01f800c600;
    decBuf[5705] = 256'hcf002a019701e001ee01990136010e014a01ad010b02480253025d0266026e02;
    decBuf[5706] = 256'h67022902ad010c01a00065007700a800f1001a013e017501e3014a02c302f302;
    decBuf[5707] = 256'he502a2027d0272029002ac02b4027f023402c6015f010101c4008d006f007800;
    decBuf[5708] = 256'ha200f4006d01ff01b0025603c203d603c4035203eb028e023902ec01a6015401;
    decBuf[5709] = 256'h1d01ff000801310165019601c101e9010d023f0270028f02ab02ba02bf02cc02;
    decBuf[5710] = 256'hc802a8028202540235023a025e029102b302ba029e026f023702e50198013e01;
    decBuf[5711] = 256'h0101e000fe003e01990106026d02cb0220036d039f0395034b03f10284023a02;
    decBuf[5712] = 256'h2d0221020002e201a20189019101c101120249023f02ff01c501be01fc016702;
    decBuf[5713] = 256'hec0221031103aa024c024002a3021c036d034103ad02d6014601f7003f01ab01;
    decBuf[5714] = 256'he601f801c701b801e0016602060347033403da0289023f02320256024b022d02;
    decBuf[5715] = 256'h0002e701ee01110249026f0283029602b202c102b4027402eb0189012f014001;
    decBuf[5716] = 256'ha7011f029102bd02cb02bf02ca02e802f102e802a5024102e301a6019b01cd01;
    decBuf[5717] = 256'h0d0247025d023b020f02f301f8012b024e0247020902af0172016701c1012e02;
    decBuf[5718] = 256'hb3020c031d03490356037b0386035403cb02a4017d00beff9bfffaff89000c01;
    decBuf[5719] = 256'h8301ef015102f202b40337044f04b70307033102db01c101d801c30188012f01;
    decBuf[5720] = 256'hfe006501f801a902f0028402d301fe006e008800cf001001fc00eb001b01be01;
    decBuf[5721] = 256'hd702e30392047204e203f702590276025c024402ad01ad00b9ff5aff77ffc6ff;
    decBuf[5722] = 256'h3c00a800e3003d01ef01c5028e031104f9038d03040387023502ec01a9015401;
    decBuf[5723] = 256'h1d0127016701c20116022102ef017901e70084004f005f006e009600ba00c500;
    decBuf[5724] = 256'he3004801f601cb02950317042f04c3033903bc026b022102a901d600d3ffdffe;
    decBuf[5725] = 256'h80fe9dfe1fffc6ff88000b01b101740293035304bc045d045a032002f900edff;
    decBuf[5726] = 256'h3effdffec3fe45ff1b0057017e028b03f3039403cb02e00103013900b7ff11ff;
    decBuf[5727] = 256'ha4fe91feeafebdffc000b40152026f0255020e0223028602bb02ab020902f000;
    decBuf[5728] = 256'he3ff35ff15ff6bff85ff9dff87ff9bff3c002a0146020603e3024502b601ff00;
    decBuf[5729] = 256'hb70077008a0055002400f8ff20007500c200cc008c0052002c00410054003800;
    decBuf[5730] = 256'hebff46ffcffe10ffe8ff24014b020b03e8028902f901ab016401f800470012ff;
    decBuf[5731] = 256'h40fe80fda3fd80fe49ff000047005d004900a3003501be01d0013e0166009dff;
    decBuf[5732] = 256'h4eff66ffa7ffbbff3eff0dff57ff1f00ce017f034703e201e3ff07fe4efdf7fd;
    decBuf[5733] = 256'h2afe42fd72fbc2f9faf92bfcf7ff9603f0058305910382023002100354031f02;
    decBuf[5734] = 256'hd5fe8bfb8cf8f0f8b4fa98fd8aff2fff39feeefd42ff6e017903bd031601e7fd;
    decBuf[5735] = 256'hc4fb60fb70fcaffe90ff4cff92fe5afe59ffb4014f030503a10061feebfca7fc;
    decBuf[5736] = 256'hdcfd14fe7bfd7dfba1f9dff9d8fbc4feb5001001190039ff7dffb100ab02ef02;
    decBuf[5737] = 256'hc30022fea9fb56fbccfca8feddffc4fef9fcc4fbfdfb2efece002901320091fd;
    decBuf[5738] = 256'h18fbc6faa6fb82fd3bfe93fd2efca3fbc9fc09ffed0118030802c9ff53fe0ffe;
    decBuf[5739] = 256'hc8fe00ffcdfecffc6bfad0f81bf9f7fa22fd03febffd05fd3dfd3cfedeff6701;
    decBuf[5740] = 256'h3401efff74fe0ffde1fc0bfd98fca3fb87fa7af929fac4fbbdfd11ff4fffa6fe;
    decBuf[5741] = 256'h0dfedffd09fe2ffec7fd6bfc26fb54fac7fa46fcabfd36fe64fd57fca9fb08fc;
    decBuf[5742] = 256'h44fdbffef2fe0afe8ffc2afbfcfa7afb3afca3fc04fc75fb26fbcdfbe6fcf2fd;
    decBuf[5743] = 256'h5bfefcfd33fdb0fcf7fc64fd9efd45fd51fcd2fa39fa67fa3afbfafb1cfcbefb;
    decBuf[5744] = 256'ha1fbbbfb32fcf4fc43fdfbfc64fcdbfbedfb9ffc16fd2cfda2fcdefb5bfbd2fb;
    decBuf[5745] = 256'hc0fcdcfd4ffee7fd09fd40fcbefba6fb90fb07fb1efa41f9b1f8cbf8d1f90bfb;
    decBuf[5746] = 256'h31fc3efd32fed0fe9aff1c00040017ffbbfd19fc01fb68faddf9b2f98cf9aff9;
    decBuf[5747] = 256'hcff95efa49fbe8fb77fc5dfc45fc5bfc96fceffc61fd70fdf7fc24fc5bfb0dfb;
    decBuf[5748] = 256'hf5fa61fb12fc88fcf4fc57fdb0fde1fdd2fd5afd86fc84fb8ffab2f922f9d4f8;
    decBuf[5749] = 256'hecf858f908fa3dfbb8fcb7fd42fe6dfef9fdd7fdb7fd61fd12fd6cfca9fb27fb;
    decBuf[5750] = 256'h0ffb7bfb05fc82fc51fcaffb17fbdcfa12fb84fbebfbdefba1fb54fb5efbe7fb;
    decBuf[5751] = 256'h98fc0efd4ffd3cfd06fd16fd7dfd11fe4bfe16fe63fd5efc6afbccfaaffa95fa;
    decBuf[5752] = 256'hdcfaf2fa2cfbaafb7dfc80fd2efe8dfe70feedfd18fd4efc98fb50fb66fba1fb;
    decBuf[5753] = 256'h42fc30fdcefd97fee5fefdfee7fe5efe99fdaefcd1fb7bfb2cfb44fbb0fb12fc;
    decBuf[5754] = 256'h6cfcddfc80fd42fe2dffccffafff2cff56fe54fda5fc86fc69fc83fc3cfcfbfb;
    decBuf[5755] = 256'h0ffcaffcc9fd22ff0a008800150021ff04fe91fd29fd48fd2bfdddfcc5fcdbfc;
    decBuf[5756] = 256'h64fd70fe7dffe6ff0500affff8fe52fee6fdabfd75fd24fdf8fcd0fc0cfd9bfd;
    decBuf[5757] = 256'h73fe3cfff3ff6a00ab00bf0089003800b3ff12ff4ffecdfd56fd40fd7bfdd5fd;
    decBuf[5758] = 256'h46feaefe26ff98ffffff42003600e9ff8fff22fff5fe03ff27ff5effa4fff6ff;
    decBuf[5759] = 256'h43009d00f200fd00cb006700d4ff72ff3cff4cff5bff68ff5cff51ff6fffc1ff;
    decBuf[5760] = 256'h5000b200e800b70050000d0001004e00d00029015a012e01eb00f70018014a01;
    decBuf[5761] = 256'h53012a01e700b900d20024018701af017301e4005a00010032007b00f4004501;
    decBuf[5762] = 256'h7101b401f10128025a0251021702d30194018b01c0010b0251029102cb02e202;
    decBuf[5763] = 256'he802bd026802b201c70068004c009a0011015201b401e9015b02fd02c0034304;
    decBuf[5764] = 256'h8a044904c0034303d102a50297028b023e02f801dd01f5014802c1025303b503;
    decBuf[5765] = 256'h0f041f041004b3032d038c02f5016c0136016701b00144021b031e0412052f06;
    decBuf[5766] = 256'hef06cc062e062b05ab03ac02c5019a0174019701b7014602fd0202043c050f06;
    decBuf[5767] = 256'he9058005e2041904fe03460487049a046504d20370038203b30338049104c204;
    decBuf[5768] = 256'hb304db0418059105e205f1057805e6045d04e0038e0380038d03b10314048d04;
    decBuf[5769] = 256'h1f05a80502061206e605d805e405d905bb057c050005a6047604a20400053c05;
    decBuf[5770] = 256'h3105ff04f6041f05900563062c077b076307f70646067005a70425047e033d03;
    decBuf[5771] = 256'h5103ce03a104a40598067607050854086c082b08a107b9069c05dc042e040e04;
    decBuf[5772] = 256'h2b04ae045405c0054a06a306150741074e072a07c7064f06fd05ef05c6058a05;
    decBuf[5773] = 256'h53050d052805a40569061f07c607db07a0078f077e07ab079d07180753063405;
    decBuf[5774] = 256'h74040b046a043305ea05320647068206b8064a07d3072d081c089807d3065006;
    decBuf[5775] = 256'hda05c405d805ea05fa0509064b06a0061907ac070e08430813088e07ed062a06;
    decBuf[5776] = 256'h7305fd04bc04cf042905dc0582064407c7070e08f907be074107cf064a06f105;
    decBuf[5777] = 256'ha0059105d4052906a2061307400732072607ef06e506b7067e062b06b2056105;
    decBuf[5778] = 256'h52057a05b705ee05f80501062a069b062d07b6071008bf073a0799062d06f205;
    decBuf[5779] = 256'hbc056b050405a6049a04290501060407b20792073c078506df0548050d059004;
    decBuf[5780] = 256'hfd03c303d40367048d05b406c1072908ca073b07b8064106aa05f9045304bc03;
    decBuf[5781] = 256'h8103b6032804e8046a05b205c705b405a205920565052205e604af047d046104;
    decBuf[5782] = 256'h49042304f303c703d8032504ca04a00530067e0637069f05ef04190450039902;
    decBuf[5783] = 256'hf301b2019e013f022d03490456050406e5058f050c056604ce0345038002c901;
    decBuf[5784] = 256'h82019801fa01e202c0038904a3045c041b04b903830352032603e3027602f101;
    decBuf[5785] = 256'h9801670176019e01f3015602b402f00211030703da02a0025c02f80180010e01;
    decBuf[5786] = 256'ha7007f00bb0060013602ff0282039a035903cf027602e4015a019600abffcdfe;
    decBuf[5787] = 256'h3dfe23fe6bfe58ff7500820176021403a4038a034203800295017800b8ffc4fe;
    decBuf[5788] = 256'h26fed0fd81fd99fd05feddfee0ff1a01ec015f023c029e01d500eaffcdfe0dfe;
    decBuf[5789] = 256'h19fdbafc9efcb8fc8efd90fecafff100b1011a02bb01f1000600aafe66fd93fc;
    decBuf[5790] = 256'hd3fbb0fb91fb21fca3fc79fd42fe2dffcbffe8ffcefff8fe2ffe78fdd2fc91fc;
    decBuf[5791] = 256'ha5fcb7fcc7fcb8fcc5fceafc37fd91fde6fdf1fdd3fd5cfdcafc19fc73fb07fb;
    decBuf[5792] = 256'hf3fa29fb9bfb1ffc9cfc0efd58fd65fd71fd50fdf6fc71fcf4fb41fbcafab5fa;
    decBuf[5793] = 256'ha1fa8ffa7ffa70fa98faedfa7cfb06fc83fc73fceefb71fbfffad3fac5faa1fa;
    decBuf[5794] = 256'h54fafaf9d6f9f7f979faf6fa26fbbffa2cfaa3f9b5f926fac9fa09fb80fa98f9;
    decBuf[5795] = 256'hbaf864f8e7f88df950fa6afa52fae6f9f9f953faa4fab3fa20faf9f8d2f75ff7;
    decBuf[5796] = 256'h3cf79bf72bf879f8c1f8d6f838f9b6f907fa16fad3f935f972f8f0f7a9f768f7;
    decBuf[5797] = 256'h2df71bf72bf775f7edf75ff8c6f8d4f897f876f880f8aef8b6f872f8eaf7c3f6;
    decBuf[5798] = 256'hf1f57df5e6f584f614f762f7aaf7eaf725f87ff88ff845f87df740f6c2f59cf5;
    decBuf[5799] = 256'h4af627f77ef763f7edf655f6f3f529f67af66bf60ef6a1f557f5b4f56af68af7;
    decBuf[5800] = 256'hfdf720f882f7b8f66af652f611f6aff5c7f429f4d2f321f456f57cf689f7f2f7;
    decBuf[5801] = 256'h11f8bbf76df725f78ef6b6f5b3f405f4e5f33cf4f3f499f505f619f607f637f6;
    decBuf[5802] = 256'h64f68cf698f64bf6ddf576f54ef55af57bf571f568f55ff576f5cff524f65bf6;
    decBuf[5803] = 256'h3df6ebf588f560f584f5a5f5c3f596f52af5c3f4d0f425f5caf5d0f6f2f6d3f6;
    decBuf[5804] = 256'h7df6faf5b3f59df5b1f57bf52af5c3f49af4eff494f59af648f768f7d8f655f6;
    decBuf[5805] = 256'haff518f5ddf4eff4fff42bf553f5a8f5f5f54ff6a4f607f74af76ef74df7dff6;
    decBuf[5806] = 256'h3df67af5f8f4e0f44cf5fdf573f6e0f6f3f605f7f5f604f711f7d4f671f6f9f5;
    decBuf[5807] = 256'hc8f5d7f56af642f7d2f7ecf7a5f738f7fef60ff740f76cf75ff70af7d3f6c9f6;
    decBuf[5808] = 256'he5f63ff794f79ff76df740f737f78af703f875f8a1f85ef809f8bcf7daf73ef8;
    decBuf[5809] = 256'h9cf8d9f8b8f85ef821f842f8b0f835f98ef97ef934f986f810f8faf7e6f740f8;
    decBuf[5810] = 256'h91f8bdf81bf988f90dfaaefa1afb55fb43fbf1fa8afa12fac1f959f931f9f5f8;
    decBuf[5811] = 256'hd4f8caf8f7f841f9c3f988fa3ffbe5fb51fc8cfc57fc26fcfafb9cfb5ffbfcfa;
    decBuf[5812] = 256'h9ffa7afa85faf3fa78fbf5fb26fc35fc42fc66fcc9fc42fd73fd46fdb3fc03fc;
    decBuf[5813] = 256'h8cfb76fbb1fb2efc5ffc8bfccefc3bfdddfda0fe23ff3afffafe97fe1afeeafd;
    decBuf[5814] = 256'hdbfdb3fd8efd41fd0ffd2bfd85fd23febafe44ffc1fff2ff0000f3ffb6ff69ff;
    decBuf[5815] = 256'h23fff6fefefe42ffb8ff2a00af00e4001501240131012501d8006a00e5ff68ff;
    decBuf[5816] = 256'h17ff43ffd6ffae0077012e027602b602ca02dc02ab027f023c02cf0185017801;
    decBuf[5817] = 256'hb4012d02c002220357036803590366035a0365036f0342030803d302bf02ea02;
    decBuf[5818] = 256'h3f03f503ac045205be05f9050b06da0590053305ad043004df03b303c0031504;
    decBuf[5819] = 256'h8e0441051606a606290740072b07f006ba064906ff05d7059a058f059905eb05;
    decBuf[5820] = 256'h64063707c7077e08c508b00875081b08eb07dc07cf07aa079f07a907c507fe07;
    decBuf[5821] = 256'h42085d0876087d0869088808d1082b099809e209ef09fc09f109d309c909c109;
    decBuf[5822] = 256'h8d09780972098309bb09f009040a170a110a0c0a3f0a8b0ad10a110b290b040b;
    decBuf[5823] = 256'hfd0a100b2c0b6e0b9c0b830b6d0b3d0b2a0b5d0ba80bee0b1c0c240cf00bcd0b;
    decBuf[5824] = 256'hae0b920bb60bdf0b120c500c8a0cbe0c0a0d3c0d330d1a0dd60c600c0e0ce20b;
    decBuf[5825] = 256'hd50b2a0c8d0cea0c3f0d760d940dd40dfd0d140e1b0ed60d5f0dee0cc10cb40c;
    decBuf[5826] = 256'hd80c0f0d190d220d1a0d220d7b0de80d4f0ead0eb90e820e780e810e9a0ecf0e;
    decBuf[5827] = 256'hc80e6a0ed70d260d800c6a0c7e0cd70c290d900d080e9a0e4b0ff10f5d104a10;
    decBuf[5828] = 256'ha90fbb0e9e0ddf0c760c560c3a0c880cff0c960d950e890f2710b7109d10f70f;
    decBuf[5829] = 256'h090f2c0e620dab0c350c9d0b8a0b9c0b2e0c2d0d670e390ff90f621042105f10;
    decBuf[5830] = 256'hdc0f360f480e2c0dd20b470bc90aef0a580b350cfe0cb50d8b0e540fd70fef0f;
    decBuf[5831] = 256'h570f580e1e0d4c0c8c0b230b040b5a0b740beb0b820c5a0dea0da10eb80e4c0e;
    decBuf[5832] = 256'hc30dfe0c130cb40b240bd60aee0ad80a130b490b9a0bc60b090c2d0c220c2c0c;
    decBuf[5833] = 256'h110cd70bd00bc90baa0b990b600b0e0bd70aa50a770a6f0a3b0a0a0af809e709;
    decBuf[5834] = 256'hec091f0a330a2d0a1c0a030af5091b0a490a680a630a350ad709940957092009;
    decBuf[5835] = 256'hee08af0854082f083a085808ab08cc08d608ba0880083d082208f807c407a107;
    decBuf[5836] = 256'h690735072e0734073a0753075807540750074c07430740071e07e20698063e06;
    decBuf[5837] = 256'hd005870544051f05fe04f404100539056e05ab05f60514060b06d1056f05f704;
    decBuf[5838] = 256'ha6045c043404f703d603a40377035e038303a603c503bf039b0356032403f602;
    decBuf[5839] = 256'hee02d802b5027d0249022602130219021e02100204020002fc010c021a020302;
    decBuf[5840] = 256'hd4016d0105018d003c00d4ffacff88ff7dff9bffdbff36008a00d700cd00b200;
    decBuf[5841] = 256'h89002700caff75fffcfeabfe61fe39fe45fe7cfe86fe7dfe53fe10febefd87fd;
    decBuf[5842] = 256'h69fd60fd78fd80fda2fdc2fddefdedfdd6fd96fd32fdd4fc7ffc5efc40fc25fc;
    decBuf[5843] = 256'h0cfcd8fba8fb88fb8efb9dfbbefbd3fbcffbbefb95fb6efb4afb17fbd9fa9ffa;
    decBuf[5844] = 256'h5cfa1cfaf3f9cdf9d4f900fa27fa5ffa94fa9bfa6ffa31fae7f98df950f919f9;
    decBuf[5845] = 256'hbff883f836f82cf847f870f896f8aaf87ff836f804f8e8f7e0f7e7f7e1f7cef7;
    decBuf[5846] = 256'hd3f7e3f728f882f8a7f870f8eef729f772f6ccf560f54cf55ef54ef55cf5baf5;
    decBuf[5847] = 256'h27f6acf64df7b9f7cdf797f705f754f6ddf546f5bdf463f412f403f4f6f332f4;
    decBuf[5848] = 256'h95f40ef580f5e7f52af636f6fff5cdf556f5c4f43bf49af32ef3f3f2e1f2f1f2;
    decBuf[5849] = 256'h58f3b6f30bf458f48af4b7f4c0f48bf440f4faf3baf390f389f374f33cf3f9f2;
    decBuf[5850] = 256'h94f251f25df294f2eef243f34ef330f315f3fcf2f5f2eef2c2f279f233f2f3f1;
    decBuf[5851] = 256'hfbf14ef29bf2e1f20ef317f31ef325f32bf30ff3cdf244f293f11cf1dbf0eff0;
    decBuf[5852] = 256'h25f155f182f1c5f101f238f292f2cff2f0f2e6f2b8f28ff25af21df2f3f1cef1;
    decBuf[5853] = 256'habf180f158f10bf1d4f0b6f09bf0d5f045f1d8f161f2def20ff33bf32ef3f1f2;
    decBuf[5854] = 256'h8ef216f263f1bdf051f016f028f099f01ef1bff156f2b8f212f343f351f329f3;
    decBuf[5855] = 256'hedf274f2e1f17ff102f1b1f0c0f0cdf00af157f19df1eff168f2b9f220f37ef3;
    decBuf[5856] = 256'h8af369f337f3c0f26ff225f2e2f1bef1c9f1bff1daf1f3f10af21ef257f26df2;
    decBuf[5857] = 256'h9df2d5f2fbf21df349f365f389f3b3f3b8f3a9f39bf36cf341f324f3f6f2bef2;
    decBuf[5858] = 256'h8af259f253f29cf2f6f27cf3f9f34af476f49ef47af46ff465f425f4ebf3c6f3;
    decBuf[5859] = 256'ha4f3b6f30bf447f494f4daf4e3f4ecf4f3f4d1f4b2f48af448f42cf434f45af4;
    decBuf[5860] = 256'hb3f420f56af5adf5eaf50bf651f67ef676f651f605f697f54df525f501f522f5;
    decBuf[5861] = 256'h54f5a6f509f69cf625f7a2f7f4f7e5f7a2f735f7b0f657f626f617f625f649f6;
    decBuf[5862] = 256'h80f6c6f64ff7d8f755f8c7f8f3f801f9dcf8a5f873f858f83ff838f815f8eaf7;
    decBuf[5863] = 256'hcef7bef7c3f7e9f736f883f8ddf84af994f90cfa5dfa8afa97fa73fa26fae0f9;
    decBuf[5864] = 256'hd7f9cef9e5f9f9f9f3f9e2f9ddf9d9f910fa53faa5fadcfa0efb18fb30fb65fb;
    decBuf[5865] = 256'h95fbc1fbf3fbfafb00fcfbfb00fc17fc2cfc30fc34fc2afc22fc2afc44fc5cfc;
    decBuf[5866] = 256'h78fc93fcb3fceafc3dfd8afdd0fdfdfd06fe0dfe22fe34fe45fe55fe47fe21fe;
    decBuf[5867] = 256'hf2fdd3fde4fd12fe4afe8efecefe18ff72ffdfff29006c0060003f000d00dfff;
    decBuf[5868] = 256'hb6ff90ff89ff83ff94ffb8fffdff6b00f0004901bb01e701f5010102f601d801;
    decBuf[5869] = 256'haa0181015c01550167018f01c701fc013a0273029902bb02e7020e033c035c03;
    decBuf[5870] = 256'h780387039503a203c503ee030a041a040304d4039c0385037e03b70318049004;
    decBuf[5871] = 256'he204490556057b05860590059905b205b905ce05d405ce05d305e105dd05e105;
    decBuf[5872] = 256'heb05e805f705140636067c06c206ef0629074f0771079d07c407e807ff07fb07;
    decBuf[5873] = 256'hd807c107b407b007d007ee07f107fc07f907fc0723086c089e08f0083d095b09;
    decBuf[5874] = 256'h77098f099709ac09be09a2099d098f0969095a09550959098409cd09ff09510a;
    decBuf[5875] = 256'h880aa60ac10ada0ae20ae90aef0ac70ab80ab30ab80ae20a0a0b190b1e0b220b;
    decBuf[5876] = 256'h260b530b8c0bb10bd30bda0bc90bce0be50bfa0b250c410c320c2d0c200c150c;
    decBuf[5877] = 256'h1f0c1c0c020cf10bee0bf00b180c6c0ca90ce00c260d410d7b0da00d9a0d7a0d;
    decBuf[5878] = 256'h310dc30c790c510c450c7c0cae0cee0c280d5c0d710d840d890d7a0d880d950d;
    decBuf[5879] = 256'ha80ddc0d110e180e120eea0d9d0d660d340d190d110d270d2e0d5a0d8c0dca0d;
    decBuf[5880] = 256'h150e470e500e580e320e100efd0df80df30d130e200e240e350e250efa0dcf0d;
    decBuf[5881] = 256'h910d460d3c0d460d5e0da20de20d1b0e5f0e9f0ea70ebe0ec40ea50e7e0e500e;
    decBuf[5882] = 256'hfe0dc70d950d560d3d0d350d4a0d820da80dd80d040e200e2f0e460e530e470e;
    decBuf[5883] = 256'h4b0e350e100eec0db90d6d0d3b0d200d070d2d0d4f0d6e0da10dc30dd60df20d;
    decBuf[5884] = 256'hf70de00dcb0da80d750d530d330d0c0d070d020df60c010d0c0d020dff0ced0c;
    decBuf[5885] = 256'hce0cd20cee0c0d0d4d0d680d700d5a0d380dff0ccb0c9b0c560c280cff0be90b;
    decBuf[5886] = 256'hfd0b100c160c250c200c140c1f0c380c4e0c790c8b0c7b0c800c690c3a0c1b0c;
    decBuf[5887] = 256'he80b9c0b560b160bed0ae60adf0ae50a0c0b300b510b880b9e0b980b780b460b;
    decBuf[5888] = 256'h080bef0ad90ac40abe0aa20a730a540a430a340a390a3d0a310a270a0b0ae809;
    decBuf[5889] = 256'hda09c509b109bc09c509d309eb09ee09cf09a80970092c091109e808c208ae08;
    decBuf[5890] = 256'h8e087208630868086c089608b308c208d008c308a808960874083808ee079407;
    decBuf[5891] = 256'h3f07f206d406cb06e30609071007230733074d076d077a0767074007fe06ac06;
    decBuf[5892] = 256'h5f062d0611060906f205c205a305700540052e0533054305630589059905a605;
    decBuf[5893] = 256'ha205870561053205fa04b70477043d041804f503e203d203b80398037a036603;
    decBuf[5894] = 256'h55035e0367037f03a703cf03e803ed03be036d03f4028202fd01a40153012601;
    decBuf[5895] = 256'h340158018f01e9013e0275027f0264022a02e60182012401b70050000d00d1ff;
    decBuf[5896] = 256'hc6ffe4ff23006e00a000bb00c3008f005100f6ffa1ff54ff0efff3fedafec4fe;
    decBuf[5897] = 256'haffea9feaefeb4fecbfed7fedbfecafea1fe63fe19febffd6afd33fd15fd0cfd;
    decBuf[5898] = 256'h25fd59fd97fdc0fdc8fdc1fd95fd41fdecfc89fc2bfcd7fba0fb6efb64fb7dfb;
    decBuf[5899] = 256'hb2fbf0fb29fc40fc47fc1bfcd2fb8cfb3afb03fbe5fac9fab1fa9afa85fa73fa;
    decBuf[5900] = 256'h6dfa68fa63fa5ffa4cfa2cfa0efae4f9bcf9a3f979f95df958f94af94ef962f9;
    decBuf[5901] = 256'h6cf976f984f97cf962f93bf9f9f8a7f844f801f8c4f7b9f7c3f7dff708f81ef8;
    decBuf[5902] = 256'h41f86cf87df882f875f83df8ebf79ef744f707f7d0f6b2f697f68ff6a5f6c7f6;
    decBuf[5903] = 256'h0cf74cf786f79cf795f76af737f7ebf6a5f678f63ef60af6d9f5aef59df5a2f5;
    decBuf[5904] = 256'hb0f5c5f5fff528f65df68df693f68ef66af624f6caf58ef557f539f554f55cf5;
    decBuf[5905] = 256'h73f588f58ef593f599f58bf56df552f52bf512f504f5eff4ebf4fcf4fff413f5;
    decBuf[5906] = 256'h36f543f550f54cf526f5f8f4d8f4bcf4c1f4e2f4eff4f2f4f6f4e0f4ccf4c4f4;
    decBuf[5907] = 256'hb3f4a9f4abf49ff49df4aaf4acf4b8f4cbf4c8f4c6f4d5f4c7f4c2f4c0f4aaf4;
    decBuf[5908] = 256'h8df48af486f48ff4a9f4a6f4a9f4b2f49ff4a6f4c6f4d4f4d8f4e4f4c4f4a7f4;
    decBuf[5909] = 256'h93f482f478f481f479f477f492f49ef4bef4ecf4fff405f514f50ff514f51ff5;
    decBuf[5910] = 256'h0ef5fef4f6f4cef4a7f4a2f48bf486f49af4a4f4c0f4f3f415f534f545f536f5;
    decBuf[5911] = 256'h31f535f532f53cf552f54ff547f54ef53ff541f555f54df546f53bf51df5f7f4;
    decBuf[5912] = 256'hf2f4e4f402f53cf565f5a8f5e8f512f628f63df62af603f6dff5a3f569f534f5;
    decBuf[5913] = 256'h04f5fef41af53ef57af5d5f511f65ef6a4f6c0f6c8f6c1f675f61bf6c6f579f5;
    decBuf[5914] = 256'h47f53ef557f59af5ecf539f693f6d0f607f739f742f719f7e4f699f63ff602f6;
    decBuf[5915] = 256'he1f5d7f5f2f52cf661f69ff6d8f6fef62ef74df748f738f718f7e9f6bdf6b8f6;
    decBuf[5916] = 256'ha8f6bff6eef60df740f77ef7a7f7bef7d2f7c0f798f774f738f70ff7f8f6e4f6;
    decBuf[5917] = 256'heaf611f735f77bf7c1f713f84af890f899f8a1f88bf85bf816f8e8f7aef798f7;
    decBuf[5918] = 256'hadf7ccf70af854f89af8b5f8cef8b8f8a3f89df88cf872f86ef858f854f882f8;
    decBuf[5919] = 256'hbaf80df95af98cf9a7f9aff999f992f97ff963f93ff928f90af906f918f934f9;
    decBuf[5920] = 256'h57f981f99df9c1f9eaf912fa40fa52fa58fa53fa45fa38fa34fa38fa35fa38fa;
    decBuf[5921] = 256'h4afa64fa92facafafefa21fb40fb46fb41fb3cfb27fb0cfbe5fac1faaafaaefa;
    decBuf[5922] = 256'hbafad9fa08fb40fb75fbcefb0bfc58fc8afca5fcaefca6fc91fc72fc56fc3cfc;
    decBuf[5923] = 256'h1cfc0ffc04fc00fc16fc2afc4cfc76fc92fcc0fcecfc1ffd4ffd87fdacfdc1fd;
    decBuf[5924] = 256'hc7fdb6fda7fd99fd8cfd89fd9afda3fdacfdbefdd4fdf3fd1afe3efe55fe6afe;
    decBuf[5925] = 256'h76fe87fe90fe93fe91fe8afe7bfe79fe8cfeb3fef1fe2bff5fff90ffa2ffbeff;
    decBuf[5926] = 256'hceffdcffe0ffcdffadff87ff6dff72ff87ffb2ffd9ff070033004f0069007700;
    decBuf[5927] = 256'h83007f007c0085009900b600d90003011f0143015a016f018301860183017a01;
    decBuf[5928] = 256'h680161015f0165016a016f01730180019501ba01f3012702570283029402a302;
    decBuf[5929] = 256'hba02c702cb02ce02bf02b602a902a202b502c702d802e702f102f60202031503;
    decBuf[5930] = 256'h2703420353035c03710383039d03c403f203110438044804430436041304ea03;
    decBuf[5931] = 256'hce03b403a603b303d603f6032d047104b104da040f051505280523050905f204;
    decBuf[5932] = 256'he504c204b4049f049304a504c704e80427056705a105d605ea05f005eb05d105;
    decBuf[5933] = 256'ha8058b05720551054505500562059105cf05f8053b06690682069806ad06a706;
    decBuf[5934] = 256'ha10692067a06760672066f06720675066d066f067e069406bf06eb0607072107;
    decBuf[5935] = 256'h2f073b074f0760076a07720770076d076f07750774077f07870788079807ab07;
    decBuf[5936] = 256'hb307c407d307d507eb070808230842084f084b084f0852084f0861086d086708;
    decBuf[5937] = 256'h65085f08570868087f089508c008df08fc081f0937093b093f09340918091409;
    decBuf[5938] = 256'h0a09000914092c093c0956096709640972097a0978098f09a509b309cb09e109;
    decBuf[5939] = 256'he409f609020a080a160a1f0a1e0a310a430a460a590a660a5f0a610a5b0a410a;
    decBuf[5940] = 256'h350a2b0a1b0a240a360a500a850ab90adc0a200b4e0b670b7d0b760b570b3b0b;
    decBuf[5941] = 256'h0d0bee0ae80aed0af20a0f0b1b0b260b3b0b500b5d0b720b750b630b600b620b;
    decBuf[5942] = 256'h6c0b870bb10bc20bdc0bea0be50b000c0b0c080c100c090cee0bf90b020c050c;
    decBuf[5943] = 256'h220c2e0c1c0c190c0b0ce90bdb0bd60bc30bce0bdd0bec0b130c460c680ca00c;
    decBuf[5944] = 256'hd50ce90c090d0e0df50cdd0caf0c760c510c210ce90bd20bcb0bb80bd50bf80b;
    decBuf[5945] = 256'h220c600c9a0ca10cb60cbc0cab0cbb0cc80cc40cd00ccc0caa0c930c750c520c;
    decBuf[5946] = 256'h4e0c410c1e0c100cfb0be70bf90b090c170c2f0c320c230c260c240c190c270c;
    decBuf[5947] = 256'h250c1a0c240c2b0c2a0c3b0c500c4d0c4b0c350c0a0ceb0bb80b7a0b510b2c0b;
    decBuf[5948] = 256'h090b030b090b040b1b0b380b4c0b720b8c0b9a0baf0bbb0ba90ba60b860b580b;
    decBuf[5949] = 256'h2c0bf90abb0a920a7c0a590a530a420a290a240a200a1c0a260a230a150a170a;
    decBuf[5950] = 256'h100a0a0a140a1d0a1e0a2c0a2e0a220a150afa09c00987094309f108ba089c08;
    decBuf[5951] = 256'h6e0866085f086508850896089b089f088a086f0856084108270823081a081108;
    decBuf[5952] = 256'h0f080708fd07f307d9079e0765072107cf069806660638062006090602060906;
    decBuf[5953] = 256'h0e061e063e065c066f06730669064a062306eb05a70555051e05d80498046f04;
    decBuf[5954] = 256'h5904520458045204580453043e042a041204e903c20394036803410327031903;
    decBuf[5955] = 256'h0c030103fd02fa02f702ea02d902ba0287024902ff01b90179012e01e800bb00;
    decBuf[5956] = 256'ha2009b00af00c200e900f90007010201ef00cf00980055001500cbff99ff59ff;
    decBuf[5957] = 256'h40ff29ff15ff02ffe6fed7febffea2fe77fe50fe22fef6fdcefdabfd93fd87fd;
    decBuf[5958] = 256'h7bfd71fd6dfd65fd4dfd31fd16fdf6fcd9fcb6fc8cfc5afc1cfcd1fb9ffb72fb;
    decBuf[5959] = 256'h49fb23fb0efbfcfaf6fafbfa00fb15fb11fb00fbd7fa99fa3efa02fab5f983f9;
    decBuf[5960] = 256'h67f94ff947f94ef954f965f96af966f948f916f9bcf867f81af8d4f7a7f78ef7;
    decBuf[5961] = 256'h77f77ef791f797f7a6f7bdf7b0f795f76ff722f7d5f68ff64ff615f6fff5f8f5;
    decBuf[5962] = 256'hfef50ff61ef62cf631f615f6f6f5d0f58df53bf504f5aaf46df44cf442f44bf4;
    decBuf[5963] = 256'h64f47bf482f494f48ff48af485f45ff426f4f2f3a6f360f345f32cf325f32bf3;
    decBuf[5964] = 256'h25f320f325f30ef301f305f3e5f2b6f297f259f220f218f2f6f1eff100f2fbf1;
    decBuf[5965] = 256'hf7f10cf208f204f214f200f2e8f1d9f1b3f18ff178f152f12ef12af10cf1f8f0;
    decBuf[5966] = 256'hfcf0e0f0d4f0d1f0bbf0a7f0a9f08ff085f088f079f081f09bf0a6f0aff0c9f0;
    decBuf[5967] = 256'hbff0aff0a6f07ff058f048f015f0e5efd3efabef9cefaaefbfefd2eff9effeef;
    decBuf[5968] = 256'h03f00ff00bf016f026f01df015f01cf005f0fbef0af0fdeff1efeaefccefafef;
    decBuf[5969] = 256'habef92ef8fef98ef90ef9cefb7efbbefcdefefefebefefeffaeff0eff9ef19f0;
    decBuf[5970] = 256'h1df029f041f03ef041f04ef034f02af020f001f0ebefe7efcfefccefe6eff0ef;
    decBuf[5971] = 256'h13f045f05af079f095f0a5f0bcf0daf0def0e8f0f1f0ddf0dbf0f0f0edf0f5f0;
    decBuf[5972] = 256'h0af102f1f5f0f7f0e0f0d6f0e5f0ddf0e4f004f112f127f152f16ef192f1cef1;
    decBuf[5973] = 256'he6f10cf22ef235f23af24af23cf237f243f232f228f22bf213f210f21ff21cf2;
    decBuf[5974] = 256'h28f248f24cf26af28df2adf2d4f216f344f36df393f3a7f3baf3d6f3d1f3d6f3;
    decBuf[5975] = 256'he2f3dff3cdf3d0f3b6f3acf3b5f3adf3aff3c5f3c7f3daf3fdf32cf464f4a7f4;
    decBuf[5976] = 256'hd5f4eef413f528f53bf54bf551f55ef56bf567f572f58ef59af5abf5c7f5cbf5;
    decBuf[5977] = 256'hc8f5c4f5b6f5a9f5b0f5aef5c0f5e4f512f64af67ef6aff6e7f61bf73ef75df7;
    decBuf[5978] = 256'h79f774f779f77df779f77cf786f783f786f791f794f7a2f7bcf7cff7e8f704f8;
    decBuf[5979] = 256'h0ff828f857f879f8b1f8e6f808f928f944f949f957f96cf978f982f992f99af9;
    decBuf[5980] = 256'ha2f9b8f9c6f9d8f9eef9f6f9f9f9fbf9f5f9fff916fa32fa55fa88fab8fae3fa;
    decBuf[5981] = 256'h16fb46fb65fb82fb9bfba9fbadfba2fb97fb8efb7ffb82fb8efba1fbb9fbd5fb;
    decBuf[5982] = 256'he8fbfafb1cfc3cfc5afc7dfc8bfc98fca3fca7fcbdfcd7fceffc11fd32fd47fd;
    decBuf[5983] = 256'h62fd82fd97fdaafdaefd9efd90fd88fd81fd87fd99fdaafdcafdf3fd26fe56fe;
    decBuf[5984] = 256'h82fea9fec3fed1feccfec9fec5fec2fec5fecdfeddfefdfe30ff6effa8ffdcff;
    decBuf[5985] = 256'hffff110022001d000f00faffe7ffd5ffd2ffe0ff080046007f00c30003013c01;
    decBuf[5986] = 256'h620177018901780169015b014e014b015c017e01b101e1010d02350258027002;
    decBuf[5987] = 256'h74027f027502650262026a027b029b02c402ec021a033903610384039c03b103;
    decBuf[5988] = 256'hc403cf03d203e003f803140437044e0452045604530449044c044f0451046404;
    decBuf[5989] = 256'h77048704a704ec041e055e059805be05ee050d0613062c063a06470662067a06;
    decBuf[5990] = 256'h8a069e06ab06ae06c106d306e40604072407310754077d07a507d3070b083108;
    decBuf[5991] = 256'h61088c08a908eb08190953098709c509de09030a260a380a490a4e0a400a450a;
    decBuf[5992] = 256'h410a440a600a830aa40ae30a230b5d0bb00be70b190c6b0ca20cc00ced0c060d;
    decBuf[5993] = 256'h1d0d4d0d5f0d700d8a0d980d940d9f0d9c0d8c0d8f0d8c0d8a0d9d0db50dd10d;
    decBuf[5994] = 256'h0b0e450e6a0eb60efc0e290f630f890f9d0fb00fb60fb10fbe0fb20f970f8c0f;
    decBuf[5995] = 256'h760f570f5b0f570f4c0f560f590f510f740f980fb90ff00f241047107f10a510;
    decBuf[5996] = 256'hc710ff1025113911591169116411691165114a1138112211f710fd10ec10dd10;
    decBuf[5997] = 256'hfd1024113d118311dd1119127c12da12fe124b137d139913c213d813c413e313;
    decBuf[5998] = 256'he913ee130e142c14301456146614611476148a149414c314e51405155915ae15;
    decBuf[5999] = 256'hfb156916d0162e179b1702182a187f18a0189618b218991873186c185a183e18;
    decBuf[6000] = 256'h571878188418be1819195619b919161a531aa01ad21aed1a271b5c1b701ba91b;
    decBuf[6001] = 256'hdd1bf21b2a1c5e1c731c9f1cb01c961c9b1c851c4b1c431c2d1c0a1c1d1c441c;
    decBuf[6002] = 256'h541c991c071d331dac1dfd1d0c1e4f1e5b1e501e461e2a1ef11de91dd41db51d;
    decBuf[6003] = 256'hc61dd51dc81ddd1de11dc81dd81dcf1da81dad1da81d881d9d1da91d971db31d;
    decBuf[6004] = 256'hbf1dae1dbd1dba1d931d8d1d5f1d0e1dd71c911c1a1cc91b621b041baf1a781a;
    decBuf[6005] = 256'h1e1afa19d919bb19c419bc19a519ac19991967194419f31890183318ad170c17;
    decBuf[6006] = 256'ha016171676150a15a8144e14fd1396131d13ac124412b1112811ab1019108f0f;
    decBuf[6007] = 256'h120fa00e570e2e0ef20dd10d9f0d5f0d150da70c220c810bbe0a080a32096908;
    decBuf[6008] = 256'h7d07df06160693054c05e0047e042504d3038a032c03d7025e02ec0185010d01;
    decBuf[6009] = 256'h9b003400f1ff9cff4fff1dffeffeb6fe72fe32fed7fd83fd0afd77fceefb71fb;
    decBuf[6010] = 256'hdffa7cfafff9cff9a2f97af96ef98ff999f9a2f9bbf995f965f914f9b1f839f8;
    decBuf[6011] = 256'hc7f742f7e9f698f64ef626f61af6f9f5eff5e5f5bcf588f54af5eff482f438f4;
    decBuf[6012] = 256'hc0f34ef322f3dff2a2f297f28df284f28cf267f21bf2d5f15ff1acf035f073ef;
    decBuf[6013] = 256'hbcee15ee7eedf5ecbfec6eec24ec31ec0dececebceeb6aeb0ceb9feafde93ae9;
    decBuf[6014] = 256'hb7e8e2e752e7cfe629e6bde582e505e5b4e44ce4d4e321e3abe2e8e131e18be0;
    decBuf[6015] = 256'hf3df43dffcdebbde80de92de81de90deb8de94de5dde2bdea2dd19dd9cdce9db;
    decBuf[6016] = 256'h43dbd6da26daafd96ed933d9fed8edd8dfd8d1d8f6d8d5d8cbd8d4d8bbd8b4d8;
    decBuf[6017] = 256'hd6d8d0d8ecd82ed94ad973d9c6d9d1d9efd90adae1d99dd982d917d9cdd88ad8;
    decBuf[6018] = 256'h35d814d81ed803d81bd86ed8a5d8d7d83bd963d9a0d9edd90bda26da60da68da;
    decBuf[6019] = 256'h7cdac1dacada04db56db77db95dbd5dbcddbd5dbdbdba3db6fdb4cdbefdaacda;
    decBuf[6020] = 256'h87da50da5ada88daa1dae4da49db8bdbf9db7ddcb3dc04dd4edd41dd4ddd58dd;
    decBuf[6021] = 256'h4edd57dd70dd77ddb5dd10de65dedede70dff9df9ae05de1dfe1b5e27ee301e4;
    decBuf[6022] = 256'hd7e4a0e557e62de7f6e778e84ee9dee995ea3bebfeebb5ecbaedaeee8bef01f1;
    decBuf[6023] = 256'h66f2abf37af52af7b3f87efa2efcb7fd82ff33012c038004300649071409480a;
    decBuf[6024] = 256'h610b600ca50d770ed10fb810df1139137d14a4154a17d318381ada1b621dc71e;
    decBuf[6025] = 256'hc6201a22ca235325b8265928e229472b8c2cb22dbf2eb32f913020316f31b631;
    decBuf[6026] = 256'ha031b4317e312d31e330a03064306f3079308230dd3032316931c331e731dc31;
    decBuf[6027] = 256'hbe3147317430ab2f8b2e322ded2b722a0d292528ff26f225fe2420241e232a22;
    decBuf[6028] = 256'h4c211020e91e901dee1b651a00195f17d615d71436131d121e11da0fb30e590d;
    decBuf[6029] = 256'hb80b2f0afe07f3051704eb01750099fe65fd4cfc19fc8efb64fb8afb67fb08fb;
    decBuf[6030] = 256'hecfa35fa5ff923f8fcf656f5cdf368f223f1fcef3cef8eee2feed9edbfedd7ed;
    decBuf[6031] = 256'hc1edaded9bedaced9dedaaedb6ed03ee5deee3ee84ef1bf0ccf072f109f293f2;
    decBuf[6032] = 256'hc8f2d9f2acf284f217f2b0f152f116f10bf13df18ff11ef2f6f2bff376f44bf5;
    decBuf[6033] = 256'hdbf52af641f600f69ef521f54ef44bf39df2bff1f6f074f0cdef8cef79ef43ef;
    decBuf[6034] = 256'h33ef42efffeec2ee8bee09ee68edfcec24ec22eb73ea96e993e8e5e7c8e608e6;
    decBuf[6035] = 256'h14e537e434e340e223e1cadfe2de67dd68dc23dbfcd9f0d841d864d7d4d652d6;
    decBuf[6036] = 256'hdbd56fd534d5b7d445d4c0d3fcd245d26fd16cd078cf9bced1cde6cc87ccf8cb;
    decBuf[6037] = 256'hdecbf5cb0bcc46cc9fccd0cc37cd7acd9ecdbfcdddcdc2cdbacdd0cdbccde7cd;
    decBuf[6038] = 256'h3ccea9ce4bcf39d016d153d2ced333d577d647d8f7d980db4bddfbde84e0e9e1;
    decBuf[6039] = 256'h2ee355e4aee539e60ce7cce7eee70ee82be811e8f9e7e3e7a8e773e783e774e7;
    decBuf[6040] = 256'hb7e724e8a9e86ee98dea9aebd4ec4fee4eef92f0b9f1c6f274f352f4a8f4c2f4;
    decBuf[6041] = 256'haaf413f462f38cf250f129f01def9ded9eecb6ebe4ea24ea01eae1e9c4e9dfe9;
    decBuf[6042] = 256'hc7e95be9f9e810e833e7f7e5d0e476e332e25fe19fe037e017e034e0b6e0fee0;
    decBuf[6043] = 256'h95e1f7e150e281e272e24ae226e2d9e1a7e18ce183e17ce190e197e17be157e1;
    decBuf[6044] = 256'h11e17be062df56de61dd03ddacdc63ddc7de5ee142e5eae98def5ff6cafca002;
    decBuf[6045] = 256'h7209dd0f0814d217e319831a151b901a2719ba188f17ea173c18b2198e1b351e;
    decBuf[6046] = 256'h632162241a27492a6c2c252fe9302933ca354338cc3b173fcb436e49bc4e8e53;
    decBuf[6047] = 256'hf057105d826062623b65c0654765da647664676314635f632b64606559673569;
    decBuf[6048] = 256'h616bd76ca36de06d386d076b666838655e61bf5d655b66583c57e156d8574e59;
    decBuf[6049] = 256'ha25ace5cd95e2d606b60a360a45fa65d425b5d58de549351ba4d1a4ac047e743;
    decBuf[6050] = 256'h4740fd3c23397b341930f92a27268420361b64160212290f9c0d330ca00c040d;
    decBuf[6051] = 256'h7d0f18112413001534166c169f16b815e81338123f10630eb30c2a0bc509dd08;
    decBuf[6052] = 256'h0a08fe064f06f30452035901f5fe11fc1ffaa6f766f586f442f47ff478f6dcf8;
    decBuf[6053] = 256'hc1fb07000304ac080e0d0a11a013eb160f19001bc51c601e401f1c21cc22e523;
    decBuf[6054] = 256'h16262128fd29292c9f2df32e27304031733145316f31fc301f317d310d322d33;
    decBuf[6055] = 256'h1f35fb361e3a1d3dd53f04430246bb48344bcf4c454e114fca4f7350a6507750;
    decBuf[6056] = 256'h4d50da4fe64ec94d234c2a4a3e47864457417e3dde3994369533dd30182f212e;
    decBuf[6057] = 256'h6c2e382fe830e132bd34e9365f382b396939c0385b375d35f932702f262c2729;
    decBuf[6058] = 256'h6f26f523b621151f501db51b3f1a6318b3164a146511ad0e330cf4095307d904;
    decBuf[6059] = 256'h3e035e020a01cc009400c7009900c3009c007a001b00c4ff42ff2affe9fefdfe;
    decBuf[6060] = 256'h56ffe8ff7200360185019d015c0184000eff43fd9cfa22f8e3f5d7f3fbf142f1;
    decBuf[6061] = 256'h7af113f2b5f3aef59af852fb81fe7f01710380047705c205f6043c04b4024f01;
    decBuf[6062] = 256'h0a008ffe2afd42fc6ffbaffa47faa9f9a6f8b2f756f6b5f4bbf257f0bceeb1ec;
    decBuf[6063] = 256'hd5ea25e97ce87de74fe725e74be76ee78ee771e7eee678e68ae56de460e3e1e1;
    decBuf[6064] = 256'h7ce094df6dde60dd6cdcd1da48d97dd7d6d4a8d1a9ce2acbeec615c46dbf4cbc;
    decBuf[6065] = 256'h73b9e5b77cb634b597b53db534b614b7e0b71eb8e5b7b2b7cbb64fb5eab3a6b2;
    decBuf[6066] = 256'hd6b0a2aff9aefaadccad4aae71aed9ae77af07b021b098b057b01cb02eb0ddaf;
    decBuf[6067] = 256'hecaf7fb008b1f1b14cb391b460b611b89ab999baddbb07bc2ebc0bbc6dbbddba;
    decBuf[6068] = 256'h8fbae8b9feb960ba96ba28bb27bc90bc2ebdf7bdddbd96bd80bdcfbc29bc14bc;
    decBuf[6069] = 256'hb1bbc3bb97bc26bd7abebfbf91c051c1ffc161c125c0aabe13bce4b8e6b52db3;
    decBuf[6070] = 256'hffafb6aec5acb5ab08ac52ac1eadcfae77af10b09bb071b0b1af77aefcac31ab;
    decBuf[6071] = 256'h81a9f8a793a608a635a50fa578a597a5b4a5cea528a565a446a3a0a117a04c9e;
    decBuf[6072] = 256'h9c9c139b149a2c99ad9887981e98ff976f978496a795dd945b94d1941696cd98;
    decBuf[6073] = 256'ha29e22a637af32ba88c44cd30fe191edf0f846034d07670d830e810deb08c004;
    decBuf[6074] = 256'h72ff9ffa7ef7a5f418f381f480f7fffa2b005f06340c06139c17721dc0229227;
    decBuf[6075] = 256'h342d8232b63836404647874f83593960c3684f6e5f751f78a07ade792d794c77;
    decBuf[6076] = 256'h97750a74917324734e7413765378f37a6d7d087f537f877e5b7c257970740f70;
    decBuf[6077] = 256'h126c6a674964b76332638c658b68d16cf1716375c5799d7c2b7eb27db47a6d76;
    decBuf[6078] = 256'h4e71ba69aa62695aa55291497743b33ba8363c30672a95232a1d54178210170a;
    decBuf[6079] = 256'h41047700a4fb83f8aaf526f5aef4f6f521f730f8cbf9acfaf0fa36fa1ef9edf6;
    decBuf[6080] = 256'h4cf41df144eda4e969e56de1cddd83daced56cd170cdc8c866c446bf74ba12b6;
    decBuf[6081] = 256'h39b3a3b039afa7afd1b0b5b45db900bfd2c512ced6d5e6dc27e5b3eabeef7ef2;
    decBuf[6082] = 256'hfff445f7f5f755f7e6f762f7eaf67cf6a7f701f89cf912fbeefc1aff25018903;
    decBuf[6083] = 256'hc905d407380a780c190f471246158c19881d3122d327212d54332a39fc3f9244;
    decBuf[6084] = 256'h674ab54f275389573e59d55b4d5ce05bb55aa659665730543151794e954aff47;
    decBuf[6085] = 256'hb444b641c43f4b3d543c743bb83bf53b0e3d733e71404d427944ef45cb478448;
    decBuf[6086] = 256'hbc482348de466644ed41c03dc3391b35b930992bc7266522691ec91a7f17a513;
    decBuf[6087] = 256'h0610bb0cbd0904078b04a601b5ff3bfdfcfa1bfac7f88af8c2f8f5f8ddf903fb;
    decBuf[6088] = 256'h10fc04fd21fee1fe49ff69ff13ff90febafd7efc03fb38f90cf701f59df2b9ef;
    decBuf[6089] = 256'h00ed87eaa2e7eae425e38ae114e0d0df0ee0b7e082e2ade44ee77dea7bed34f0;
    decBuf[6090] = 256'hadf2edf4f8f64cf805f93df970f942f9c4f851f8e8f7c8f772f78cf7a4f7baf7;
    decBuf[6091] = 256'hf4f72af81af8eef7abf725f7a8f616f665f5bff47ef443f455f4c7f487f5a6f6;
    decBuf[6092] = 256'hfff7a1f99afbfefd3e00490225045a0572060b07dd060a066404fb0117ff97fb;
    decBuf[6093] = 256'h5cf75ff3c0ef85ebace815e6bbe398e16de013e0c1df0be0d7e015e14de180e1;
    decBuf[6094] = 256'h52e1d4e060e06cdf8fde8cdd98dcfadb6adb1cdb04dbeeda02db14db04dbbada;
    decBuf[6095] = 256'h42da4ed914d899d6ced4a2d201d088cd48cbd2c96ec7d3c588c5bcc4fac413c6;
    decBuf[6096] = 256'h78c719c9f3cbabcedad1b3d553d99ddc9cdf54e2cee40ee783e84fe984eabcea;
    decBuf[6097] = 256'hefeac1ea42ea83e9d4e8b8e75ee61ae54ae39ae111e046de11ddf9db60db8edb;
    decBuf[6098] = 256'h61dc6dddedde1ee129e38de571e863ea27ecc3ed0deed9ee9ceef3ed5aedcfec;
    decBuf[6099] = 256'ha8eb9ceaa8e98be832e7ede51ee46de274e088dd97db1dd939d647d483d28cd1;
    decBuf[6100] = 256'hacd0f0d02ed1d6d1d5d2bdd390d44fd5b8d598d57cd5f9d453d465d388d24bd1;
    decBuf[6101] = 256'h24d018cf24cec8cc83cb08ca3dc88dc604c5d3c25dc181bf4cbe34bd35bcaabb;
    decBuf[6102] = 256'h2bbb05bb9cba3dbae7b999b9b1b973bafbbb45bf80c3e7cafbd3f7de41ecc3f8;
    decBuf[6103] = 256'h620725153a250a30de39ce426d44f3429c41823bbe33ae2c6d24a91c9e17de14;
    decBuf[6104] = 256'h09144f16c019631f3526a02c20342c39973fc2430846da4afc4d1b53ee57905d;
    decBuf[6105] = 256'h6264cd6aa370f175c47ae57d777efb7ea17ca3792376e871c86c56697667c065;
    decBuf[6106] = 256'h3c65a566c868816bfa6ddf70d0722b73d8726371876fdf6c666a2668b0666c66;
    decBuf[6107] = 256'h2667af68e06a806dfa6ff1703b71e76f406da8680563af5aeb52d7494c418839;
    decBuf[6108] = 256'h79320d2c3826ea20b61a8c163e116b0c09080d045bfe91fa20f7fef326f1a1f0;
    decBuf[6109] = 256'h19f187f178f33df534f6a9f7ddf6a9f5cff289ee69e935e3b5dba5d43ace64c8;
    decBuf[6110] = 256'h16c344be23bb4ab8b3b559b336b144af80ad40abcaa976a8bda766a831aa53ad;
    decBuf[6111] = 256'h08b2ebb856bf81c80cd1d0d8dfdf4be675ea3feef0ee50ee9aec04eab9e6bbe3;
    decBuf[6112] = 256'h02e189deeddc38dd7cdd2cdf96e1d6e30ce7e5ea7cedc6f0a0f448f96afc8901;
    decBuf[6113] = 256'h5c06fe0bd0123c19111fe3254e2c7930c735d837b9396e3bf33b7b3b0d3be339;
    decBuf[6114] = 256'h8839da39253a793bae3c373e363f1e409c40dc3fa23e7f3c48394a3691336330;
    decBuf[6115] = 256'h3f2e152dba2cb12dbc2fa83261358f38b33aa43c4a3c533bb238cf342630842a;
    decBuf[6116] = 256'h3625031f2d19df136d104c0d730ae6088c06430552038d014effadfc33faf4f7;
    decBuf[6117] = 256'he8f594f460f327f3c0f3a8f423f622f7c4f86cf905fa7af9a7f8b5f651f46cf1;
    decBuf[6118] = 256'hb4ee85eb87e895e61ce4dce166e012df62ddd9db74dad3d84ad7e5d5fdd47fd4;
    decBuf[6119] = 256'hf2d4e6d581d7ead973ddbee0bce33ce796e9b9ebe4ec3eed47ecd2eaf6e84ee6;
    decBuf[6120] = 256'hd5e395e11fe053df9aded2de6bdfb0e0d7e197e28be329e47fe4cee415e556e5;
    decBuf[6121] = 256'h06e63be7b6e8e7ea88ed01f0e6f29ef518f8b3f929fbf5fbb7fb7ffb80fa3bf9;
    decBuf[6122] = 256'h69f8a9f740f720f704f71ef765f74ff7c6f601f67af480f2a4f0fded84eb44e9;
    decBuf[6123] = 256'hcee77ae6c1e5f9e592e633e8bce921ebc3ecdbed74eea3ee79ee6cedeceb87ea;
    decBuf[6124] = 256'h89e835e785e56ce46de3e2e264e23de2d5e176e1e6e02fe05adf57de63dd85dc;
    decBuf[6125] = 256'h2fdcacdb95db01dc8adc2bdd44de04dfb2df90e059e1dce1b1e27be366e482e5;
    decBuf[6126] = 256'hdce67de806ea6bebb0ec82eda9ed40ed63ecb3ea0ce893e5aee22fdfd5dcb2da;
    decBuf[6127] = 256'h87d978d825d870d83cd971da89db54dd0edeb6de4fdf7ddfffde8cde98ddbadc;
    decBuf[6128] = 256'hb8db7eda57d94ad810d795d530d48fd206d13bcf8bcd92cb3eca09c961c8c8c7;
    decBuf[6129] = 256'h99c7c3c736c89fc8fec854c93ac9c3c82cc806c78ac525c484c2fbc096bf52be;
    decBuf[6130] = 256'h2bbd6bbc77bbd9ba49ba92b9bcb8f3b79fb65bb5e0b315b264b0dbae10addcab;
    decBuf[6131] = 256'hc3aa2aaa58aa2bab6badf3b02fb572bbf2c207cc02d758e16dedccf81606050f;
    decBuf[6132] = 256'h2517931b9a1fd220b61faf1c191844127a0ea709c60711069606e009950e3714;
    decBuf[6133] = 256'h8d1c5124612bcc31a237743e09433447fe4ad14f33542f58e05daa61de67096c;
    decBuf[6134] = 256'h5771c974a9765f78da7762773e758672a26e036ba9686067c4678869c86bfe6e;
    decBuf[6135] = 256'hd8727776c279c07cb27e0c7f5f7f7e7ea27c6e7b75799977df76567557747073;
    decBuf[6136] = 256'hf4712970826d9f69ed639f5e6c58eb50dc499b410f3cff3469303f2c75286326;
    decBuf[6137] = 256'h42238d21f61e9d1c9e19e616b713b910000e870b47093c0760052b04a202d700;
    decBuf[6138] = 256'h27ffbdfc35f9eaf535f193eb45e612e03cdaeed41cd079caafc69ec47dc1c8bf;
    decBuf[6139] = 256'h3abec2bd54bdf1bc96bce9bc33bdffbd34bfbdc0eec28fc5bdc8bccb3bcf77d3;
    decBuf[6140] = 256'h4fd6e6d840db88dcb3dd0ddebbdddbdc0fdcdada32daffd98adab1dba3dd8fe0;
    decBuf[6141] = 256'h0fe43be90eeeb0f382faed00c306950d2b1200184e1d21228326a22b142f3532;
    decBuf[6142] = 256'h0e35a5370e39563aba3a143bc23a4c39f83748364f34fb32c6318e3127328234;
    decBuf[6143] = 256'h0b38463c89425f48314f7257fe5c09629f667467366825660463075f56590854;
    decBuf[6144] = 256'hd54dff473544c340a23ded3b5f3af638d236a8352e33ef304e2ed42b95298927;
    decBuf[6145] = 256'had25f4249d253626d727d029ac2b5c2d052ed22d8d2c152a32268921271d0818;
    decBuf[6146] = 256'hd411a90ddf096e068d04fb036e02f50188012401ca00d3ff5dfe09fd59fb40fa;
    decBuf[6147] = 256'h41f959f82ff8a2f80bf9a9f972fa8dfaa4fa0dfae7f86bf73af52ff343f052ee;
    decBuf[6148] = 256'hd8eb3dea5de909e84fe7a7e60ee626e5abe346e2a5e01cdf51dd1cdc74dba7db;
    decBuf[6149] = 256'h8fdc5ede05e134e432e7b2eafced20f011f221f3cff2eef19af06fee63ec87ea;
    decBuf[6150] = 256'h5ce8e6e692e5d9e4c0e327e39ce2c9e1bde083df5cde02dd1bdc48db22dbffda;
    decBuf[6151] = 256'hdcdb18dd93de5ee08ae295e4e9e51ee7c7e7fae76ee748e6eee4aae3dae12ae0;
    decBuf[6152] = 256'ha1ded6dca1db18dab3d812d7f9d5c8d353d277d0c6ce3ecda5cc19cc44cc9dcd;
    decBuf[6153] = 256'h3ecfa8d1e7d31ed741d9fadb09dd00de4bde7fddcedb46da15d809d62dd47dd2;
    decBuf[6154] = 256'hf4d0c1d036d0b4d028d190d12ed2bed20cd324d365d379d3aed320d4a5d48dd5;
    decBuf[6155] = 256'haad603d848d96fda7bdb6fdc0eddf1dc6edcf7dbdedad2d9ded882d73dd66ad5;
    decBuf[6156] = 256'h5ed4afd311d30fd21ad13dd03acf00ce82cd75ccc7cba7cb8bcba5cb1ccc5ccc;
    decBuf[6157] = 256'hbfcc3ccd0bcda4cc11cceaca1bc96bc701c5c1c24cc1e8bef1bd7bbcafbb71bb;
    decBuf[6158] = 256'haabb77bb48bb1ebbabbafdb91fb91cb8e3b6bcb5afb401b463b3d3b2b9b271b2;
    decBuf[6159] = 256'h31b2f6b19cb10ab159b0b3afc5ae27aed1ad83ad9aaddbad16aedbae92af38b0;
    decBuf[6160] = 256'h7cb11eb317b58bb8c6bc09c38acaa2d5f8df0dec6cf7b6043911981cfa230128;
    decBuf[6161] = 256'haa2b8e2a87271c219b199014250e4f088d073e085f0ba21123193722322d8837;
    decBuf[6162] = 256'hee40e94b4b5352576c5d885e8e614f64cf66996a0b6e6c726976117bf27ca77e;
    decBuf[6163] = 256'h237ed87aff764d71ff6bcc65a161d75dc65b665c1b5ebb61e766b96b5c71aa76;
    decBuf[6164] = 256'h1c7a3d7df27e777f0d7ec57c0c7a487864757273ae711270726df86a14680663;
    decBuf[6165] = 256'h345e9258c0517f49bb41b03c44366f30292eb72a172a6128dd27642741254f23;
    decBuf[6166] = 256'h2120471c9f173d131d0e4b09e90434039d002500dcfe40ffe5fe4afdd4fbe8f8;
    decBuf[6167] = 256'ha2f482ef4fe979e32bdef8d7cdd303d0f2cd52cde3cd5fcdc8ce35cf99cf3ecf;
    decBuf[6168] = 256'h48ce67cd8bcb57ca3ec90bc9f3c9c2cb6ace4dd2f6d657db54dff3e24de570e7;
    decBuf[6169] = 256'h9be840e8eee70ee742e689e5c1e5c0e661e8cbeaafed67f096f394f64df911fb;
    decBuf[6170] = 256'h51fdf2ff6b025005cf080a0d2a12fd169f1c71230728322cfc2f6e334e35e035;
    decBuf[6171] = 256'h5c35d4354136a5366938a93a4a3d2d41cd441848164b084d174ec54dba4b5649;
    decBuf[6172] = 256'h7146f242a73fa93cb73aa839fa39703b4c3d773f83415f439344cc4433449142;
    decBuf[6173] = 256'h2840e83db23ab337fb3481324230cc2e682c282a1d283125b121761d7a19d114;
    decBuf[6174] = 256'h6f10970df7098e084607a907b908af09bb0b970dcb0e030f360ff20dce0b2d09;
    decBuf[6175] = 256'hff0500034800cefd8ffb19fac5f80cf8f3f6f4f553f4caf299f0f8ed7feb9ae8;
    decBuf[6176] = 256'ha9e6e4e449e394e360e495e58ee76ae995eba1edf5ee29f062f02ff0a3ef7dee;
    decBuf[6177] = 256'h70ed7cecdeeb4eeb34eb4ceb8ceba0ebd6ebe6eb9ceb3febb9ea18ead7e99de9;
    decBuf[6178] = 256'haee961ea37ebadec78eeacef35f100f3baf3f2f325f4f6f324f364f270f1d2f0;
    decBuf[6179] = 256'h7bf02df015f081f0e3f03df1aff1bdf160f1f3f015f038ef35ee41eda3ec86ec;
    decBuf[6180] = 256'ha0ec17edaeed86ee16ef99ef81ef15ef16ee96ec65ea5ae8f6e5b6e3abe1cfdf;
    decBuf[6181] = 256'h1fde76dd77dc8fdb11db04dacad8a4d74ad606d58ad38bd200d2d6d149d23dd3;
    decBuf[6182] = 256'hd9d461d692d808dae4db9ddcd6dca3dcbbdb94daa1d84dd79dd584d485d357d3;
    decBuf[6183] = 256'h2dd353d3bcd31ad471d4bfd4a7d492d47ed448d49ad477d594d63ad8a3dae3dc;
    decBuf[6184] = 256'h19e018e309e519e60fe7c5e671e5c0e3e7e02edeb5dbd0d8dfd61ad5c8d47dd4;
    decBuf[6185] = 256'h49d57ed697d7fcd8e4d962da88da20da42d9ecd835d8bfd7ffd762d802d947da;
    decBuf[6186] = 256'h2fdb01dc74dc0cdcb0da0fd935d67cd34ed04fcd97ca1dc827c7dcc620c755c8;
    decBuf[6187] = 256'hdec9a9cb59cd71ce0acfdcce5ece51cd17ccf0cae4c935c9d6c8bac8d4c81bc9;
    decBuf[6188] = 256'h05c955c850c78ac5e3c269c0e1bc96b973b781b527b579b5efb653b9dbbc26c0;
    decBuf[6189] = 256'hffc39fc7f9c91cccd5ce4ed133d479d899ddcce3f7ec82f57eff930bb213081e;
    decBuf[6190] = 256'hbe24f62512270c24761ff617e610a50819030efe23fd4e0120086110951cf427;
    decBuf[6191] = 256'h3e35c0411f4d8154385be15efd5ffa5ee55f105f4e5e9d5d7e5f3361c1623963;
    decBuf[6192] = 256'h82641e645a621a60e45c0a597456295306516951e353b458e85ebd648f6bd073;
    decBuf[6193] = 256'h5c79637c237f4e7e8c7d1a7af976d971676e056ae6647461525e565aae554c51;
    decBuf[6194] = 256'h094b3345e53f51384633b02e852ac3291329f32acc2d6c31c633c436ef37df36;
    decBuf[6195] = 256'hfb33ed2eba288f1f0417080d5206c7fd3bf830f39aee1aec58eba8eac7e835e8;
    decBuf[6196] = 256'ha8e64ee42be239e0c0dd24dc44db00dbc2da6bdb04dc32dc08dcfbdaf0d8bad5;
    decBuf[6197] = 256'hbbd275ce79cad9c67fc437c3d3c2e3c323c659c932cdd2d01cd41bd7d3d998db;
    decBuf[6198] = 256'h33dd13dedfde14e00de2e9e391e6bfe9beec3df088f3abf5d6f6e5f793f7b3f6;
    decBuf[6199] = 256'he7f5b2f47af413f557f6cff868fdca010d08e20db414201b4b1f152386262727;
    decBuf[6200] = 256'hdc285728df277227d527e528802a212d0431ad350e3a2e3f01442247d7485c49;
    decBuf[6201] = 256'he348e54565422a3e0a39983537315e2ed92d612d842f04333f373c3be43f0543;
    decBuf[6202] = 256'hde456c47f346d0448940693b9736b42f1e2b4925fb1f891c68198f160a16a114;
    decBuf[6203] = 256'h0f15ab145114fe13b4137013b6127e127f11f41076100310540f380ede0c3d0b;
    decBuf[6204] = 256'h4409e006fc03430115fe16fb97f73df53ef286efc1ed81eb76e99ae765e64de5;
    decBuf[6205] = 256'hb4e4e2e461e5bae615e9f9eb79efc3f2c2f57af8f4fa46fb66fa02f879f44def;
    decBuf[6206] = 256'h7aea97e302df2cd962d5f0d10fd07ecf0bd165d364d6e3d91ede1be2bae505e9;
    decBuf[6207] = 256'h03ecbceeeaf10ef438f548f69af64ff683f558f321f023eddce8e0e438e0d6db;
    decBuf[6208] = 256'hfdd867d60dd47ad4ded4a2d6e2d818dcf2df91e3dce6dae95aedb4efd7f190f4;
    decBuf[6209] = 256'h54f64bf72bf86ff8b6f7bdf559f3d0ef95eb75e6a2e100dcb2d640d31fd06ace;
    decBuf[6210] = 256'he5cd4ecf72d1b8d5b5d95ddebfe298e537e9a0eae9eb4cec3debfde8f2e616e5;
    decBuf[6211] = 256'h6ee2aae06adef4dca0dbf0d9d8d873d72ed607d5aed369d296d170d193d170d2;
    decBuf[6212] = 256'he6d317d6b8d831dbbade14e112e4cbe68fe82bea75ea41eb04ebcceacde9e5e8;
    decBuf[6213] = 256'hbee764e620e5a5e340e2fbe080dfe7de5cde32dea5dedfdf5ae18be32ce6a5e8;
    decBuf[6214] = 256'he5ea86ed4aef41f08cf0c0ef8bee02ed6beaf1e7b2e511e34ce156e075df31df;
    decBuf[6215] = 256'hebdf23e056e03ee114e13ae1d1e0f4df2bdf40de23dd63dcfadb9cdbb8db6fdc;
    decBuf[6216] = 256'h15ddaddd85dedbdef5deddde1bde30ddd4db8fda14d9afd76ad643d5d0d422d4;
    decBuf[6217] = 256'hc3d3a6d324d3dcd270d2e7d146d1afd025d0cccfbccfcacf5ed00ed113d24dd3;
    decBuf[6218] = 256'h74d481d500d765d864da50ddcfe00ae52aeabef1cef80f01d308e711721afe1f;
    decBuf[6219] = 256'h0423ef231a23501f1c194713750cdf07b4036e017f03e107240efa185023652f;
    decBuf[6220] = 256'hc43a1a457f4e9954255a275b125c3d5b7b5aca59ea575857d3565b56c9562c57;
    decBuf[6221] = 256'hd256db5590553c5483534b537e531f55f957785ba460d866ad6cfb712f78af7a;
    decBuf[6222] = 256'h797e297f897ed47c3d7a027606725d6dfb68dc636a60c75afd568c53e94d1f4a;
    decBuf[6223] = 256'had464c42733fe53d6d3ddb3d053f7f416344544619486b48f546f942da3d4536;
    decBuf[6224] = 256'h312da72473185310fd0547ff2df9d9f5d2f2e8f1bdf27ff32ff4d0f461f5ddf4;
    decBuf[6225] = 256'h65f41cf3f2f12df092ee87ecabea03e8d5e4fbe053dcb1d663d12fcb5ac590c1;
    decBuf[6226] = 256'hbdbc9cb9e6b76bb8d4b9f8bb3ec05ec530ca92ce8ed237d758da0ddca4de0de0;
    decBuf[6227] = 256'h7be0a5e100e252e29de259e29fe187e088df43dec8dcc9db9bdb19dc59dee1e1;
    decBuf[6228] = 256'h0de741edc1f4d5fd6006240e3415751d012307269d2a722b342ce52c042b722a;
    decBuf[6229] = 256'he5288b264225182453225d211221ce2087218023e4256d29992e6c330e39e03f;
    decBuf[6230] = 256'h76444b4a154e2750c75035509f4d544a9f453e411e3c4b37ea3211307a2d202b;
    decBuf[6231] = 256'hd829ad289e27a7263125dd23a9222021bb1f761e4f1d8f1c271cc81bab1b911b;
    decBuf[6232] = 256'h1a1b831a8419be179315f2120e0f6f0b340737038ffe2dfa31f691f237f039ed;
    decBuf[6233] = 256'h47eb38eae6e930ea84ebb9ecb2ee8ef0baf230f4fcf43af521f456f233ef5aeb;
    decBuf[6234] = 256'hb1e64fe230ddbed99dd6c4d33fd3c7d20fd4c8d6f6d9f5dc74e0bfe3bee6afe8;
    decBuf[6235] = 256'hbfe911eac6e9fae841e8b8e653e50ee493e22ee146e074df01df98deb8de0edf;
    decBuf[6236] = 256'h2de087e128e321e585e769ea5becd4ee14f18af2def397f43ff50cf5def4b4f4;
    decBuf[6237] = 256'hf4f38bf36cf3dcf28ef246f2daf12af183f0c1efd6ee38ee6eedecec03ed19ed;
    decBuf[6238] = 256'hcaedcfee09f030f189f271f344f46af401f424f3aef17def72ed0eebcee82de6;
    decBuf[6239] = 256'h69e429e2b3e05fdf2bde82dd4fdd7eddfcddbcdeb0df0ce1ade2c6e32be513e6;
    decBuf[6240] = 256'h91e66be602e667e46ee292e0ebdd71db8dd89bd6d7d4e0d300d3bcd275d31ed4;
    decBuf[6241] = 256'h1dd561d6dcd7a7d9d3db49dd25df51e15ce3b0e460e679e712e89de873e8b3e7;
    decBuf[6242] = 256'h04e7e8e58ee44ae323e216e1aee04fe06ce022e1c9e1e2e23be480e5fbe660e8;
    decBuf[6243] = 256'ha5e9cbead8eb12ed39ee45ef3af017f1e0f12ff2e7f17bf155f031ee26ec3ae9;
    decBuf[6244] = 256'hbae570e271dfb9dcf4dafed9b3d97fdab4dbaddd99e08ae204e5e8e712e922ea;
    decBuf[6245] = 256'h74ea94e9c8e818e71fe5bbe27be0dadd61db21d916d73ad505d45cd3c3d295d2;
    decBuf[6246] = 256'hbfd232d39bd3bbd3d7d3bdd3e7d2e5d1abd030cfcbcd86cc5fcb86cbeecb89cd;
    decBuf[6247] = 256'hf3cf32d269d542d9d9db23df22e2dae454e738eaf1ec89f1ebf52efc0402d608;
    decBuf[6248] = 256'h410f6c1336174719a718f1164912e70dc708f503140282011904360ab611ca1a;
    decBuf[6249] = 256'hc6251c30303c5044be48c54cfd4de14cdf4b1e49494803465345f345a8472d48;
    decBuf[6250] = 256'h874af44a1f4c794ccb4c164de24d174f805109554459885f5d65ab6adf700975;
    decBuf[6251] = 256'h4f77007860778774e770bb6be96687628b5eeb5a91589355a15392525250b14d;
    decBuf[6252] = 256'h384baf4764444142883f793e273e073f5b400b422443574312429a3f4d3af731;
    decBuf[6253] = 256'hfb27951e9a134409dfff54f700f4f5ee0aeedfeea1efb2f193f348f5c4f44cf4;
    decBuf[6254] = 256'h28f270ef41ec68e8c8e48de090dcf1d8b6d496cfc3ca21c5d3bfa0b975b5abb1;
    decBuf[6255] = 256'h9aaff9aeafb045b380b7a0bc73c115c7dfca51ce32d0c3d03fd0d6ce8dcd9ccb;
    decBuf[6256] = 256'hd7c9e1c896c862c997ca1fcc84cd26cf3ed03dd125d2a0d36bd513d841dbd1e0;
    decBuf[6257] = 256'h1fe6b3edc3f42efbae02b9074f0ccf0e910f4210610eac0c1e0ba60a130b3e0c;
    decBuf[6258] = 256'h6c0f2114c31995200027812e9035d13d5d436848294b544f1650c6502650704e;
    decBuf[6259] = 256'he34c894a8b47d2445942bd40483f7c3eb93ed23f9d4144447347714a2a4d5850;
    decBuf[6260] = 256'ha151cb5226538a517f4f934c4d485044a83f063a3c366931072d0b296c251223;
    decBuf[6261] = 256'hee20fd1eed1df61c161cd21b101cd81b0b1cdc1b5e1beb1ab1198d17ed14be11;
    decBuf[6262] = 256'he50d450a0a06ea0017fcf6f8faf463f2faf0b2ef87ee2dee7feecaee96efd4ef;
    decBuf[6263] = 256'h0cf0d9ef4eef7bee6eeda9ebf9e98fe7abe4f3e179df95dcdcd918d87dd69cd5;
    decBuf[6264] = 256'h58d596d5afd614d8b5d93edb09ddb9ded2df6be0f6e074e19be178e197e141e1;
    decBuf[6265] = 256'h27e1e0e074e0eadf26df3bde1edd11dc1ddb7fda62dab1dab6db7bdda7df48e2;
    decBuf[6266] = 256'h76e550e9e6eb31ef2ff2e8f4acf6a3f783f8c7f88af871f772f674f498f26cf0;
    decBuf[6267] = 256'h61ee85ecd5eabce923e951e9d0e9dcea16ece6ed96ef1ff1eaf2a3f3bcf4eff4;
    decBuf[6268] = 256'hc0f4eef394f2f3f0faee96ec56ea4be86fe6bfe4a6e30de33be3bae3c6e400e6;
    decBuf[6269] = 256'h7be77ae862e98ce919e925e88ae691e4b5e289e07edea2dce9dbd0da9dda6fda;
    decBuf[6270] = 256'h99dabfda28db87db16dc65dcacdc18ddc9dd3fde02dfeddf8be055e140e2dee2;
    decBuf[6271] = 256'h6ee3f0e308e4f2e3b7e3f3e23ce237e143e0e7deffdd2cdd6cdc49dc69dcf9dc;
    decBuf[6272] = 256'he4dd01df5ae0fbe114e379e461e5dfe5b9e596e5f8e4f5e301e3a5e160e08edf;
    decBuf[6273] = 256'hcede20de00de1dde6bde11dfd4df8be061e12ae2e1e2b6e30de4c4e46ae501e6;
    decBuf[6274] = 256'h8be64fe79ee7b5e774e7c4e68fe568e4c2e2c9e075dfc5dd1cdd83dcb2dcdcdc;
    decBuf[6275] = 256'h4fddb8dd16de33de7cdda7dc6adbefd924d874d65bd55cd4d1d3a7d367d415d5;
    decBuf[6276] = 256'h71d613d89bd966db17dda0de6be096e20ce470e654e90decf0ef99f43bfa0d01;
    decBuf[6277] = 256'h7807f90e04146f1aef1c351f241d031ae314b00eda081005ff029f039c075f0f;
    decBuf[6278] = 256'h5b1970250f34e33d654a8552f3564a58125786517b4ce547ba43f03fdf3dfe3b;
    decBuf[6279] = 256'h903c263f90408e430e476749414de0502b54e058415d61623467956b6e6e0571;
    decBuf[6280] = 256'h7d7110711e6fa56c1c69e0640862715f175daa5c0d5d1d5eb85f9860ec612a62;
    decBuf[6281] = 256'h1161ac5ff55c3c5a0e570f541e525950634f184fd44e1b4e024dd14a05475441;
    decBuf[6282] = 256'h823a41324528e01e5516c910b909f9067904b70367040705bd064a08c3083009;
    decBuf[6283] = 256'h3f07c504e1019afd7bf8a8f306eeb8e884e2afdcddd547d171cba7c796c575c2;
    decBuf[6284] = 256'h07c394c4eec6c8ca70cf12d5dcd8afddd0e062e1dde074df9bdbf2d650d102cc;
    decBuf[6285] = 256'h2fc70ec459c2ddc247c445c78ccbabd07ed520dbeadebde3dee693e82aeb93ec;
    decBuf[6286] = 256'hb6eea8f021f361f56cf7c0f871fafafb93fcd7fd52ff8301ba046e09100fe215;
    decBuf[6287] = 256'h4e1c2322f528602fe1312734d734f6326432d7305f30cc30be32ec357c3bca40;
    decBuf[6288] = 256'h9c453e4b084f1a51ba510550774e2c4b5347bc4463423f40a340fd403d434845;
    decBuf[6289] = 256'hac47ec49f74bc34c7c4dd44cd54b7a493a476f43cf3f943b9737ef328d2e6d29;
    decBuf[6290] = 256'hfc25da220220741efc1d691e941fa320f520d6210a21591ff01cc318a313700d;
    decBuf[6291] = 256'h9a07c8005dfa32f668f257f0b7ef25efb2f00cf355f446f6a1f6aaf59ff32bf0;
    decBuf[6292] = 256'hefebd0e69ce0c7dafdd68bd369d0b4ce30cea8cef1cfe2d15cd440d731d9f6da;
    decBuf[6293] = 256'heddb37dc6bdbbbd952d76dd4eed0b3ccb6c820c6d5c28dc129c139c278c4afc7;
    decBuf[6294] = 256'h88cb31d092d48fd82edc88ded1df6ddfa9dd69dbc8d84fd60fd499d2cdd186d2;
    decBuf[6295] = 256'h0fd4a6d6d5d9aedd4ee198e472e811ec7aed9eef01f05cf00af0bfef6bee36ed;
    decBuf[6296] = 256'h1eec1feb37ea0dea33eae1ea3decdfed48f088f293f46ff61ff857f824f8e0f6;
    decBuf[6297] = 256'h10f569f2f0efb0eda5ebd9ea1fea57ea56ebf8ecf1ee55f1f0f266f432f5f4f4;
    decBuf[6298] = 256'h6bf3a0f17eee7feb00e8b5e4b6e1fede39dd43dc8ddc59dd13de9cdf01e1a2e2;
    decBuf[6299] = 256'hbbe3eee31ce4f2e332e3f8e1d1e0dede02dd52dbc9d964d820d7a4d50bd580d4;
    decBuf[6300] = 256'h56d47dd471d5cdd6cbd8a7da4eddc7df07e27de3d1e40fe566e401e3a6e067de;
    decBuf[6301] = 256'h30db32d840d67cd42ad474d4c8d570d89edb9dde55e1cfe36ae5b5e571e5c0e3;
    decBuf[6302] = 256'hc7e163df7fdc8edac9d8d2d788d7ccd700d989daeedbecddc8df79e101e366e4;
    decBuf[6303] = 256'habe5d2e62be8b6e889e9afe98de92ee964e845e7ece54ae4c1e25ce175e0a2df;
    decBuf[6304] = 256'h7cdf59dfb8df0ee090e0d8e019e153e11ee1ede068e0a4dfeddee8ddaedc87db;
    decBuf[6305] = 256'h2dda8cd803d704d61cd59ed411d54bd61ad846dae7dc60dfa0e1abe3ffe4b9e5;
    decBuf[6306] = 256'h61e6c6e7c4e938ed64f298f8c3014d0a4914ff1a192135222f1f991a6e117206;
    decBuf[6307] = 256'h10ffabf502f2e6f0f1f50700cb0e7c2023314540084e64534458ca561450fa49;
    decBuf[6308] = 256'hfe3f99367f30f32aec27012781294b2d1e32c0370e3d42431749e94f5456d55d;
    decBuf[6309] = 256'he564506b7b6f4573f57355737c70d46b3166e360b05a3058ea5539555b58335b;
    decBuf[6310] = 256'hdc5f3e645d696f6b4f6de16d546cfa69d66757640c610e5e555b9159f5578056;
    decBuf[6311] = 256'ha454f3528a50a64d264aeb45cb40f83b5636842fee2ac4267621041e231c4a19;
    decBuf[6312] = 256'hc6185d17ef168c167c1585147a128e0f0f0cd307b30280fcaaf6d8ef6de998e3;
    decBuf[6313] = 256'hc6dc30d8b0d5e6d135d195d027d1b4d20ed557d648d858d9aad9cad866d681d3;
    decBuf[6314] = 256'h3bcf1bca49c5a6bfdcbb6ab88ab6f8b57cb6c7b9a1bd49c2ebc739cdabd0ccd3;
    decBuf[6315] = 256'h82d50fd797d64ed55dd34dd2b2d067d0abd05cd2c5d4a9d729db73de72e1f1e4;
    decBuf[6316] = 256'h3ce815ecb5eff0f310f9e3fdc504310bb112bc17521c7d20c32213227221e120;
    decBuf[6317] = 256'h531fea1d7c1da71e2021f225c52aa8311338e83dba445049d04b924c434da24c;
    decBuf[6318] = 256'h114c7a492047d845e643224287403c40f83f36404e41b34255444e462a48da49;
    decBuf[6319] = 256'h824a4f4a0b499346af42103fe43972361032372fa12c282c962cf92c092e5b2e;
    decBuf[6320] = 256'h102e442d9d2a6f279523e41d9618c313610f420ad006ef043a03b5023d02cf01;
    decBuf[6321] = 256'h6c011101bf00dfff03fe5cfb78f7d9f3aceedae938e4eade17dab5d5dcd24fd1;
    decBuf[6322] = 256'hd7d044d136d3afd593d84cdb10ddacdef6dea2ddfbda63d601d2becbe8c51ec2;
    decBuf[6323] = 256'h4bbd6bbbd9ba5dbbb7bdb6c035c471c86dcc0cd066d2afd3d9d4cad3d3d2c8d0;
    decBuf[6324] = 256'h64ce24cc83c9bfc723c6d9c51dc6cdc717cb61cef1d33fd912de73e270e606e9;
    decBuf[6325] = 256'h7ee911e9e6e76de589e2d0df57dd60dc15dc69dd95dfcbe2a5e64debafefabf3;
    decBuf[6326] = 256'h54f875fb4efedbff63fff5fe04fd8afa02f7b7f3b8f000ee3bece9ebc9eca5ee;
    decBuf[6327] = 256'hd1f007f406f7bef938fcd3fd1efe52fd1dfcb4f974f7d3f4a5f1a6eeb5ecf0ea;
    decBuf[6328] = 256'hfae9afe97beab0eba9ed85ef2cf2f0f38cf56cf628f6f3f4faf20ef08fec44e9;
    decBuf[6329] = 256'h6ae5d4e26be1fde061e170e20ce417e6f3e71fea94eb60ec1aed52ed1fed37ec;
    decBuf[6330] = 256'h64eb0beac6e89fe7f9e5e1e4e2e3fae27be2a2e20ae327e480e522e71be96fea;
    decBuf[6331] = 256'ha4eb4cec7fecf4ebcdeadae876e636e42be24fe01adfe2de15df5ae07de289e4;
    decBuf[6332] = 256'h75e72deaf2eb31ee12ef56ef18ef8fed90ecefea66e967e87fe701e78de6b0e6;
    decBuf[6333] = 256'h51e635e6e6e59fe533e5f8e4c2e4b2e419e5c7e59de6a0e74ee8ece809e9bbe8;
    decBuf[6334] = 256'he5e7e2e663e5fee35ce244e1dfdf53dfd5de62de3fde1fde3cde8bde01dfefdf;
    decBuf[6335] = 256'h0ce165e2aae37ce43ce5ebe5cbe5aee5fde5a3e6e7e79fea73f0f4f708019309;
    decBuf[6336] = 256'h5711621622194d188314ef0cda03dff87df1c7ea8fe9e3ecf7f563037813ee26;
    decBuf[6337] = 256'h0334a944254b1d4d534b73461d3cb832bd275b20a519fb1517171e1ab41e8a24;
    decBuf[6338] = 256'h5c2bc73147395740c246984ce651b856da598f5b0a5bb158d7542f508c4a3e45;
    decBuf[6339] = 256'hcc41ec3fa1413744544a2a50fc56675d3d630767186937678265d960785c5857;
    decBuf[6340] = 256'h8552644f8b4cfe4a854af34a564b1b4db64e964fda4f214fb84c2f49f444b03e;
    decBuf[6341] = 256'hdb3809329e2bc8257a20691e881cf61b7b1cf31c3c1e9f1efa1e031e621b3418;
    decBuf[6342] = 256'h7f13dd0d0b07a000cafaf8f38ded62e998e587e3a6e114e199e111e25ae384e4;
    decBuf[6343] = 256'hdfe48ce4ace3d0e1added4da34d708d236cd93c7c9c358c077bec2bc4fbeb8bf;
    decBuf[6344] = 256'hb7c2fdc61dcc8fcff1d3a6d52ad6b2d58ed30fd0d4cbfbc85bc501c394c2bec3;
    decBuf[6345] = 256'hedc6a1cb44d192d626de36e576ed3af546fab100dc0422077106d105f80259ff;
    decBuf[6346] = 256'h1dfb21f794f51bf51af827fdbb04d40f2a1a3f269e310039b63f5f437b447441;
    decBuf[6347] = 256'hdf3cb4386633932e312a7c2801295b2b342fe634b83bf843bc4bc85033575e5b;
    decBuf[6348] = 256'h205cd05caf59b3550150b34a804455408b3c19397938e7377439ce3bcd3e8541;
    decBuf[6349] = 256'hb444d746024811491b480f461342f43cc036402f3028c521ef1b2518b3141314;
    decBuf[6350] = 256'ha5143b179519b91baa1d051e691c33197f14dc0e0a089f011ffa14f57ef0feed;
    decBuf[6351] = 256'hb8eb07eba8eb16eb9aeb13ec80ec1dec0deb16ea76e7fce473e138dd18d8a6d4;
    decBuf[6352] = 256'h45d048ccb2c949c8dbc73fc84ec9eacaf5ccd1ce81d029d15cd12ed1b3cfe8cd;
    decBuf[6353] = 256'hbccb1bc9a2c607c591c34dc306c48fc526c8a0ca28ce73d196d34fd65ed755d8;
    decBuf[6354] = 256'h0ad8c6d70dd7f5d5c2d5f0d5c3d61cd81ada7edcbede5fe18de4b1e669e9e3eb;
    decBuf[6355] = 256'h22ee2ef00af23ef3e7f34ef3c3f29cf142f0feee2bee51ee8bef03f232f50bf9;
    decBuf[6356] = 256'hb4fd15021206a8082109b308c2064804bf0075fd9bf905f79cf553f4b7f4c6f5;
    decBuf[6357] = 256'h61f76df9d1fb6cfde2feaeffebffb3ff1aff79fd0ffbd0f899f5c0f129efdfeb;
    decBuf[6358] = 256'he0e828e618e522e46ce4c0e5ece7f7e95becf7edd7ee1befe6ededeb89e900e6;
    decBuf[6359] = 256'hb6e2dcde46dcecd9a3d840d89ad891d907dbe3dc93de1ce081e1afe1d9e119e1;
    decBuf[6360] = 256'he0df64de99dcf2d92ed8eed578d4acd3ead392d491d58fd76bd997dba2dd6ede;
    decBuf[6361] = 256'ha3dfdbdf42df5ade34dddadb96da17da57d934d993d95dda7cdb22dd1bdff7e0;
    decBuf[6362] = 256'h23e32ee50ae73fe8e7e880e9f5e8cee775e630e561e3a8e2ffe1cce157e27ee3;
    decBuf[6363] = 256'h8be40be6d6e70ae9b3e94cea7aeafce989e9dae8fde734e748e6aae554e506e5;
    decBuf[6364] = 256'h1de55ee599e516e688e6d2e665e7eee76be8fee8aee984ea87eb35ec13ed69ed;
    decBuf[6365] = 256'h1aed45ec08eb8de98ee819e9e9ea87ee39f48ffc5304670df11545194c1c8c19;
    decBuf[6366] = 256'h0c12f708fcfdb2f0c2e7e3e25de464e85ff39d03c01271241735e63fde41a743;
    decBuf[6367] = 256'hc83e72345d28fe1ca812f20b49082d07330a9f107416ca1ec6287c2f0738933d;
    decBuf[6368] = 256'h9e423447b449764ac649e547e943403f9e395034de30fd2e6c2e02312e36623c;
    decBuf[6369] = 256'he243f64c10539c58a35b8e5cb85b7259a054fd4eaf49dd44bb41e33e553ddd3c;
    decBuf[6370] = 256'h4a3d3c3f6a42694521489b4a924bb14ad5483745863fb4387330af289f21341b;
    decBuf[6371] = 256'h0917c31473151416ec18831bdd1d00209d1f8d1e041bd815a50f25081501aafa;
    decBuf[6372] = 256'hd4f486ef14ec33ea7ee8fae772e804e82fe989e937e9ece820e870e607e423e1;
    decBuf[6373] = 256'ha3dd58da7fd6d6d1b5ceb9ca22c8b9c64cc676c73bc91fccd8ce06d205d5f6d6;
    decBuf[6374] = 256'h51d7fed6f3d47fd144cd47c9b1c657c4eac314c543c8f7cc99d2e7d71bdef0e3;
    decBuf[6375] = 256'hbae78dec6eee46f1d4f23df4abf4d5f530f682f637f6f3f5b5f55ef6c3f77afa;
    decBuf[6376] = 256'h88ffbb05e60ee21938244c306c38ce3fd5439c42103d0036ea2b8522fa19a616;
    decBuf[6377] = 256'h9f133518b61fca283636b842184e6e58245fcd62b161aa5e6956a54e9647553f;
    decBuf[6378] = 256'hc939be342830522f9831aa330b382b3d5e433449824e5553765608577154454f;
    decBuf[6379] = 256'hb1479d3e1236162cb122261ad216d015bb16e51a3320c827d32c932f1332cd2f;
    decBuf[6380] = 256'h5b2c7925381d3c13d6094c0188f97df4e7ef11ef4fee00ef21f2d6f36df6d6f7;
    decBuf[6381] = 256'h1ef9f4f77af5f2f1c6ec92e6bde0ebd97fd3aacd5cc84bc66ac4fcc492c7ddca;
    decBuf[6382] = 256'hb6ce56d2a0d5e9d64cd73dd659d34bce78c9d6c388be16bbf5b763b7f1b84bbb;
    decBuf[6383] = 256'h24bfc4c2f0c7c2cce4cfbcd241d3b9d34cd321d2a8cf0dce01ccadcaf4c92cca;
    decBuf[6384] = 256'h91cbeccd75d1b0d5d0da03e1d9e627ec99efbaf26ff4f4f47bf458f266f0eded;
    decBuf[6385] = 256'h52ec71ebb5eb66edb0f0faf3aff810fd0d01b505d6088c0a190c820d150db10c;
    decBuf[6386] = 256'h570cbc0a4609f2074206b904ba038b035e0404066d08520bd10e1c121a150c17;
    decBuf[6387] = 256'h1b182517af15c312430f080b0c07630242ff8dfdfffb87fbf4fb1ffd98ffd801;
    decBuf[6388] = 256'he303bf05790640064105e7020200bcfbc0f717f3f6ef1ded90eb17ebaaea0deb;
    decBuf[6389] = 256'h1dec13edf4ed38eefaedc2edc3ec7eeb03ea9ee8fde604e528e377e17edf2ade;
    decBuf[6390] = 256'hf5dc4ddc1adc48dcc7dc3adde8dd08deebdd00dda4db03da0ad8b6d681d5d9d4;
    decBuf[6391] = 256'h0cd53ad50dd666d7abd87dd93ddaa6da86da30da4ada03daedd928daf2d9e2d9;
    decBuf[6392] = 256'hd3d9abd9e8d977da27db2ddc67dd8dde9adfd4e0fee0d8e0e4df48dec0dc5bdb;
    decBuf[6393] = 256'h16da98d90bda45db14dd40dfe0e15ae4f5e56be737e875e83de8a4e75fe6e4e4;
    decBuf[6394] = 256'h7fe381e1a5dff4dd4cdd19dd01de25e0c5e2a9e648ea84ee5cf1eaf253f4e6f3;
    decBuf[6395] = 256'h82f3ddf3d3f474f70dfcef025b09300f7e148f16ef15f3112f0a6b0257f9ccf0;
    decBuf[6396] = 256'h78ed7beee6f4bcff060d1b1d3e2c013af04290441643b1392631f22493193d0f;
    decBuf[6397] = 256'h360bfe09520d5d129e1a9a24ff2dfa385c40c2496b4dbf50c653db520552bf4f;
    decBuf[6398] = 256'hed4a4b45fd3f2a3b09387737fb37463bb141f149b551ca5a5463e068e76bfc6a;
    decBuf[6399] = 256'h7c68b2647f5ea958d751414dc14a7b48cb47ac49844c24506e534857d5583f5a;
    decBuf[6400] = 256'hd159e057fc534b4e79470d418d397d323c2ab024aa21bf20ea1f3022a1258227;
    decBuf[6401] = 256'h5b2ae82b702b4d29cd25b01f30182011df081b010cfa76f54bf105ef55eeb4ed;
    decBuf[6402] = 256'h6aeff7f06ff1b8f254f290f0aced2cea00e52de08bda3dd5cbd16acd91cafac7;
    decBuf[6403] = 256'h91c6ffc662c7bdc7fcc908cce4cd94cf1dd150d1c5d04acf19cde2c909c669c2;
    decBuf[6404] = 256'h1fbf20bcf6ba05bc45bea6c248c81acf86d55bdba9e07ce59de82fe9aae841e7;
    decBuf[6405] = 256'h1ee52ce31de226e171e14de3f4e58dea2ff001f76cfdec04fc0b3d14c919d41e;
    decBuf[6406] = 256'h94211524d724262405212c1e961b2d1ae41848190c1b951ec123f42975318438;
    decBuf[6407] = 256'hf03e1b43e5469547f5463f45a9425e3f603ca7399838463826398a3bca3d6a40;
    decBuf[6408] = 256'he4427f44f545c1460846ef448a43e941ef3f133e633cda3a0f395f37d6357134;
    decBuf[6409] = 256'h2d33063246315230742f1e2f332e162d702b97281725dc20df1c3718d513b50e;
    decBuf[6410] = 256'h440b6309ae072907b1064306e0051b04db013bff57fbb8f77cf380efe1eb96e8;
    decBuf[6411] = 256'h72e681e471e37be29ae146e096de9ddcc1da95d8f5d530d4f0d17bd027cff2cd;
    decBuf[6412] = 256'hd9ccdacb4fcb7cca09caa1c942c95fc9adc9f4c935ca21caecc95ac982c87fc7;
    decBuf[6413] = 256'h45c61ec512c4a9c389c319c46dc50ec777c9b7cbc2cdaed0a0d264d400d6e0d6;
    decBuf[6414] = 256'hacd7ead792d82bd913dae6daa5dbdfdc5adebfdf61e15ae336e5e6e6dfe843eb;
    decBuf[6415] = 256'h83ed8eef6af11bf333f4ccf457f581f5a8f585f526f509f523f59af55df67cf7;
    decBuf[6416] = 256'hd6f81afa41fb9afc82fda9fe69ffd2fff1ff9bff4dff05ff99fe10feb7fd24fd;
    decBuf[6417] = 256'h9bfc1efccdfb83fb75fb82fb77fb81fb9cfb94fb8cfb4efbd3fa0efa23f906f8;
    decBuf[6418] = 256'hadf6c5f59ef491f39df2c0f1f7f074f0ceef8def52eff9eea7ee40ee92edbdec;
    decBuf[6419] = 256'h80eb05ea3ae80ee603e4afe27ae162e095e020e1f3e1ffe239e460e5d3e5b0e5;
    decBuf[6420] = 256'hd3e424e373e10adfcadcbfda6bd92dd9f5d88ed9d3da4edcb3ddf7decadff0df;
    decBuf[6421] = 256'hcedfaedfabdeb7dd9adc41dbfcd92ad9b7d894d8f3d882d96eda8adb97dcd1dd;
    decBuf[6422] = 256'hf8de6bdf8edf2fdf9fdee8dd42dd7fdc31dceadba9dbbcdb39dcabdc6bdd56de;
    decBuf[6423] = 256'hf4debddfa9e086e189e2c3e395e455e578e558e502e517e4bbe276e1fbdf96de;
    decBuf[6424] = 256'haedd84dd91de56e0fee22ce606ea9cecf6ee3ef0a2f092eff7ed56eb92e940e9;
    decBuf[6425] = 256'h20ea94edb1f331fb4504d00c5c12671752182714d90e84042efac8f01fedcbe9;
    decBuf[6426] = 256'hd6ee17f7830546135b237e32523caf410f40a13b3b324027f6190611270cad0a;
    decBuf[6427] = 256'h040c8f148b1ef0275d354c3e6b46cd4d254f5d50414f3f4e7f4b54470642943e;
    decBuf[6428] = 256'h733b9a3816387f39583d0142e4482451e858fd6116683269356a74674a63785c;
    decBuf[6429] = 256'h0c568c4e8149c046404402457448954bb5508855a958825b0f5d975c735af456;
    decBuf[6430] = 256'hc851f54c1246a73fd2398434502e252adf272f278f264428da2a342d7d2ea72f;
    decBuf[6431] = 256'h4d2f0d2d41299023be1c5316d20ec2072d0302ffbcfc0bfcacfc3dfdc2fd4afd;
    decBuf[6432] = 256'h01fc10fae1f608f35feefde9dee46ce14ade72dbdbd863d81ad7b7d65cd60ad6;
    decBuf[6433] = 256'h2ad55ed4a5d38cd259d2ced1a4d17dd115d177d074cff4cd29ccfdc9f2c79ec6;
    decBuf[6434] = 256'he5c58dc658c87bcb55cffdd35fd85bdcf2de4be1b9e18ee07fdfe4dd6edc2adc;
    decBuf[6435] = 256'he3dc4ddf31e2e9e418e816eb41ec05eefceedcefb8f157f5fff92202e609fb12;
    decBuf[6436] = 256'h851b492350263b27bb24e91da815e40dd4063e021403de06d30fce1a18289a34;
    decBuf[6437] = 256'hfa3f504a564e8f4f734e6347f84077396832d22d522b902a402b212d1d31bd34;
    decBuf[6438] = 256'hda3aaf40fd45d04af14dca504e51e54fe74cd94745403539f530312925243b23;
    decBuf[6439] = 256'h10245626292b0b3277384c3e1642c7422642073dd336a82d1d25591d4a16de0f;
    decBuf[6440] = 256'h5e0d9c0cec0bcd0da5103c13a5141315af14a01360112a0e500ab1068401b2fc;
    decBuf[6441] = 256'h50f830f3beef5deb60e7cae452e4e4e30fe5d3e66ee8e4e928ea6fe976e78ae4;
    decBuf[6442] = 256'h43e023db51d6afd0e5ccd3ca33cae8cb76cdd0cff3d1e5d3a9d5fcd51bd5c7d3;
    decBuf[6443] = 256'h17d21ed042ce89cdc1cd5acee5ce63cfd6cf3fd05fd0b5d038d1ded1f7d29dd4;
    decBuf[6444] = 256'h96d682d93bdcb4def4e06ae236e3efe327e4f4e322e4a1e414e594e65fe806eb;
    decBuf[6445] = 256'h7fed64f055f21af459f6cff723f94ffb5afd36ffe600ff0164039203c0026601;
    decBuf[6446] = 256'h0bffccfc56fb8afabffb28feb101ec05e809880dd310f612931283119f0e1f0b;
    decBuf[6447] = 256'hd507d6041e020e01bc000701d30107030105dd068d08160a150ba00bca0bf00b;
    decBuf[6448] = 256'h880baa0afb08d805ff0156fdf5f8f8f462f208f09aeffeef77f200f63cfa38fe;
    decBuf[6449] = 256'hce003702ca01d8fff5fb4cf7aaf1d8ea42e66de0a3dc92da32dbc4db5adeb4e0;
    decBuf[6450] = 256'hb3e36be630e826e971e9a5e8f5e68be44ce2abdf31ddf2da51d8d7d53cd431d2;
    decBuf[6451] = 256'hddd09fd0d7d0d6d178d3e1d5c5d87edb8ddc84dda4dcc8da21d8f2d4f4d13bcf;
    decBuf[6452] = 256'h77cddbcb26ccf2cca2ce0cd14bd3c1d48dd5cbd523d58ad4a2d37bd221d1ddcf;
    decBuf[6453] = 256'hb6ce43ce66ce85ce4fcf3ad056d163d228d4d9d561d72cd9e6d98edac1da36da;
    decBuf[6454] = 256'h0cdae5d9c3d9e2d9ffd919da60daa1da2bdb13dcaedd17e045e464e9f9f00dfa;
    decBuf[6455] = 256'h97025b0a670f2712a70f590a640169f613ecade204dfe8ddf3e2dfee7efd2f0f;
    decBuf[6456] = 256'h9724fb32104070429a44b43e32329323d0154e096e0400000704210a5516b421;
    decBuf[6457] = 256'hf231c13c9646854f2551ab4f534e394875406639fa32d02e062bf428d52ad12e;
    decBuf[6458] = 256'h8334d93c9d44b14d3c56c85bcf5e8f610f5f455b1155914d8146403eec3ae637;
    decBuf[6459] = 256'hfb36d0379a3b6d400f465d4bcf4ef0518252f550aa4dd0491f444d3de2360c31;
    decBuf[6460] = 256'h3a2aa4257921af1d9e1b3f1cd01c5e1eb8200022f2234c2455231f20461c9416;
    decBuf[6461] = 256'h4611130b3d05efff7dfc5cf9a7f722f7aaf617f77bf720f7cef658f5f4f2b5f0;
    decBuf[6462] = 256'h7eed80eac7e74ee50ee303e1afdfffdd76dcabda7fd874d620d5ebd3d2d29fd2;
    decBuf[6463] = 256'hced2a0d3fad43ed665d7d8d7fbd75dd721d652d426d21bd0b7cd1bcc3bcb7fcb;
    decBuf[6464] = 256'h2fcd99cf7dd2c3d6c0da5fde9be273e50ae873e9bbea1febc4ea72ea92e94ee9;
    decBuf[6465] = 256'h10e9b9e9eaeb20efd4f377f94900b406890cd711aa16cb195d1ad9196f187115;
    decBuf[6466] = 256'hb812f410fd0fdd10c9134917661d3b230d2a7930a434f239033ca33cee3a6039;
    decBuf[6467] = 256'h063708341632523000304a30263249352339c23cfd40fa449047ea49584af449;
    decBuf[6468] = 256'h3048f045ba42e03e4a3cff38db36b135a134f434d43528375d3875390e3a3d3a;
    decBuf[6469] = 256'h6a39c4375b35d231962d9a29f2249020941cfd19a3175b16f715e81496144b14;
    decBuf[6470] = 256'hf7124711dd0e540b19071d0374fe13fa16f680f326f102ef9fee44eef2eda7ed;
    decBuf[6471] = 256'h53eca3ea3ae856e50fe113dd73d938d55fd2c9cf6fcd26ccfcca56cb04cbe4cb;
    decBuf[6472] = 256'ha0cb5acc92ccc5cc50cd7acd54cda5ccc8cb8cca10c945c711c688c489c3a1c2;
    decBuf[6473] = 256'hcbc23ec332c4cdc556c721c9d2ca5accbfcd04cf2bd038d171d244d39dd4e2d5;
    decBuf[6474] = 256'h09d762d8a7d9ceda27dc6cdde7de18e123e387e5c7e768eae1ecc5efb7f130f4;
    decBuf[6475] = 256'hccf5d7f72bf9e4f9fdfa30fb5efb34fbc1fae4fa43fb45fc0bfeb200e103ba07;
    decBuf[6476] = 256'h5a0ba40ec810b912c9131b143b135f11ae0f260ef50b7f0a2b09f607be07f107;
    decBuf[6477] = 256'hd908540a1f0c4b0e5610321267130f14dc1397122010f10cf309730628032a00;
    decBuf[6478] = 256'h38fe29fdd7fc21fdedfd9eff27018c0273039e037703c902ac01530055fe69fb;
    decBuf[6479] = 256'hb0f882f583f2cbef9cec79ea4ee93fe891e871e93dea72eb8bec24ed98ecc6eb;
    decBuf[6480] = 256'h20eab6e777e5d6e25ce078dd87db0dd916d836d76ad6a8d650d74fd837d95eda;
    decBuf[6481] = 256'h1edbccdbecdbcfdb81dbabdaa8d96ed8f3d628d578d3efd124d06bcf52ce85ce;
    decBuf[6482] = 256'h10cfe3cf89d112d3ddd48dd6a6d73fd810d892d739d697d40ed3a9d165d03bd0;
    decBuf[6483] = 256'haed0e8d1b7d3e3d584d848da88dcfeddcade8cde54de21de39ddbadc47dc24dc;
    decBuf[6484] = 256'h83dc13ddfedd99df92e16ee316e6dae71aeafaea3eeb00eb58ea25ea53eacfeb;
    decBuf[6485] = 256'hccee80f322f9f4ff3508c10dcc12b713e212940d6007e0ffd0f865f2e5ef2bf2;
    decBuf[6486] = 256'h5ef88901f50e781b172aeb334839e73a6d39b7322d2a31207b19611345124b15;
    decBuf[6487] = 256'he1196221762a7135d33c8943c244de45e0462044f53f2b3c1a3af8364335bf34;
    decBuf[6488] = 256'h28367037293a0c3eb5421747364ca84f0a54bf553b55d253f84f504b6d44023e;
    decBuf[6489] = 256'hd7390d365c35fd35d5387e3de041ff46714a924d014d734b194965440340e33a;
    decBuf[6490] = 256'h1136af31d62e402ce6299d28732763266d258c2448240b24d2233923ae22df20;
    decBuf[6491] = 256'hb31ee71a48171c12490de708c803b70195fee0fc65fdddfd6ffdd3fd78fd39fb;
    decBuf[6492] = 256'h98f8b4f40cf0aaebaee717e5bee275e1d9e133e2e1e12ce260e134df93dc65d9;
    decBuf[6493] = 256'h66d6aed3e9d197d177d2cbd3f7d502d8ded913dbdbdadcd9ded77ad595d2a4d0;
    decBuf[6494] = 256'hdfce8dced8ce2cd058d28ed58cd80cdc56df55e20de53ce85fea8aeb4eed45ee;
    decBuf[6495] = 256'h90ee4cee0eeed6ed3ded0fed39ed92ee34f09df226f670f925fe8702a607da0d;
    decBuf[6496] = 256'haf13fd18311f0625d028e12a822ba9280925ed1e1719c913b8111811f013ab1a;
    decBuf[6497] = 256'hc124d630353c8b46f04f0a5626572456b94f3848243f9936d52eca290a278a29;
    decBuf[6498] = 256'h542d8733083b1c44364afa510155c157eb56a554724ef246e23fa137dd2fcd28;
    decBuf[6499] = 256'h0d268d234f24c127232c66323c38063c173e763d9e3af535122fd2260e1ffe17;
    decBuf[6500] = 256'h9311bd0b77096607c6063406c1072b09730ad70a310b3a0a2f084305c40197fc;
    decBuf[6501] = 256'hc5f723f2d5ec02e860e212dda0d97fd6c9d43cd3b4d3fdd427d6ecd7e2d898d8;
    decBuf[6502] = 256'h44d718d5e2d108ce69ca1ec745c3aec045bffcbd99bda8befbbe70c03cc1f6c1;
    decBuf[6503] = 256'h9ec2d1c2a3c279c252c275c252c3e2c3cdc4abc53ac620c6aac5e7c464c41dc4;
    decBuf[6504] = 256'hb4c4dbc553c8ebcc4dd149d5f2d953de2ce1bae223e4b5e352e342e2f0e110e1;
    decBuf[6505] = 256'h54e189e282e46ee7edea29ef25f3c4f60ffa0dfdc6ff8a0126039b0467052106;
    decBuf[6506] = 256'h590626069b057105fd0466054306b907ea09200d1f109e13e9160d19371a921a;
    decBuf[6507] = 256'h9b199017b4150c134811ad0f370ef30d310ed90e3e1083115512621310143014;
    decBuf[6508] = 256'h13149013ea12d111c410450f7a0dca0b600920071505390304025c012901fb00;
    decBuf[6509] = 256'h79019f013701d80062ff31fd26fb3af881f508f36df161ef0dee54ed3ceca3eb;
    decBuf[6510] = 256'hbbeae8e9dbe85ce7f7e555e4cde202e1cddf44dedfdc3edbb5d950d80bd738d6;
    decBuf[6511] = 256'hdfd4f7d3d0d210d262d1c4d034d01ad0d3cfbdcff8cf51d0c3d02ad102d17dd0;
    decBuf[6512] = 256'h95cff9cd00cc24ca74c85bc728c7b4c72fc960cb00ce2fd152d344d59ed54cd5;
    decBuf[6513] = 256'hd6d3fad153cfdacc3ecbc9c985c935cb2ecda2d0edd3c6d766dbc0ddbee0e9e1;
    decBuf[6514] = 256'h8ee13ce1c6dfeaddbedbdeda9adad8da61dc92de32e161e45fe718ea91ecd1ee;
    decBuf[6515] = 256'h72f1ebf3d0f616fb360009056a09430cd10d670c69095b0428fea8f6a1f3e1f0;
    decBuf[6516] = 256'h61f3b7fbb305c7116620292e1937f83b723d6b39e130ad244e19ec11350bfd09;
    decBuf[6517] = 256'h510d65166121b72bcb37eb3f4d47544b1b4ac746bc41263d513787337531d530;
    decBuf[6518] = 256'h6731f4323f36193ac13e63442d48004d62511753a4542c540952894e4e4a5146;
    decBuf[6519] = 256'hb242673f1f3ebb3d803fc04160448f47b249a44bfe4b634a58486c45b342853f;
    decBuf[6520] = 256'h613d703bab396c37f6351a34ee31e32f7f2d3f2b9e288f279826b8257425bb24;
    decBuf[6521] = 256'h32230121601e7c1add169213b90f220dd809b4078a062f063805c3036f024300;
    decBuf[6522] = 256'ha2fd29fb44f8c5f46bf26def42ee7eec87eb3ceb70ea3be9b2e71be5ede1eede;
    decBuf[6523] = 256'h36dcbcd921d8abd6efd624d81dda81dcc1de37e003e14ae031df9adc6bd992d5;
    decBuf[6524] = 256'hfbd2b1cf68ce05cec9cfaed22dd668da65de0de32ee607e995ea0deba0ea3cea;
    decBuf[6525] = 256'h2de936e8ebe71fe75de705e8d0e977eca6ef5af4fdf94bff7e05a909f70e0811;
    decBuf[6526] = 256'he9127b13ed118410600e360d260c790c840ef8113316531b86215c27262bf92f;
    decBuf[6527] = 256'hd9316b32e7316e312630fb2eec2d9a2d7a2ece2f7e31e733cc368439493be43c;
    decBuf[6528] = 256'h5a3e163ed83dbf3c5a3b5c3908385836b0357d35ab3529369c360537a6361636;
    decBuf[6529] = 256'hc33421332831c42e852c792a15287a260425b0230022e7201c1f6c1de31b7e1a;
    decBuf[6530] = 256'h8018a41678146d120910250d6c0a3e073f04c00075fd77fa85f8c1f6caf5eaf4;
    decBuf[6531] = 256'ha6f4edf3d4f26ff171ef0ded84e939e660e2c0de76db52d928d818d7c6d67bd6;
    decBuf[6532] = 256'hbfd682d649d616d62fd508d4fbd2c1d19ad041cf59ce86cdc7cc5eccffcba9cb;
    decBuf[6533] = 256'hc3cbabcb96cb82cb94cbc5cb2cccbfcc97cd9ace8ecfaad004d248d36fd4c9d5;
    decBuf[6534] = 256'h0dd734d841d935da51db5edc98dd13df78e019e213e4efe51ae890e96ceba1ec;
    decBuf[6535] = 256'h2aee29ef11f037f1f7f1ebf208f461f5a6f6cdf773f98cfa57fc8bfd14ff7900;
    decBuf[6536] = 256'h1b02a4036f059a071009ec0a9c0c450dde0d690eea0dc40d5b0dfd0ce00c620d;
    decBuf[6537] = 256'h090ef70e131020111412f1120e13c01249125b113e10320f3e0e210dae0c000c;
    decBuf[6538] = 256'ha10b840b360bbf0a270a2809ee07c8066e05cd03b402b50171004aff3dfebdfc;
    decBuf[6539] = 256'h58fb5af97ef753f5b2f238f09dee92ec3eeb09ea61e9c8e83de812e853e75ee6;
    decBuf[6540] = 256'h03e5a8e268e032dd0edb56d891d6f6d4abd4efd42dd5d5d508d637d6b8d55fd4;
    decBuf[6541] = 256'h61d2fdcfbdcd1ccba3c808c727c66bc625c73dc86eca79ccddce79d059d115d1;
    decBuf[6542] = 256'h5cd0d3ce3cccc2c983c777c523c4e6c38ec459c685c825cb54ce52d10bd4cfd5;
    decBuf[6543] = 256'hc6d611d7cdd698d580d481d3f5d2cbd28bd3c5d494d6c0d861dbdadd1ae025e2;
    decBuf[6544] = 256'h01e436e54fe64ee7d9e7afe73ce748e62be51ee470e350e3e0e368e5d1e7b6ea;
    decBuf[6545] = 256'h35ee70f26df60cfa66fcaffdd9fe7ffe88fd3dfdf9fc2efeb7ffb4028d062409;
    decBuf[6546] = 256'h7e0bc60c630ce909050785032b0199018a03d808aa0fc0192623b02b3c313e32;
    decBuf[6547] = 256'h2933542d82261620eb16d110b50fb30e4913c91add23682c64361a3dc3401744;
    decBuf[6548] = 256'h1141503e253ad7340530a32bee296929e229052c852fc033bc376e3d38410a46;
    decBuf[6549] = 256'h2c49e14a654bfc49fe467e43433f233ab1369033fe328333ec34c538653ca040;
    decBuf[6550] = 256'h9d4433479c480a4918479f447140753cd6388b358d329b30d72ee02d952dc92c;
    decBuf[6551] = 256'h942bec2a872942281b270f26d524ae235522b320ba1e561ccd188315a9110a0e;
    decBuf[6552] = 256'hbf0a9c08aa06e60493044904050442040a0471032d025d0032fe91fb17f9d8f6;
    decBuf[6553] = 256'h37f472f2d7f0cceef0ec40ebd6e8f2e500e487e190e045e089e03ae2a3e487e7;
    decBuf[6554] = 256'h79e93deb90ebafea4be8c3e487e08bdcebd892d649d5add526d8afdbeadfe6e3;
    decBuf[6555] = 256'h8fe8b0eb89ee0def86ef18efeeeddeece8eb32ecfeec33eebcefedf18ef452f6;
    decBuf[6556] = 256'h36f9effb1dff1c029b05e608c00c5f10aa13a816d317e2189018b017e416a616;
    decBuf[6557] = 256'h6e1607170519691bf21e2d230626a529f02c132f3e3098304630fb2f3f300230;
    decBuf[6558] = 256'h3a30d3300131d730b1300230642f612eb32d542daa2d612ec62f2b316f32ea33;
    decBuf[6559] = 256'h8334b2343334da3239313f2fdb2c402b35295927a9252024bb2276214f20431f;
    decBuf[6560] = 256'h4f1eb01dae1cff1b221b1f1ae518be177f153f1309100a0d8b09400642038900;
    decBuf[6561] = 256'h10fed0fbc5f9f9f8c4f71cf7e9f65df68bf5cbf44bf380f1d9eeabebace866e4;
    decBuf[6562] = 256'h8de1eddd93db70d945d8ebd799d7e3d727d865d89dd8d0d8a2d824d8b0d748d7;
    decBuf[6563] = 256'he9d659d6a2d59dd4a9d38cd280d1d1d072d056d0d8d0ded15dd328d554d75fd9;
    decBuf[6564] = 256'h3bdbebdc04de9ddecbdea1de2edec6dda6dd50dd9edd74deb0df7fe1abe3b6e5;
    decBuf[6565] = 256'ha2e85bebd4edb9f071f336f5d1f647f88bf844f97cf949f9d4f953fac6fa00fc;
    decBuf[6566] = 256'h7bfd46fff6005f039f054008040a440c4f0ea30fd810f1118a12b812e212bc12;
    decBuf[6567] = 256'h53127611e610fb0f1e0f540e060ebf0dd40d360e900e430fb90ffa0f0e10b40f;
    decBuf[6568] = 256'hc10e410d760b4a09aa063004f00150ff8bfdf0fb10fb44fa8af952f9b9f82ef8;
    decBuf[6569] = 256'hb0f7a3f669f5eef323f2f7efeced88eba4e8ebe5bde299e0e1dd1cdc81da36da;
    decBuf[6570] = 256'hf2d9acda54dbeddb78dcf6dcd0dc96dbc7d920d73cd39dcf52cc78c8e2c588c3;
    decBuf[6571] = 256'h40c2a3c2b3c3a9c4b5c609c83dc956ca89ca5bcadcc9d0c850c7ebc54ac4c1c2;
    decBuf[6572] = 256'h5cc174c04ac00ac1fec199c392c5f6c736ca41cc95cd4ecef7cec4ce95ce17ce;
    decBuf[6573] = 256'ha4cd81cda0cd30ce1bcf77d019d212d4eed59ed727d98cdad0db4cddb1de52e0;
    decBuf[6574] = 256'hdbe10ce482e55ee70ee926ea25ebb1ebdbeb4eecb6ec15eddfedfeee0bf0d0f1;
    decBuf[6575] = 256'h80f3eaf5cef886fb00fee400d6024f0546062607f2073008d8083d0a3b0c9f0e;
    decBuf[6576] = 256'h28126316601af61c501fbe1f931e1a1c911837161314b0137415461a7a20fa27;
    decBuf[6577] = 256'h0a2f75354b3b0d3c5c3bfa36b730e22a10247a1fa41e661f3924db29ad301937;
    decBuf[6578] = 256'hee3cb840c9426a43b4411e3fe23a0a3873351933d1316d3113310a321534f135;
    decBuf[6579] = 256'h1439123c923fdc42db45054760476946c8439a40e53b8337ab341432ab301931;
    decBuf[6580] = 256'h0a3339363739f03b693e0440ba3fde3db23b7c38a2340c32c12e9d2cac2ae728;
    decBuf[6581] = 256'h4c27d62582245722e120051fd01d281d291cfa1bd01b101b1c1a8118a815ef12;
    decBuf[6582] = 256'h0c0f630a0106290389ff2ffdc2fc5efcb9fc0bfdebfda7fd69fd70fb0cf928f6;
    decBuf[6583] = 256'h70f341f043ed8aeac6e8cfe759e68de558e4cfe26ae16cdf90dd5cdc43dbaada;
    decBuf[6584] = 256'h35db08dcaedd37df36e01ee1f3e0e7df67de36dc95d91cd725d645d589d539d7;
    decBuf[6585] = 256'ha3d987dc06e060e25fe589e64ee844e98fe95bea90eb38ec37ed7ceea3ef63f0;
    decBuf[6586] = 256'h11f170f1c6f1b1f24cf4b6f63ffa7afebd04930ae10f5313b4174618c2175916;
    decBuf[6587] = 256'h5a13a210730d2b0c8e0c530edb1107173b1d1023da26ad2bce2e8430ff2f872f;
    decBuf[6588] = 256'h632d392c742a7d293329ef28a829502a4f2bf12c7a2edf2f803109330834f034;
    decBuf[6589] = 256'hc235e9358035a3342d33c831ca2f762e412d282c8f2bbe2b942bba2b972bf92a;
    decBuf[6590] = 256'hf6297728ac268024df211b20db1d651c111bdc19c4185f171a169f146e126310;
    decBuf[6591] = 256'h770dbe0a90079104a00226008bfeabfd57fc9efbf5fa90f94cf828f687f30ef1;
    decBuf[6592] = 256'h85ed3aea3ce783e40ae2cadfbfdd6bdcb2db09dbd6daa8da7eda57daefd951d9;
    decBuf[6593] = 256'hc1d80ad805d7cbd550d4ebd249d1c0cfc1ce36ce0cceccce06d0d5d101d4a2d6;
    decBuf[6594] = 256'h66d802dae2da9eda60dab8d953d86bd741d71ad783d7dfd880daeadccedfbfe1;
    decBuf[6595] = 256'heee411e703e9c7ea63ec43ed87ed40eee8eee7efcff0a2f148f3d1f49cf64cf8;
    decBuf[6596] = 256'h45fa21fcd2fdeafee9ffd1004f017601de013d0294027f039b04f50596071f09;
    decBuf[6597] = 256'h1e0a060b300b0a0b5b0a7e097b088707e90620069d05850544050905f804a604;
    decBuf[6598] = 256'h3f04e1032c0375029f019c00a8ff4cfeabfcb2fad6f8aaf69ff4c3f212f1faef;
    decBuf[6599] = 256'h61efd6eeacee85ee1dee7eed42ec73ea47e8a6e52de3ede077df23dee6dd1ede;
    decBuf[6600] = 256'h51de7fde55dee2ddeedcd1db78dad6d8bed759d614d541d482d3d3d2f6d12dd1;
    decBuf[6601] = 256'h41d0e3cf8ccf72cf18d085d00ed1afd1c4d1b1d134d160d05ecf6ace8ccd36cd;
    decBuf[6602] = 256'h84cd2bce6fcfb4d0dad1e7d295d3b5d3d2d383d36cd381d30bd417d5bdd6b6d8;
    decBuf[6603] = 256'h92da42dc5bdd5ade42dfc0df33e09ce03ae1cae1b5e2d2e3dee418e63fe74ce8;
    decBuf[6604] = 256'hcbe930ebd2eccbeea7f0dbf164f363f4eef46df52df621f73df897f938fb31fd;
    decBuf[6605] = 256'h95ff31011102dd021b035303ba028b02b502750369040506fe07da098a0b130d;
    decBuf[6606] = 256'h780e600f32103f110413b5148e17471ac01c5b1ea61e521dab1a7c17c812a70f;
    decBuf[6607] = 256'hf10d6d0db8104716191d5a251e2d2e34ee36c3377d354a2fc927ba2079182515;
    decBuf[6608] = 256'h1e1209133417821c1624262b9131bc350238b238d136f93359301e2c22288b25;
    decBuf[6609] = 256'h3123e921be20ce2169230a26ed298d2dd730b1344737b03843381837ea331030;
    decBuf[6610] = 256'h712c36283924ac223322a1225925d3275c2ba62eca30f4319a31a330982eac2b;
    decBuf[6611] = 256'hf328c525a123e920d91fe31e021ebe1d051d5d1c5e1b191a9e189f175a168815;
    decBuf[6612] = 256'hc8145f148213f2129e11fd0f040ea00bbc0803068a03a5007bffb6fdc0fc75fc;
    decBuf[6613] = 256'h31fc6ffc37fc38fb50fa29f983f7faf52ff47ff266f101f0bcee95ed3cec9bea;
    decBuf[6614] = 256'h12e9ade70be6f3e45ae488e45be501e78ae8efe933ebb2eb8beb97eabde859e6;
    decBuf[6615] = 256'h19e478e1b4df19de63de2fdfd7e105e504e883ebceeeccf1f7f206f459f40ef4;
    decBuf[6616] = 256'hcaf395f2edf154f125f14ff1c3f171f2cdf328f667f833fcd3ff0e040a08aa0b;
    decBuf[6617] = 256'hf40e18114212e811f110e60e0a0dde0afe09ba09ef0a580de1101c153c1a0f1f;
    decBuf[6618] = 256'h70234926d7274029d228a827e3254824d2227e21c5201d20b6209d211923e424;
    decBuf[6619] = 256'h0f271b29f72aa72c4f2d4e2e202ea12de22ca82b2d2ac82883270826a3245e23;
    decBuf[6620] = 256'h8c22cc211d21fe201a2135217c21bd21822128215520df1e141de91add187916;
    decBuf[6621] = 256'h3a149911d40f390ec30cf70bc30aaa09ab08c3079c064305fe03d7027e013900;
    decBuf[6622] = 256'h13ffb9fd18fc1ffa43f89bf522f3e2f041ee7dece2ea01eabde980e928ea5bea;
    decBuf[6623] = 256'he6ea10eb9dea35ea18e9bfe71de694e4c9e295e10ce073df44df1adf8ddf81e0;
    decBuf[6624] = 256'h5fe128e213e3f1e380e403e51be55ce596e585e595e5a4e596e5d3e520e67ae6;
    decBuf[6625] = 256'h17e7dae791e867e969ea5eeb7aecd4ed18ef3ff098f180f253f313f4c1f420f5;
    decBuf[6626] = 256'h76f5f9f59ff662f781f8dbf91ffb9afcfffd44ff1700d6008501a40188013901;
    decBuf[6627] = 256'hc3002b00a2ff25ffd3fec5feedfe42ffe7ffbc00bf016e020c032803da02d501;
    decBuf[6628] = 256'h9b00ccfe1bfd22fb46f91af7a5f5d9f41ff4e7f3b4f386f3b0f38af321f3c2f2;
    decBuf[6629] = 256'hf9f1daf080ef3cee6cec40ea35e859e6a9e420e3bbe130e1b2e08be023e042e0;
    decBuf[6630] = 256'h5fe045e05de047e0e5df8bdfd9de03de00dd81dbb6d905d80cd6b8d483d3dbd2;
    decBuf[6631] = 256'h74d35cd42bd657d862dab6dbebdc23dd8adc46db76d9c6d73dd63ed5b3d431d5;
    decBuf[6632] = 256'h3ed603d8b4d91ddcb8ddc3df8fe049e111e144e1b8e08ee0b5e0d8e076e13fe2;
    decBuf[6633] = 256'h2ae347e4ede576e7a7e91cebf8ec2deed6ee09efdaee5cee9ced33ed53ede3ed;
    decBuf[6634] = 256'h6bef64f1c8f307f6a8f8b8f9aefaf9fab5fa80f968f8cff744f7c2f7cff894fa;
    decBuf[6635] = 256'h44fc3dfe1900ca0172020b03dd025e023802cf01b001cc01e701cf01b9015701;
    decBuf[6636] = 256'hfe00cd00f900c201380369057407d809180cf80c3c0d070c7e0a4d08d7068305;
    decBuf[6637] = 256'h3d06c607c30ac10d41119a130814dd12af0fd50b3608dc059404be05ed087c0e;
    decBuf[6638] = 256'hca13fd19281e6e205d1e3c1b1c16e90f130a49063804d804b1075a0c3c13d217;
    decBuf[6639] = 256'ha81dee1fff215f21a91f1c1ec21b9e19ad1752170017b516f916b317cb18301a;
    decBuf[6640] = 256'h2e1c921e77212f24a926e8285e2aa22a642adc28ab269f24c3228f21c7216022;
    decBuf[6641] = 256'h01246a26aa284b2b0f2d622dac2de02c302b37295b27ab259224f923cb23a123;
    decBuf[6642] = 256'h14247c249c24b92436249023cd22ae21a120671f411e341dfa1bd31ac719d218;
    decBuf[6643] = 256'h771732160b156513dc111110dc0ec40dc50c800bad0a3a0a460969086607e605;
    decBuf[6644] = 256'h1b04f001e4ff80fde5fbdaf9fef7c9f6b1f5b2f426f4a8f3e8f23af29cf1d2f0;
    decBuf[6645] = 256'h50f0d9ef98ef85ef73ef42efdbee12eed6ec5beb90e9dfe757e6bee5ece567e7;
    decBuf[6646] = 256'hfee92ded2bf0abf304f672f6d5f67bf6e0f46af316f25df195f194f292f47ef7;
    decBuf[6647] = 256'h36fab0fc4bfec1ff1501ce01060205034a04c5059007370ab10cf10e66103211;
    decBuf[6648] = 256'hec11b31180115211d01190121014db150718a71a6c1c071e7d1fc11fff1f3720;
    decBuf[6649] = 256'h6a203b2066208c20f5205321e3216622ad22ee22da22ec22dc22eb2213234f23;
    decBuf[6650] = 256'h8623e0230524e4239e231523ef21c8206e1f2a1e031df61b481baa1a1a1a9719;
    decBuf[6651] = 256'h801913198a180d183a1737164315e713a212d310a70e060c8d094d0742056603;
    decBuf[6652] = 256'h31021901e6005a0030000a00a1ff03ff00fec7fc4bfb80f955f749f56df3c6f0;
    decBuf[6653] = 256'h4deeb1eca6eadae921e959e98ce974ea47eb06ecb5ec95eccceb78ea7ae816e6;
    decBuf[6654] = 256'hd6e361e20de1cfe007e1a0e188e25be367e4d0e42fe54be531e51ae52fe5b9e5;
    decBuf[6655] = 256'ha1e6bee7cae8bee91dea00eab2e90ce91ee880e72ae70fe7b6e7cfe875ea6eec;
    decBuf[6656] = 256'hd2ee12f11df3f9f42ef646f745f8d1f84ff975f952f972f955f93bf923f939f9;
    decBuf[6657] = 256'h4df9a6f99afad4fba3fd53ff4c0128035d049504fc031403450195ff9cfd48fc;
    decBuf[6658] = 256'h0afc42fcdbfc7cfe95fffa0085015b014e00cffe9efc93fab7f806f7eef5bbf5;
    decBuf[6659] = 256'he9f513f686f6eff6cff606f61bf5bff3c1f16df041eecbecffebcbea22eaefe9;
    decBuf[6660] = 256'h64e93ae914e9f1e892e83ce851e734e627e5a8e3dde1a8e01fdf20de38ddbadc;
    decBuf[6661] = 256'h47dc24dc04dce7dbcddb86db70db84db72dba3dbeddbdfdbbbdb84dbeeda2bda;
    decBuf[6662] = 256'h74d99fd848d82ed876d863d980da8ddb81dc5eddeedd3cde84de99defbde78df;
    decBuf[6663] = 256'hcadf4ee0a8e0d9e022e180e1d5e14ee221e324e4a3e56ee79ae9a5eb81edb6ee;
    decBuf[6664] = 256'h5fef2ceffdeed3eeadee8aeea9ee00ef82ef88f07cf198f2a5f353f4f1f4bbf5;
    decBuf[6665] = 256'h0ef70cf9e8fa14fd8afe56ff18ff70fe71fd2cfc05fbf9f94af9a9f9acfab7fc;
    decBuf[6666] = 256'hc2fe9e004f0267039a03c9034a03d70229024b01bc0039002100e400cf012b03;
    decBuf[6667] = 256'h6f049605f006340807092d09c508a8070206e904ea035f0332043e0578064808;
    decBuf[6668] = 256'h7c09950a2e0ba30a28095d073105bb03ff03b0051908a20bdd0fb6125516be17;
    decBuf[6669] = 256'h2c183a160c13570ef6091d078f0508062b08ab0be60fe2138b18ed1ca21e2f20;
    decBuf[6670] = 256'hb71f6f1e7d1c6e1bc01b0b1cd71c901d191f18205c21d722d62362248c244c25;
    decBuf[6671] = 256'h40261a287e2abe2c342e782ebe2da62c412bfc2929296a2801289f28152a462c;
    decBuf[6672] = 256'he72eab30a231c230f62f452ebc2cbd2b792afa29ee2885286628bc280a292229;
    decBuf[6673] = 256'h342899261025452310226821cf20e71fc01e1a1d011c021b1b1af4189a179c15;
    decBuf[6674] = 256'hc0131012f710920faa0e2f0d640bb4092b082c07a106230616059603cb019700;
    decBuf[6675] = 256'h7eff7ffe3afd14fcd4f994f71ef6caf496f37df2e4f1b6f1e0f139f337f59bf7;
    decBuf[6676] = 256'h37f917fad3f99ef8c4f50cf328ef89eb3ee81be6b7e57ce705eb31f064f68ffa;
    decBuf[6677] = 256'h59fe6a000a0155ffc8fd6efb94f7fef495f302f42df5a6f7e6f987fc00ff4001;
    decBuf[6678] = 256'he1035a069a08100aec0b200dc90d620e900e660ea60db20c950b220b8b0b260d;
    decBuf[6679] = 256'h8f0f181363163c1ad31c1d20662190228121411fa01c271a8c18ab17ef172419;
    decBuf[6680] = 256'had1ade1c7f1ff821dc2407261627c4264e25fa234a22c120f61e461d4d1b7119;
    decBuf[6681] = 256'hb8180f18a81833195a1a1a1bc91b271c441cc21b5d1a2c188c151213d210c70e;
    decBuf[6682] = 256'h730d3e0cb50aea083a07b1054c0408038d01c2ff8dfe74fddbfcadfc83fc76fb;
    decBuf[6683] = 256'hf6f92bf884f50bf36ff1cfee0aed6feb64e910e8d2e72ae7f7e66be645e538e4;
    decBuf[6684] = 256'hfee2d7e164e141e122e105e1b6e040e0a8dfd0de5bdd90db64d959d705d64bd5;
    decBuf[6685] = 256'h13d5acd594d60fd874d916db9fdc04de8fdeb9def9dd79dc14db2cda06d9dfd8;
    decBuf[6686] = 256'h02d9a0d9a3da23dceedd9edf07e2a2e3aee502e736e8dfe878e9a6e928e9b5e8;
    decBuf[6687] = 256'h06e868e74be731e7d8e71ce9bdea27ed66ef07f281f4c0f6a1f7e5f722f87af7;
    decBuf[6688] = 256'he1f6b3f6e0f56df504f5e5f401f584f52af618f735f8f5f8a3f9c0fa80fbb9fc;
    decBuf[6689] = 256'he0fdedfe9bffbbff2bff40fea5fcacfa48f808f692f4c6f304f41df582f623f8;
    decBuf[6690] = 256'hacf9abfa36fb0cfb99faeaf98ff8edf6f4f418f3e3f1cbf098f0c6f0f0f017f1;
    decBuf[6691] = 256'h39f159f13cf1eef018f0a2eed7ecacea36e9e2e729e7f1e6bee649e7c7e720e9;
    decBuf[6692] = 256'h65ea34eceeec96edfdec15ec46ea96e80de742e591e309e2d6e104e22be31ee5;
    decBuf[6693] = 256'hfae6aae833ea32eb1aecececacedcfed70ede0ec2aecb3eb72eb10ebb6ea24ea;
    decBuf[6694] = 256'he9e91fead2ea36ec01ee2df0a2f1f6f22bf444f543f62bf7a9f783f760f701f7;
    decBuf[6695] = 256'he4f6fef646f7b2f714f86df8dff846f9a4f9c8f97bf90df9a6f899f84ef9a2fa;
    decBuf[6696] = 256'h43fcccfd31ff76004901bc019901fb00beff43fe78fcc8fa20fa87f9b5f9dff9;
    decBuf[6697] = 256'h52fa01fbdefb54fd1fffcf00c8021c045105f9052c06fe052b0538034c0094fd;
    decBuf[6698] = 256'h1afb24fad9f9b5fbe1fd170115049507ef09370bd40ac40929081e06ca048c04;
    decBuf[6699] = 256'h1506e007870ab60db410a612b51307142713d31123102a0e5e0d9c0db40e7f10;
    decBuf[6700] = 256'hab124c157a18791b311e60218323ae24bd256b258b2437230b21001f241def1b;
    decBuf[6701] = 256'h471be01bde1dca2010250c29b52dd630af333c35c4347c33fc2fb12cb3293326;
    decBuf[6702] = 256'hca245d24c024852620289629722ba72c4f2d822df72c782cb92bc42a69292428;
    decBuf[6703] = 256'h5526202507246e23e322b9229322e42185212f21ac2036201d1f761d7d1ba119;
    decBuf[6704] = 256'h76170016ac147713cf12d0114511c6105310a50f880ee20c790a39082e065204;
    decBuf[6705] = 256'h1d039401950050ff7efe0bfee8fdc8fdabfdc0fca4fbfdf975f810f7cbf5a4f4;
    decBuf[6706] = 256'h4bf363f2e4f1bef127f2c5f255f33af394f2a6f14af0a9ee90ed91ec06ec30ec;
    decBuf[6707] = 256'h3dedbdeeeef063f2b7f371f4c8f3c9f228f19fefa0eeb8ed8eed4eee13f0bbf2;
    decBuf[6708] = 256'he9f5e8f8a0fb1afeb5ff9500d9009b00d300a00072004800bb002401c201c502;
    decBuf[6709] = 256'hb90396049905d3064e087f0a8a0cee0e8910ff11cb120913d1129e126f12ee12;
    decBuf[6710] = 256'hfa133415af161418fc187b195419a61889177d1688156915861571168d17e718;
    decBuf[6711] = 256'h881a111c101d9b1d1d1d771b0d1929167013f710b70e410ded0bb90a100a7709;
    decBuf[6712] = 256'ha609780ad20b730d8c0e250ff60ecf0ddd0bf1087105360139fd9af94ff651f3;
    decBuf[6713] = 256'h26f217f169f1b4f108f3c1f369f49cf411f496f2cbf01bef02ee9decb5ebe3ea;
    decBuf[6714] = 256'hd6e957e8f2e6ade586e4c6e318e37ae2eae1ffe021e058dfd6debede2adf02e0;
    decBuf[6715] = 256'h3ee1b9e284e4b9e542e7dbe709e837e72ae665e439e22ee0dadea5dd6ddd06de;
    decBuf[6716] = 256'h4adfc5e090e2bce45de721e961ebd7ec2bee69eea1ee6eeee3edbcecafeb75ea;
    decBuf[6717] = 256'ha3e9c9e9bdea98ec84ef03f34ef671f82afb39fce7fb9cfb48fa13f98bf726f6;
    decBuf[6718] = 256'h3ef5bff4e6f44ef56bf6c4f766f95ffbb3fc63fe7cffafffddff070094ff2bff;
    decBuf[6719] = 256'h8dfe8bfd96fcf8fba2fb88fbcffb67fc17fdbdfd2afe8cfec1fef2fe1eff7cff;
    decBuf[6720] = 256'ha0ff69ffd3fe8ffd34fbf4f8e9f685f48ef3aef26af2a8f250f34ff494f50ff7;
    decBuf[6721] = 256'h0ef853f97df956f962f846f79ff517f4b2f210f187ef22ee81ecf8ea2de97de7;
    decBuf[6722] = 256'h64e631e676e745e9eceb1bef3ef130f33ff492f41cf340f11dee44eaa4e65ae3;
    decBuf[6723] = 256'h5be031dfd6decddf43e1a7e3e6e51de91becd4ee4df1e8f233f3eff2baf131f0;
    decBuf[6724] = 256'h66ee3bec2fea53e81fe776e6a9e64be8b4ea98ed18f172f370f69bf7f5f7fef6;
    decBuf[6725] = 256'h1ef642f416f20bf0b7eefeed36ee9beff6f1daf45af8a4fb7eff0b017402e202;
    decBuf[6726] = 256'hf00077fe93fbdaf861f621f441f385f3b9f4b3f627fa71fd4b01ea0444078d08;
    decBuf[6727] = 256'h2908cf0733062804c40184ff79fd9dfb68fac0f9bffa60fc3affb902f506f10a;
    decBuf[6728] = 256'h880d000e6d0e430d330c980ab8096408ab070207cf06fe067c0789087d09990a;
    decBuf[6729] = 256'h590bc20be20b380cba0c900d3f0f6b11761352150317ab171217cd15fe134e12;
    decBuf[6730] = 256'h35119c1027114e12a813a615fa162e18b7191c1b611c881d941e431fe11f7120;
    decBuf[6731] = 256'hbf200621f120b6203920861fe01e9f1e8b1e9d1e0f1fcf1fba2016225a238124;
    decBuf[6732] = 256'h4125aa254b25812462230922c420f11f321f541ff31fbc2044223d2491254127;
    decBuf[6733] = 256'h5a28f328682841270125c1228b1f8d1c0d19b31690142c14d213c814d4163819;
    decBuf[6734] = 256'h1c1c0d1e1d1f6f1f241fd01da51b6e18701529112d0d970a3d08f40691063606;
    decBuf[6735] = 256'h2d070d086109120b9a0c990d250e4f0e8f0d9b0c000b06091a069b0250ff77fb;
    decBuf[6736] = 256'hd7f77df535f498f45df69df83dfbb7fdf7ff6c013802f20249024a014cffe8fc;
    decBuf[6737] = 256'h04fa84f62bf407f2a4f1b3f2f3f429f828fbe0fdf0fee6ff9cffd0fe9bfd82fc;
    decBuf[6738] = 256'h83fbf8fa22fbe2fb1cfdebfe9c00b401b302e202b7024402dc01bc01d9019002;
    decBuf[6739] = 256'hf403bf056f07f808f709250a500a760adf0abc0bbf0c6d0d0b0e610eb00e270f;
    decBuf[6740] = 256'h3c0f500fd30eff0dfd0c090c6a0b870b0a0ce00c1c0e430f9c10841157127d12;
    decBuf[6741] = 256'h1412f8109e0ffd0d740c0f0b270a55092e095109b009060a550a9c0a860afd09;
    decBuf[6742] = 256'h3809190873067a0416027a006ffea3fdeafc41fc0efc83fbb1fa3efad5f9b5f9;
    decBuf[6743] = 256'h99f94af9a4f88bf7e5f5ecf310f25ff047ef48ee60ed8dec1aecb1eb92ebafeb;
    decBuf[6744] = 256'hfdeb74ece0ec1bede5ec32ecfeea82e9b7e783e6dae50de6dfe5b5e58ee59ae4;
    decBuf[6745] = 256'hfce3dfe32ee463e5dee6dde768e83ee817e8afe7cee7ebe739e822e8b6e753e7;
    decBuf[6746] = 256'h65e718e87ce947eb7cec95ed2eeeffed2dedbaec0bececeb7bec66ed02effbf0;
    decBuf[6747] = 256'hd7f287f4a0f539f620f7f3f766f8cff8aff8acf773f6f7f45ef48df45ff552f7;
    decBuf[6748] = 256'h2ef95afb65fdb9fe73ff1b00e8ff5dff8afecafd62fd42fdd2fd54fe6cfe2bfe;
    decBuf[6749] = 256'h7bfd75fc81fb22fbccfae6fa8dfb24fcfcfcc5fd7cfec3feaefe24fe3cfd1ffc;
    decBuf[6750] = 256'h13fbd9f906f946f852f7f3f663f6e1f56af5a7f4f1f31bf352f2cff188f147f1;
    decBuf[6751] = 256'h0cf1faf0a9f05ff087f0f4f079f13ef28cf215f2fcf009efa5ec66ea5ae87ee6;
    decBuf[6752] = 256'h41e679e678e719e912ebeeec23eecbee98eeb0ed35ec6aea36e9ade714e7e5e6;
    decBuf[6753] = 256'h0fe736e79ee7fde754e8a2e819e9dbe92febd0ec59ee58ef2aefabee9fedabec;
    decBuf[6754] = 256'h0decb6eb9ceb55ebbeea0dea96e9ace9d2eaa2ec49efc2f102f40df651f614f6;
    decBuf[6755] = 256'hfbf4caf2bff0e3eeaeed76ed75eeb9ef89f139f3c2f427f66cf73ef84bf9b3f9;
    decBuf[6756] = 256'h52fae1fa98fb0ffc7bfc67fc7ffb23fa82f889f635f500f4c8f3c7f468f6d2f8;
    decBuf[6757] = 256'h5afca5ffa3029504a4055205dc0388025401ab00de00c601ed0246042e05ad05;
    decBuf[6758] = 256'hd3056a05cc040304800398030404030583064e087a0a1b0d940f8b106b112711;
    decBuf[6759] = 256'hf20fda0edb0d500d250dff0c220d020d1f0dd60ddb0e151090115b139014a915;
    decBuf[6760] = 256'ha8168f17621888186618461829180f1827183c185018cd188019851a791b171c;
    decBuf[6761] = 256'hc11ba21a48190418da17e618f11a921d0c200221e321272264222c22f9211121;
    decBuf[6762] = 256'h3f20321fb31db41ccc1b4d1b271b4a1b691bf91bb01c561d9b1edf1fb2200b22;
    decBuf[6763] = 256'h9622c1224d221421f01e4f1cd6193a185a178e164717f01789181419ea182a18;
    decBuf[6764] = 256'h361719160d15d31300134012d8117911e9106610f00faf0f740f860f750f670f;
    decBuf[6765] = 256'h090f530ecb0c420b7709c707af0616068a050c05e60437045a039102da01c201;
    decBuf[6766] = 256'h0302db02de038c04eb04ce0417041203d801b100a5ffb0fed3fd43fd29fd70fd;
    decBuf[6767] = 256'hddfd17fe06feb4fd6bfd5dfde3fdeffe9500ad0112039e03c8035503ec024e02;
    decBuf[6768] = 256'hbe010701610020003400b100640139020303b9038f04580544062107b107cb07;
    decBuf[6769] = 256'hb30772075f0794070608c608b1098e0a570bda0b210c0c0c5b0b850a49092208;
    decBuf[6770] = 256'h62078507e407e708660acb0b100d8e0db50d4c0ded0c240c6d0b550b400b7b0b;
    decBuf[6771] = 256'h690bb60a8109b20786051004440307031f04ea051f073808d1084608c707bb06;
    decBuf[6772] = 256'h8105ae04a103ad02d001cd0093ff6cfe60fde0fb7bfa37f964f8f1f714f8b2f8;
    decBuf[6773] = 256'h42f9c4f9acf915f9eff7cbf5c0f3e4f1aff096effdee72ee9cee10ef78ef16f0;
    decBuf[6774] = 256'h6df01ef0a7ef8eee35edf0eb75ea76e98ee810e89de734e7d5e6b9e63be7b2e7;
    decBuf[6775] = 256'h75e860e9fee954ea6eeac8e9dae8bde7b1e677e5a4e4e4e37ce39be3f2e3a9e4;
    decBuf[6776] = 256'haee5e8e6b7e8e3ea59ec35eeeeee26ef8dee02eedbecceeb20ebc1eadeea60eb;
    decBuf[6777] = 256'h66ece5edb0ef61f179f212f3e4f265f2f2f1cff1eff1b8f2a3f381f411f5c7f5;
    decBuf[6778] = 256'h9df6a0f7daf801fac1fae3fa85fa2efa48fabffaadfbcafcd6fdcafe29ff0dff;
    decBuf[6779] = 256'h8afee4fdf6fc18fc16fb67fa08fa5ffa7efb24fd1dff81011d039204d6049904;
    decBuf[6780] = 256'h1003df00d3fef7fcc3fb1afb81fab0fadafab3fa1cfbbafb83fc6ffd4cfea2fe;
    decBuf[6781] = 256'hf1fea9fe3dfedbfd3afd4cfcf0fa4ff9c6f761f679f5a3f5b0f6eaf711f9d1f9;
    decBuf[6782] = 256'h39fa5cf920f8a5f6daf4a5f31cf21df1eff019f1d9f112f3e2f417f6bff6f2f6;
    decBuf[6783] = 256'hadf5def32ef235f0e1ee27ee5fee92ee1eef9cefc2ef9fef01efabee5dee74ee;
    decBuf[6784] = 256'h0cef0bf0fff05ef17bf12cf186f01af006f0f4ef05f0d8ef60efceee1deea6ed;
    decBuf[6785] = 256'h3aed27ed80ed74ee39f065f206f57ff7bff935fb79fb3bfb93fa2ef9e9f76ef6;
    decBuf[6786] = 256'h09f5c4f3f2f2cbf27af396f4f0f591f78af966fb92fd9dff79012903d2036b04;
    decBuf[6787] = 256'h3c04be034b039c02bf012f01e100f900bb010f03b00439060408b4093d0b080d;
    decBuf[6788] = 256'h3d0ee50e180fea0e170e580da90c0b0cee0b080cde0c1a0eea0f1612b6147b16;
    decBuf[6789] = 256'h721752180e1855173c16a31518159615091643176a18c319ab1a7e1bf11b5a1c;
    decBuf[6790] = 256'h791c961c191dbf1d821e381f0e209e20ec200421c32088205320e11ff01f3320;
    decBuf[6791] = 256'hb820a0217e228023e9234824b82301232c22622114215b21f321192340240025;
    decBuf[6792] = 256'h6825092507248722bc200c1ff31d5a1d2c1d021d281d051d251dcf1cb41cfc1c;
    decBuf[6793] = 256'h681df11d6e1e5e1ebc1da31cfd1a9318531648146c12bc10a30f700f9f0fc90f;
    decBuf[6794] = 256'hef0f1210f20f9c0f4e0fd70e140e290dcd0b2c0aa308a407bc06e6065a077c07;
    decBuf[6795] = 256'h5d07cd067905d803df010300cefeb6fd83fdb1fd2ffeeffe9eff7b00d1002001;
    decBuf[6796] = 256'hd80016002bff0efe68fc4ffb50fa68f93ef965f9cdf96bfafbfa7efbf4fbb7fc;
    decBuf[6797] = 256'h3afdb0fdf1fdb6fd39fd66fcd6fb54fb3cfb26fb61fb97fbe8fb4ffcc8fc5afd;
    decBuf[6798] = 256'hbcfd15fe46fe37fe45fe20fe41fe73feeafe7cff06008300b400a5006200ddff;
    decBuf[6799] = 256'h83ff52ff61ffa4ffe1ff2e008800dd0040018201a701860118017600b3ff30ff;
    decBuf[6800] = 256'he9fed3fe0eff44ff75ffa1ff94ff6fff0cff79fec8fd52fd11fd24fd36fd88fd;
    decBuf[6801] = 256'h79fd00fd6efc96fbcdfae2f944f97bf8f8f781f715f7daf6c8f698f66bf643f6;
    decBuf[6802] = 256'h1ff614f6f6f5a4f515f516f496f231f1ecef1aeff3ee16eff7eedaee23ee1eed;
    decBuf[6803] = 256'h2aec0deb4deae4e986e9f6e8dce8c4e8dae863e904ea9beafdeaebea59ea81e9;
    decBuf[6804] = 256'h45e81ee7c5e580e4aee33ae35de3fbe3fee438e60be731e70ee770e6a7e5bce4;
    decBuf[6805] = 256'h9fe392e2e4e185e1dbe1c7e222e4c4e56ce605e734e7b5e642e6d9e5bae564e5;
    decBuf[6806] = 256'h15e5cee4e4e4bbe5bee6b2e7cfe8f5e88de82ee89ee784e7fbe792e8b8e9dfea;
    decBuf[6807] = 256'hecebe0ec7eed61ed13ed6decaaeb5ceba3eb3aec3aed2eee8deea9ee8fee48ee;
    decBuf[6808] = 256'h32ee46ee7ceecdeeaaef06f1a7f211f5acf6b7f8fbf8bdf815f84af61ef4a9f2;
    decBuf[6809] = 256'h55f19bf063f062f1a7f2cef327f56cf693f79ff893f9b0fabdfb6bfc09fd26fd;
    decBuf[6810] = 256'hd7fc31fc18fbbff91df875f7dcf60af731f88bf9cffaf6fb69fc8cfc2dfc10fc;
    decBuf[6811] = 256'hf6fb6dfc04fddcfda6fe28ff10ffa4fea5fd6bfcf0faf1f9adf8daf767f78af7;
    decBuf[6812] = 256'h67f8ddf9a8fb58fd51ff1d00d6000f0176008eff13fe48fc1cfa11f8bdf603f6;
    decBuf[6813] = 256'h5bf58ef576f648f7a2f843faccfb31fd76fe48ff22ff2efe93fc9afa36f8f6f5;
    decBuf[6814] = 256'h80f4b4f3f2f30af5d5f686f80ffaa8fa33fb5dfb36fb59fb79fb5cfbdafa33fa;
    decBuf[6815] = 256'h9cf961f997f949fa1ffbaffbc9fb82fbbffa08faf1f931fa31fb6afce6fd4bff;
    decBuf[6816] = 256'h8f000a0209039403bf03ff020b02ee0095ffadfe2efe55fe8fff5e018a032a06;
    decBuf[6817] = 256'ha4083f0ab50b090dc20dfa0d930ec20eec0ec50e170eb80d9b0dea0def0ee30f;
    decBuf[6818] = 256'hc11050119f11e611d4123014d115ca172e1ac91b3f1d931e4c1f6520fe202c21;
    decBuf[6819] = 256'hae20a11f221e231d981c6e1c2d1dad1ede207f23f825382818295c291f290628;
    decBuf[6820] = 256'h6d27e226b826de264727a6273528b8282f2970293529db288a2840289e285429;
    decBuf[6821] = 256'h0b2ae02a372b1d2bd52a3e2a3f29902874271a2633250c244c23e322c4226d22;
    decBuf[6822] = 256'h53223b22fb21e7218e211c217a208c1f301eeb1c701b0b1a2319a51832185518;
    decBuf[6823] = 256'hb31897187d18d61792164d157e13ce114510460f5e0ee00db90d960db60dd30d;
    decBuf[6824] = 256'h840dde0cf00b550acc089b0690043c0307025f0192017a024c03a6048e056006;
    decBuf[6825] = 256'h870664060506750556044903c90164007dffaafed0fef3fe52ff6fff20ffaafe;
    decBuf[6826] = 256'h69fe07fe19fe49feb1fe0eff63ffdcff6e001f01c50131029302a50295024b02;
    decBuf[6827] = 256'hd301610117010a015f010402da026903b803a0033403ab022d021d026702fa02;
    decBuf[6828] = 256'hd2039b045205f80564067806d7059304f102690104001cff46ff9f0041023a04;
    decBuf[6829] = 256'h1606c6076e08a1087308a00794061405af030e028500bafe85fdddfcaafc35fd;
    decBuf[6830] = 256'hb3fdc0feb4ff91002101070190004cff4efdeafaaaf89ff64bf588f5c1f5c0f6;
    decBuf[6831] = 256'h04f883f8f6f8d3f874f8e4f7f9f6dcf5d0f496f3c3f2b7f17df056ef49ee9bed;
    decBuf[6832] = 256'hfdec53edd6ed7cee13ef27efceee1beee6ec6beb06ea65e84ce74de67be6fae6;
    decBuf[6833] = 256'h53e83be9b9e993e99fe843e75be631e657e6c0e65ee7eee770e888e89ee88ae8;
    decBuf[6834] = 256'h55e8e3e723e738e65be5cbe47ce4f3e48be5ede546e677e64be608e614e635e6;
    decBuf[6835] = 256'h8fe62ce799e7fbe754e844e835e842e836e86de8c7e81ce995e907ea51eaaeea;
    decBuf[6836] = 256'hebea0ceb2aeb45eb1cebbbea27ea77e9d1e890e8a3e844e989eacdeb9ded4def;
    decBuf[6837] = 256'h65f0fef08af10bf1b2ef6dee9eec69eb31eb64eba9ec78eeadefc5f0c4f1acf2;
    decBuf[6838] = 256'h2bf3eaf353f4b2f408f5baf473f4dbf303f374f225f2def1f4f12ef240f2b2f2;
    decBuf[6839] = 256'h37f3d8f3c6f421f666f78df89af948fae6fa76fbc4fbacfb40fb1afa9ff83af7;
    decBuf[6840] = 256'h52f6d4f547f63bf7d6f8cffa23fcd3fd5cff5b008a00b7ffaafe2bfd60fbaff9;
    decBuf[6841] = 256'h27f828f79cf61bf727f8edf919fc24fe00003501dd01100285010601faff7afe;
    decBuf[6842] = 256'h15fd74fbebf952f9c7f89df810f933f952f96ff9bdf934faf7fa16fc23fdd1fd;
    decBuf[6843] = 256'hf1fd9bfde4fcdefba5fa7ef971f87df7dff689f6a3f649f737f814f950fa23fb;
    decBuf[6844] = 256'h96fbfffbdffbc2fb40fbc9fa32fa33f93ef8e3f69ef577f46af3bcf2dcf2a5f3;
    decBuf[6845] = 256'hf9f4f7f65bf93ffc30fef5ff9001db019701de0055ff8afddafbe0f914f9d7f8;
    decBuf[6846] = 256'h7ff9e4fae2fcbefeea0060022c03e5038d042605b1053006a306c606a6068906;
    decBuf[6847] = 256'h6f0628066906cb069007e308850aee0c2e0fcf1193132e150f16531690163917;
    decBuf[6848] = 256'h6c179a17c417eb178217231793167916c0160117d9171519911ac21c621f2721;
    decBuf[6849] = 256'h672347241325d5242d24c82283215c209c1f341f931f5c20e4216d23d2241626;
    decBuf[6850] = 256'h952608272b2789276d271e274926d3246e2370211c206b1e531d541c6c1bee1a;
    decBuf[6851] = 256'hc71a301b4c1cf31d7b1fe0206c219621d620561f251d841a56177c13e6108c0e;
    decBuf[6852] = 256'h440de00cf00d8b0f0111dd128d1435150215be139a11f90e800c9b09e3066904;
    decBuf[6853] = 256'hce02c3006fff3afe72fe0bffad00a6028204b7055f062c06a1057a0421037f01;
    decBuf[6854] = 256'hf6ff2bfe7bfcf2faf3f968f9e6f9a6fa9afbb7fc77fd25fe84fea1fe87fee1fd;
    decBuf[6855] = 256'hc7fc6efb29fa03f943f820f8bef8faf975fbdafc7cfe94ff9300c2009800d8ff;
    decBuf[6856] = 256'h29ffcafee7fed2ffef00fc016402c3026d021e02a801670153016501d7017902;
    decBuf[6857] = 256'h92039f049305f2050f06c0051a05ae042404a70356030c033403a2037f049b05;
    decBuf[6858] = 256'ha8069c073a0857083d08f607b5072b074306e704a303d0021002330292022203;
    decBuf[6859] = 256'h3c0324038d02b501b200beffe0fe51fe02fe1afe86fe10ff69ff9aff50ff87fe;
    decBuf[6860] = 256'h4bfdd0fb05fa55f8ccf6cdf542f56cf52cf6abf7aaf892f9bcf949f955f8f9f6;
    decBuf[6861] = 256'h58f55ff30bf25af042ef43eeb8ed39ed13edf0ecd0ec27eddeede3ee1df0eff0;
    decBuf[6862] = 256'hfcf165f245f2eff104f1a8ef06ee0dec31eafce8e4e717e8a2e81dea82eb23ed;
    decBuf[6863] = 256'h3cee3bef69ef3fef7fee8bed6fec62ebb4ea94ea77ea91ea08eb74ebfeeb9fec;
    decBuf[6864] = 256'h0bed46ed7bed4aed3ced7fedecedabee97eff5ef12f0c4efbfeecaed2ced9dec;
    decBuf[6865] = 256'h4eec36ecf6ebe2ebaceb9cebe6eb79ec51ed54ee48ef25f07bf0caf082f016f0;
    decBuf[6866] = 256'h8defecee55eef3ed99ed89edd3ed4bee1eef21f0cff02ef112f1f2efe6eeaced;
    decBuf[6867] = 256'hd9ec66ec14ed31ee8aef2cf1b5f2b4f33ff469f4f6f302f366f1deef79ee34ed;
    decBuf[6868] = 256'h5eed1eee9eefcff1daf33ef6d9f7b9f8fdf8c0f817f818f7d4f501f541f493f3;
    decBuf[6869] = 256'h34f3def2f8f26ef306f4def4e0f51af741f8e7f970fbd5fcbdfde7fd74fd80fc;
    decBuf[6870] = 256'h24fbdff90df99af877f815f918fa0cfbe9fbecfce0fd7efed4fe23ff3bff50ff;
    decBuf[6871] = 256'h3dff07ffb6fe31feb4fd22fdbffc8afc9afcc6fc09fd5efdd7fd49fe93fed5fe;
    decBuf[6872] = 256'h12ff5fffb9ff57001901d0011702020251014c00ccfecdfde5fc67fcdafc43fd;
    decBuf[6873] = 256'h20feb0fefefe16ffd5fe9afe65fe54febcfe4fffffffa6003d0178016601f400;
    decBuf[6874] = 256'h1700fafeeefd3ffde1fcfdfce8fd44ffe6006f026e03550428059b0504066306;
    decBuf[6875] = 256'h0c068a0585040503a001b800e5ffa500df010304a406d209f60bae0ebe0fb410;
    decBuf[6876] = 256'h9511511197107f0f1a0e1c0cc80a93095b09c00abe0caa0f2913741672192b1c;
    decBuf[6877] = 256'hef1de61e311fed1e3d1db41be919b4180c18d917c118901abc1cc71ea3205322;
    decBuf[6878] = 256'hdc23db24c3254126b4261d27fd266e26b725e1248b243c24252491241a257425;
    decBuf[6879] = 256'h2626fc26c5271929012ad32afa2a912ab429eb28ff2722279226db2506253c24;
    decBuf[6880] = 256'h5123742257227122b9225023d92333244324f9233123f421cd20271f9e1d391c;
    decBuf[6881] = 256'h981a7f19e618ff17d41761173e17e01650166515c714fd137b139213d3130e14;
    decBuf[6882] = 256'h20146d13391269103d0e9d0b230988077d05b104f703a0049f054007c908940a;
    decBuf[6883] = 256'hd20a9a0a350993072a058f0383012f00fbfee2fd15fe43fe6affc4000802db02;
    decBuf[6884] = 256'h9b03be039e0381036703f0022e024301e7ff45febdfcbefb32fb5dfbd0fb0afd;
    decBuf[6885] = 256'h30fed7ff5f015e02ea0268038e032603c70237024c016f006cff78fe19fe36fe;
    decBuf[6886] = 256'hb8fe5eff2100d8004f01e60197023d03a903e403ae03fc0226025d01da003400;
    decBuf[6887] = 256'h9cffecfe16fe13fd65fcc7fbaafbf8fbcefcd1fdc5fee2ff55007800d9ff10ff;
    decBuf[6888] = 256'hf1fd97fc53fb2cfa1ff92bf88df770f7bff706f872f8adf877f826f8bff746f7;
    decBuf[6889] = 256'h94f6edf5d4f4c8f38ef2bbf1fbf0d8f0b9f09cf0b6f09ef0b4f079f044f0f2ef;
    decBuf[6890] = 256'h8bef2defc0ee94ee6cee48ee27eee1edb3ed9aed75ed52ed0eed85ecfbeb7eeb;
    decBuf[6891] = 256'h2deb1eeb46eb52eb1bebc1ea3ceae3e9d2e9e1e9efe9fbe998e93ae9e5e8c4e8;
    decBuf[6892] = 256'hf6e87fe908ea86eaf7ea24eb66ebbbebdceb0eec3cec23ecfeebc0eb44eba3ea;
    decBuf[6893] = 256'he1e92ae983e843e808e81ae88be8d5e84de900eaa6ea69eb20ec67ec52ec3eec;
    decBuf[6894] = 256'hc1eb90eb64eb3ceb17ebe0ea5eeae1e96fe926e933e9a0e925eaeaeaa0eb47ec;
    decBuf[6895] = 256'hb3ec3ced96eda6ed97ed39ed84eccdebc7ea19eaf9e9dde994ea69eb33ecb5ec;
    decBuf[6896] = 256'hfcecbcec81ec6fec3eec6aece3ec54ed14eeffeeddefa6f05df1a4f163f1daf0;
    decBuf[6897] = 256'hf1ef53efc4ee75ee5dee48ee0deed7edc7edb8ed4bee4bef84f054f204f41df5;
    decBuf[6898] = 256'h82f60df737f7c4f6d0f574f42ff3b4f1b5f02af0acefd2efc6f022f2c3f32df6;
    decBuf[6899] = 256'h6cf878fa44fbfdfbc5fb2cfb44fac9f8fef6d2f45cf308f2cbf103f268f309f5;
    decBuf[6900] = 256'h02f756f806fa1ffb84fc6cfd3ffe65fe42fea4fd68fc41fbe7f9a3f8d0f710f7;
    decBuf[6901] = 256'hedf60df79df754f829f92cfa20fbfefb8dfc10fd28fdbcfc5afcb9fb21fb98fa;
    decBuf[6902] = 256'h62fa73fa9ffa17fb89fb2bfceefc70fde7fd28fe3cfe2afef9fdcdfd6ffd4bfd;
    decBuf[6903] = 256'h40fd5efd79fd71fd2dfda5fccdfb76fb91fb37fc7bfd1dffa500a40130020203;
    decBuf[6904] = 256'h7503de03fe03e1035e03b8022102e6013f02d102820328041605f305f6063008;
    decBuf[6905] = 256'h5709640a120bb00b060c550c9c0c860c730c190cc80bb90be10b670c080d740d;
    decBuf[6906] = 256'h4c0e4e0f43101d12f913a915a217f618b019581a251af719cc190d19a4188418;
    decBuf[6907] = 256'ha1182419291a631b8a1c961d8a1e291f7f1f0120ea1f2b203e2009201920ed1f;
    decBuf[6908] = 256'haa1f551f1e1fec1e501ffe1fd42010228b238a242c26b427b3283f296929a928;
    decBuf[6909] = 256'h29275e2532232721d31f1a1fe21e151f431f1620d620ca21a7227023bf230624;
    decBuf[6910] = 256'hc5233c2377222421821f891dad1b781a6019c7189818c2188219bc1a371c9c1d;
    decBuf[6911] = 256'h841e031f431ec31cf81a51188c164d14d71283114e10350f9c0e6e0eec0eac0f;
    decBuf[6912] = 256'h151074101e109b0fc50ec20dce0c720b8b0a6409f108ce08ae08cb08e5089e08;
    decBuf[6913] = 256'h32085a079006da0504057404f103da031b04a404fd040e056b045203f9015700;
    decBuf[6914] = 256'hcffe6afd82fc03fc90fbb3fb12fcdbfc92fd38fea4feb8fea6fe96fe6afe5cfe;
    decBuf[6915] = 256'h07fe78fda1fc9efbeffa51fafbf915fa5cfaf4fa7dfb1efcb5fcc9fc93fc01fc;
    decBuf[6916] = 256'h29fb60fa75f9d7f847f890f719f782f647f612f601f62ef68bf6f8f67df71ef8;
    decBuf[6917] = 256'hb5f866f90cfa4dfa39fabcf90af963f8a1f71ef778f60cf682f505f573f4eaf3;
    decBuf[6918] = 256'h6cf33cf32df355f3c2f364f4fcf485f5dff5cef567f5b9f4e3f3e1f2edf14ef1;
    decBuf[6919] = 256'hf8f012f15af1c6f176f2edf259f394f33bf388f2b2f1aff001f0a2ef85efd4ef;
    decBuf[6920] = 256'h7af011f111f205f3a3f3f9f3dff309f306f2cdf051ef52ee6bed98ecd8ebfbeb;
    decBuf[6921] = 256'h5aec23ed77eebbef36f1cff15bf285f2abf2cef2aef258f2d5f15ff11ef1e3f0;
    decBuf[6922] = 256'hf5f026f134f10cf1d0f083f03df046f05ef0b1f02af19cf13ef201f3b7f35ef4;
    decBuf[6923] = 256'hf5f430f51ef50ef5c4f481f42cf4dff3adf3c9f334f411f52ef687f76ff8edf8;
    decBuf[6924] = 256'h61f93ef9dff889f806f88ff74ef713f749f7dbf7daf814fa3bfbfbfba9fc08fd;
    decBuf[6925] = 256'hecfc9dfc26fc8ffb06fb89fa37fa0bfa4efa04fb23fc7dfd1eff370036010701;
    decBuf[6926] = 256'h89007cff42fe1bfd0ffc60fb02fb1efba1fb77fcb3fd2eff9300d80156023002;
    decBuf[6927] = 256'hc701aa009eff64fe3dfd7dfc15fcb6fb0cfc5afcd1fc3dfdc7fd20feb2fe14ff;
    decBuf[6928] = 256'h4aff5afff3fe45fe6ffda6fc58fc10fc26fc61fc97fce8fc32fd8ffde4fdd9fd;
    decBuf[6929] = 256'h7ffdc9fcaafb9dfaeff90efa9efa89fba6fcb3fd1bfe3bfe1efe04fe8dfdf6fc;
    decBuf[6930] = 256'h6cfc84fba7faddf95bf914f9fef860f9ddf990fa95fb44fc21fdb1fdfffd46fe;
    decBuf[6931] = 256'h5cfe21fec8fd15fd10fc1cfb3efaaef9fdf9d3fad5fb0ffde2fda2fe0aff69ff;
    decBuf[6932] = 256'hbfffdaffc2ff2aff53fe50fd5cfc7efbeffad4fabdfa29fb01fc03fd3dfe64ff;
    decBuf[6933] = 256'hbe00a5017802eb02c8026902a001b500d8ff48ff2effa5ff670052013002f902;
    decBuf[6934] = 256'h7c03f203330447043504c3035c03e402b302df022203a70324047604dd045505;
    decBuf[6935] = 256'hc705a40682078408be09910a9e0b4c0cea0c400d5a0d430d020da00c230c700b;
    decBuf[6936] = 256'hf90ae30af70abc0bdb0c340ed60fee1053123b1362142215d0152f16d9152215;
    decBuf[6937] = 256'h4c144a13e11201139013b014bc15f616c917d6188419611a641b121cb11c071d;
    decBuf[6938] = 256'h211d391d231de81cd61cc61cb71c8f1c531cda1b681b3c1b491bff1bea1cc71d;
    decBuf[6939] = 256'hca1e331f521ffc1e451e9f1ddc1c251c7f1be81a5e1a291a5a1afc1a931b6b1c;
    decBuf[6940] = 256'hfb1c151d2d1dc11c5e1ce11b2f1b591a5619d6170b165b14d2126d11e2106410;
    decBuf[6941] = 256'h3d10a610c6101c1136114e110d11d21031106f0f830e670d0d0cc90aa2099508;
    decBuf[6942] = 256'ha1070307ad065e0647065c0670063a06e90547055904fd02b8013d003efffafd;
    decBuf[6943] = 256'h7bfdbbfc53fcb5fb25fba2fa5bfa1afa07fad1f980f918f985f8fcf77ff70df7;
    decBuf[6944] = 256'ha6f648f6dbf556f5d9f467f43bf413f41ff4fef3e0f38ef341f3e7f292f25bf2;
    decBuf[6945] = 256'h15f29ff10cf134f06bef80ee21eecbede5ed2cee6dee81ee93ee82ee56eef9ed;
    decBuf[6946] = 256'hd4edf5ed27ee9eee10ef94efeeef3ff06bf05ef052f0d9ef26ef50ee4ded9fec;
    decBuf[6947] = 256'h01ecabebc5ebddeb49ecabec6fed5beef9eec2efdcefc4ef58efcfee0aee88ed;
    decBuf[6948] = 256'h11edfbece8ecf9ec6bedf0ed6deeffee89efbeefefeffeeff0effdef08f0feef;
    decBuf[6949] = 256'hf4ef0df015f029f03cf0feef93ef0eef4aeec7ed50ed3bed75edf3eda5ee7bef;
    decBuf[6950] = 256'h44f02ff1cef124f20af2c2f182f11ff10ef11ef12df155f161f156f160f18df1;
    decBuf[6951] = 256'ha6f1aef1b5f170f130f107f1f0f020f17ef147f210f32ff4eff49ef57bf6d1f6;
    decBuf[6952] = 256'hebf6d4f63cf664f528f4adf248f103f085eff8ef32f156f361f5c5f705fa10fc;
    decBuf[6953] = 256'h64fd1dfec5fe2cfee8fcc4fab9f8cdf5dbf3ccf27af25af3aef4daf6e5f849fb;
    decBuf[6954] = 256'h89fdfefecaff0800400041fffdfd82fcb7fa82f9d9f8a6f8d5f8a7f9b4faa8fb;
    decBuf[6955] = 256'h86fc88fd7cfe99ffa6000e012e01d80021001cffe2fdbbfc61fbd6fa58fa32fa;
    decBuf[6956] = 256'he0fabdfbc0fcfafd21ff2d00dc003b011e019b00f5ff07ff2afe27fd33fc95fb;
    decBuf[6957] = 256'h92fae4f946f929f9abf9b1faebfb66fdcbfeb3ff8500f800d500b600b3ff79fe;
    decBuf[6958] = 256'haafcfafa71f90cf881f756f7caf7bef89bf99efad8fbaafc6afd19fe38fe1bfe;
    decBuf[6959] = 256'h01fe5bfd6dfc51fb44fa50f9b2f85bf876f8bdf8fef839f96ef9e0f965fa29fb;
    decBuf[6960] = 256'he0fb86fc1efd59fd6bfd3afdf0fc5dfcacfba7fab3f915f985f86bf8b2f84af9;
    decBuf[6961] = 256'h21faebfad6fbb3fc43fdc6fd0dfe22fe0ffefdfdccfda0fd5dfdf0fc6bfc12fc;
    decBuf[6962] = 256'hc1fbb2fbbffb14fc61fcf7fc8efd8efe82ff9e00ab01590279022302a0019b00;
    decBuf[6963] = 256'ha7ffc9fe00fe7dfd66fd7bfd2cfe31ffb1001602b703d0046905f405ca05a305;
    decBuf[6964] = 256'h3b05dc0413045c03b602f301a5015d01c90153025f03b804fd057807dd08c509;
    decBuf[6965] = 256'h430a1d0afa095c093f09f108d90898080f0892072007d606e4065107d5077608;
    decBuf[6966] = 256'h6409420a7e0bf90c5e0ea30f21104710df0f410fb10efa0d240d5b0cd80b620b;
    decBuf[6967] = 256'h4c0bae0b730c5e0d7a0e870fc110941107126f1250123312b0113a11cd106b10;
    decBuf[6968] = 256'h361025101710ef0ffb0f3210b4109c117912091358136f132e13cc124f12bd11;
    decBuf[6969] = 256'h34116f10ec0f460f050ff20e270f780fe00f8e103411cb11551266123612ce11;
    decBuf[6970] = 256'h3b11b21011107a0fa20ed90ded0c4f0cf90bdf0bf70b380c720ca80c1a0d640d;
    decBuf[6971] = 256'hc10dfe0df30d990d2c0d890cc70b440b6e0aa50986087907cb062d06d605f105;
    decBuf[6972] = 256'h3806cf065907d6076808f1084b097b094f09f20854089107da06d5059b047403;
    decBuf[6973] = 256'h1b0233016100edffcbff2900b9003c011202db02c603a30433054d0506054304;
    decBuf[6974] = 256'h58033c02e2009eff77fe1dfd92fc14fcedfb56fcf4fcbdfd74fe4aff13009600;
    decBuf[6975] = 256'hdd00c80065007dff21feddfcb6fbf6fa47fa67fa84fad2fa49fbb5fbf0fb26fc;
    decBuf[6976] = 256'hf5fbe6fbbefb9afb63fb31fbf1fac7faa2fa72fa53fa36fafef9d9f9a8f97df9;
    decBuf[6977] = 256'h6cf97bf99cf9dbf91bfa55fa7afa81fa62fa0efaa1f9fef867f8def784f753f7;
    decBuf[6978] = 256'h45f788f7f5f797f85af910fa87fac8fadcfa82faf0f93ff9c9f888f84df85ff8;
    decBuf[6979] = 256'h90f8d9f81cf971f9d4f932fa6efa8ffa85fa45faebf965f9e8f8b7f88bf8cef8;
    decBuf[6980] = 256'h3bf9c0f961faf8fa5afb90fbc1fbcffbf8fb1cfc27fc31fc16fcfdfbc8fb98fb;
    decBuf[6981] = 256'h79fb73fba1fbf3fb56fcb3fc08fd3ffd85fdb3fdedfd30fe70fe78fe71fe33fe;
    decBuf[6982] = 256'hc8fd60fd03fddefcd3fcf1fc1ffd59fdabfd24fef7fefaffee000b02cb02ee02;
    decBuf[6983] = 256'h8f02ff01e000d3ff25ff47feb8fd69fdb0fd1dfef4fef7ff31010402c4027203;
    decBuf[6984] = 256'h92033b03ed0247028401cd00f7ff2effacfe35fef4fd2ffef3fe13006c01b102;
    decBuf[6985] = 256'h83034304ac048c043604b3030d034b022b011f002aff4dfef7fd45feebfeaeff;
    decBuf[6986] = 256'h9900770179022803c603e303c803520364028601bd00d2ff34ff6bfee8fda1fd;
    decBuf[6987] = 256'h8bfd15feb5fe78ff63000101910114025b0271025d0204029201f0002d0076ff;
    decBuf[6988] = 256'ha0fed7fdecfc4efcf8fbddfb54fc17fdcefd74fee0fe42ff78ff68ff3bffdefe;
    decBuf[6989] = 256'h40fe52fd75fcacfb29fbe2faccfae0fa39fbabfb30fc89fcfbfc27fd4ffd73fd;
    decBuf[6990] = 256'h94fd9efd71fdf5fc30fc45fb29fa1cf96ef80ff8f2f775f81bf934fa41fb7bfc;
    decBuf[6991] = 256'h4dfdc0fde3fd84fd82fc8dfb71fa64f9b6f857f83af854f8fbf8bdf9ddfae9fb;
    decBuf[6992] = 256'hddfcfafdbafe22ff42ff5fff10ff6afea8fdbcfcdffb16fb93fa4cfa62faebfa;
    decBuf[6993] = 256'hb0fb9bfcb7fdc4feb8ff5600e60034014c0162012701cd001b0074ffb2fe2ffe;
    decBuf[6994] = 256'h47fe88fe38ff0e00d700c3011e0363048a059706b9065b0658051e04a302a401;
    decBuf[6995] = 256'h19019a007400dd003b01cb01b602940396048b0529064506600648063206f705;
    decBuf[6996] = 256'h9e054d05e5046d041c04d203c50301046404f7048105fe054f0640061806dc05;
    decBuf[6997] = 256'hbb05b105ba05e305fa05e505ad053c058904b403ea0234028d0121010e018b01;
    decBuf[6998] = 256'h7e02b80333059806dd075b083508cc07ef06b305e00420047203130383020102;
    decBuf[6999] = 256'hb9017901b3010d029f02280382039203a103c903ed033a04800489042f049103;
    decBuf[7000] = 256'hce021802a10160014c015e016e01b80116029b02f50266039303bb03af037803;
    decBuf[7001] = 256'h4603f302bc02b202bc02e5022803310308039802e5013f01a7006c0013000300;
    decBuf[7002] = 256'hd7ffaeffa2ffd9ff4700ea0081010a021c020c02c2017f015b013a0130013901;
    decBuf[7003] = 256'h31010b01cd0083002900d4ff71ff2eff0afffffe1dff5dffb8ff0d005a007800;
    decBuf[7004] = 256'h5c00e0ff1cff31fe14fd54fca6fb86fbdcfb2bfc01fdcafdb5fe53ff1c006b00;
    decBuf[7005] = 256'h82006d00e3ff43ffabfe22fec8fdb8fdc7fdd4fde0fdd5fdb7fd78fd1dfdc8fc;
    decBuf[7006] = 256'h91fc5ffc56fc6ffcc1fc24fd9cfdeefdfcfdeffdb2fd65fd1ffd04fdebfc02fd;
    decBuf[7007] = 256'h09fd1bfd43fd7bfdcefd47feb8fe20ff48ff54ff1dffc3fe56feeffd76fde4fc;
    decBuf[7008] = 256'h82fc28fc18fc44fca2fcf7fc5afd9dfdc1fdb6fd84fd57fd0cfddafcbffce8fc;
    decBuf[7009] = 256'h59fdebfd4dfea6feb7fe4ffea2fdfbfc39fc82fb3bfb25fb60fb01fcc3fce3fd;
    decBuf[7010] = 256'heffe9effbdffa1ffeafe14fe11fd63fc85fbf6fa73fa2cfaebf9d7f9e9f95bfa;
    decBuf[7011] = 256'he0fa81fbedfb28fc39fc29fcdffb9dfb60fb3ffb49fb9bfb2afcdbfc81fdedfd;
    decBuf[7012] = 256'h01fe84fdb0fcaefb74faa1f9e1f8bef89ff8f5f878f9eef95afae4fa3dfbaffb;
    decBuf[7013] = 256'hdbfbb3fb46fba4fa0cfa83f92af919f963f9dbf94dfab4fa2dfb9ffbe8fb2bfc;
    decBuf[7014] = 256'h37fc2cfcfafba8fb45fb02fbadfa76fa80fac0fa1bfb70fb91fb73fb21fbbefa;
    decBuf[7015] = 256'h96fabafa33fba5fb0cfcfffbc2fb5ffb1cfb10fb5dfbb7fb0cfc59fc9ffcdffc;
    decBuf[7016] = 256'h29fd83fda7fdb2fd80fd1cfdd9fc9dfcbefc18fd85fdecfd4afe86fed3fe2dff;
    decBuf[7017] = 256'h82ff8dff6fffe6fe0efe0cfd17fc79fb23fb3dfbb4fba2fcbefdcbfebfff5d00;
    decBuf[7018] = 256'h7a002c0085ff19ffdefef0fe83ff3300d9007101d301e5019401f100adff0cfe;
    decBuf[7019] = 256'hf3fc8efb60fb8afb4afc83fdfffefeff42016902290392037203a9025501b4ff;
    decBuf[7020] = 256'h2bfec6fcdefbb4fb8dfbf6fb94fc5dfd14feeafeedff9b00b801780226038503;
    decBuf[7021] = 256'ha20353037e02b401c900ecff23ff6cfe66fd72fc95fb05fb1ffbc6fbdffc85fe;
    decBuf[7022] = 256'h0e000d01f5017302e6020903aa0254029d019800a4ff05ff76fe27fe10fe25fe;
    decBuf[7023] = 256'h60fe96fe07ff6fff0200b200880151023d039b03b8036a039402cb0114019d00;
    decBuf[7024] = 256'h3100f6ff9dff2bfffffef1fe77ff3b00270104029402ae02670251023d027302;
    decBuf[7025] = 256'hc4020e0351035d033c03320317030e03f802e302b7027a0240020b02e901e301;
    decBuf[7026] = 256'h15026f02f40295032c048e04a0044f04ca0306031b027c01ed009e0087009c00;
    decBuf[7027] = 256'hfe00c301ae028b035504d7041f050905a70406049a0338030203d102e0020803;
    decBuf[7028] = 256'h14034b039103d103fa03e4038b03ed022a027301cd003600fbff0d003e008700;
    decBuf[7029] = 256'h1a01f201f502e903c7041d056b05f4045d04850382028e01f000600046008e00;
    decBuf[7030] = 256'hfa0083014802ff02d4039e045405cb05e1057f05de04c5036b0227010000f3fe;
    decBuf[7031] = 256'h45fea7fd50fd9ffd45fe89ff8801ec032b0637088b09c809000a010960076705;
    decBuf[7032] = 256'h0303c30022fe5efc0cfc56fcaafd5bffc40104047a05ce0602083a08d308a508;
    decBuf[7033] = 256'hd20779063405b90354026c01ee007b009e00bd0014016201d9014502f6029c03;
    decBuf[7034] = 256'h5e044a05660626078f07ae0792074307cc066006d70536051d0410031c027e01;
    decBuf[7035] = 256'h9b011d02f302f603ea04490566054c056305a405b8058205cf049b0374026701;
    decBuf[7036] = 256'hff001e01e701d302ef03af045d05bc058606d4061b073107a706070644055904;
    decBuf[7037] = 256'h7b037902ca01ed005d0043002b0097002101c20184023b031104a104ef04a804;
    decBuf[7038] = 256'he503fa02dd011e01b5009500b200cc00e400ce0009016301f5017e02b402c402;
    decBuf[7039] = 256'h980255020002c9016f011a018b00020085ff33ff25ff68ffa4ffdbfff9ff0200;
    decBuf[7040] = 256'heaffe2ffdbffe1ffe7ffd8ffa5ff59ff13ffd3fecbfee2fe3bffa8ff0f005200;
    decBuf[7041] = 256'h5e002700cdff60fff9fed1fef5fe42ff9cff22007b00ac009d005a00d5ff34ff;
    decBuf[7042] = 256'h71feeffd78fd62fd9dfd3efed5fe5fff94ff64ffdffe3efed2fd97fdf0fda3fe;
    decBuf[7043] = 256'ha8ff9c007a01d0011e0236024c025f024e02fc0178018f0073ffb3fe04fee5fd;
    decBuf[7044] = 256'h3bfef2fe69ff00006200df005101b80116023a021902bf015201eb00c300cf00;
    decBuf[7045] = 256'h0601380165018f01a501c80119027c02f4028603e9034204730481043f04ea03;
    decBuf[7046] = 256'h5b03d102540223026d02cb023803820374033803d50292029e020103af038504;
    decBuf[7047] = 256'h4e050506ab06170703073f061f05c60381025b0134019d017a02430363042305;
    decBuf[7048] = 256'h1706f406bd074008870846089607c006bd050f053204a203eb02a40263024f02;
    decBuf[7049] = 256'ha902fa024403a103de034104b9042b05cd0539064d06f4058205c2040b046503;
    decBuf[7050] = 256'hce026b0236020502d901e601230286021903ca037004dc04f00472047f03ff01;
    decBuf[7051] = 256'h340084fe6bfd6cfc3efcbcfcc9fd8effba0130038404c10489048a03e901f0ff;
    decBuf[7052] = 256'h8cfd4cfbabf8e7f695f6dff6bbf8e7fa88fd0100f800d8011c02df0136013700;
    decBuf[7053] = 256'hf3fe77fdacfb78fa5ff960f8d5f757f797f6a3f583f5d9f5c4f620f8c2f9dafa;
    decBuf[7054] = 256'h3ffc27fdfafd20fefdfd20fdaafbdff9aaf892f75ff78df763f7f0f641f6a3f5;
    decBuf[7055] = 256'h4df533f5aaf56cf623f7f9f735f9b0fa7bfca7fe87ff43ff93fd2afb45f88df5;
    decBuf[7056] = 256'hc8f376f3c1f305f4bef4f6f429f558f582f5f5f5a3f6fff7fdf9d9fb05fe7bff;
    decBuf[7057] = 256'hbfff06ff7dfd18fcd3faacf9ecf83ef861f75ef6aff5d2f4b5f438f5def5ccf6;
    decBuf[7058] = 256'he9f7f5f82ffa56fb16fcc4fc23fd06fd84fc3dfcfcfbc1fbd3fbc2fb79fbb0fa;
    decBuf[7059] = 256'h74f94df840f792f672f63cf727f883f9c7fa42fca7fd8ffeb9fe93fee5fdc8fc;
    decBuf[7060] = 256'hbbfb53fb33fb89fbd8fb1ffcb3fbdbfad8f92af949f913fa66fb08fd91fe2aff;
    decBuf[7061] = 256'h58ffdafe1afee0fc65fb66fadbf9b0f9d7f985fa63fb65fc14fd73fdc9fd17fe;
    decBuf[7062] = 256'h5efecbfe54ff1900cf0076018b010201f6ff03fe27fcfbf985f8c9f8fef987fb;
    decBuf[7063] = 256'hb8fd2efffaffbcff14ff15fe8afd0bfde5fc7cfc1dfc01fc4ffc54fdd4fe3900;
    decBuf[7064] = 256'h21019f017901ca00edff97ff7dffc4ff3000b900cb00db007400acff6ffea0fc;
    decBuf[7065] = 256'h74fa69f815f7e0f518f617f715f9f1fa1dfd93fee7ff1c01c401f7012502fb01;
    decBuf[7066] = 256'h88012001c10031007aff75fe3bfd14fcbbfa76f94ff88ff727f746f710f863f9;
    decBuf[7067] = 256'h05fb1dfc1cfdeefc1bfc0ffb60fa80fa83fb02fd67fe4fff25ff65fe2bfd04fc;
    decBuf[7068] = 256'h44fb96fa76fa20fa06faeef9d9f9ecf946fa56fa47fab4f9dcf8d9f72bf7ccf6;
    decBuf[7069] = 256'h5cf747f8a3f944fbcdfcccfd57fe2dfe07fee4fdc4fda8fd8dfd17fdfefba4fa;
    decBuf[7070] = 256'h60f98df867f8cff86df9c4f912fafaf9b9f9cdf903fa74fabefa01fb6efbf3fb;
    decBuf[7071] = 256'hb7fcd7fd30ff1800960023002fffd3fd8ffc10fc37fc2bfdc6fe4f004e017c01;
    decBuf[7072] = 256'hfe003e0004ffddfdd1fc22fc45fb7cfac5f94ef964f93bfab1fb7cfda8ff1e01;
    decBuf[7073] = 256'hea01ac0174014101cc01f3024c044a069e0758081f08ec070507de05d1045103;
    decBuf[7074] = 256'h200115ffb1fc71fafcf8b8f87af893f95efb89fd2a00a402e304ef064308fc08;
    decBuf[7075] = 256'h340901092f09590933095609f7082e084307e70545044c0270003cff93fe92ff;
    decBuf[7076] = 256'hd700a6025604ff043205a704280402042504840413056205d9054506a706dc06;
    decBuf[7077] = 256'hac0627066205ab0435041f048104fe0491051a067306c506f106340758073707;
    decBuf[7078] = 256'h05077c06a405a204680341028101180138018e0179029603a304970535068b06;
    decBuf[7079] = 256'h0806d4045903f4016801e70140033e051a074f081708180777057d032902f500;
    decBuf[7080] = 256'hdcffa9ff7bfff9ff6c0060017d028a037e041c05ac05c605ae05eb04cc037302;
    decBuf[7081] = 256'hd10048ffaffe81fe57fecafe33ff100013014d02c803c7045205d3047a03d901;
    decBuf[7082] = 256'hc0008d00bb003a0160013d011e0101014f019701d7017501d4001200f8ff6e00;
    decBuf[7083] = 256'h880194024303620345036003d60399041c05d40490033501f5fe80fdb4fcf1fc;
    decBuf[7084] = 256'h9afd33febefee8fea8ffe200090262034a04c8048805f1058f061f076d075507;
    decBuf[7085] = 256'h1407b206ee059a04f9028f004ffedafc96fccafdc4ffb002a104fc04a9049e02;
    decBuf[7086] = 256'h4a019afff1fe8affcf004a0215044a058205e904010483031003780356041f05;
    decBuf[7087] = 256'h0a066906f9067b072208b9081b09e508f207e7054603cc008dfe81fc2dfb74fa;
    decBuf[7088] = 256'hacfa45fb8afcb1fd57ffe000ab025b04c4066008d509a10a640a4b09b2082708;
    decBuf[7089] = 256'h510877089a083b08ff068405b90384026c01d3004700c9ff09ffe6fec7fe56ff;
    decBuf[7090] = 256'h0d00e300e601da023604d705f0065508e008b608f60748072b068504fc029701;
    decBuf[7091] = 256'haf002d01d4023d052108130a220bd00a850a410a7f0ab70aea0a020a33088c05;
    decBuf[7092] = 256'h5d023a000fff00feadfdf8fd3cfe7afe92fff700f6025a0599073a0aff0b9a0d;
    decBuf[7093] = 256'h7a0ebe0e800ed80d3f0db40c350cc20bce0a7209740798056c0361019500dcff;
    decBuf[7094] = 256'h34ff67fff2ffc4001e021c048006c008cb0a1f0c5d0c240c250b8409fb073006;
    decBuf[7095] = 256'h8004d8033f0310038f039b04d5055007b5089d091b0aa809b408d7070e07f306;
    decBuf[7096] = 256'h0b074c0711074d06f904b4038d028101d2007400aaff28ffe0fe21ff48001702;
    decBuf[7097] = 256'h43044e061a07d3072b072c064405c604390573069608a20a6e0b300ba7091007;
    decBuf[7098] = 256'he103be01ccff72ff20ffd5fe91fe5cfd44fcabfb7cfbfbfbbafc3afe05003102;
    decBuf[7099] = 256'hd2044b078b09010bcd0b0a0c420ca90bc20af208cf05f6014dfdecf813f68ef5;
    decBuf[7100] = 256'h07f62af8e3fa11fe35005f016f020a048005d4060009750a410b040b0a091e06;
    decBuf[7101] = 256'h9f0254ff56fc2bfbd1fa23fb6efb3afc78fcb0fc49fdd4fd52fe12ffc0ff1f00;
    decBuf[7102] = 256'h76002c01320226030304e603c702d40070fed5fcf5fbc1fcecfef8005c039b05;
    decBuf[7103] = 256'he6052a0671055804f302f50091fe51fc1bf9f8f63ff430f3ddf228f36cf325f4;
    decBuf[7104] = 256'h3ef5d7f5d5f7c1fa08ff27045b0a860ecc101b10fa0cfe08550434017ffffafe;
    decBuf[7105] = 256'h91fd49fc90f962f663f3e4ef7bee0dee71ee35f075f2abf5aaf862fbdcfd1b00;
    decBuf[7106] = 256'h2702030437056f05d60492036e0163ff97fe59fe91fe2aff59ff86fee0fc77fa;
    decBuf[7107] = 256'h92f7a1f591f43ff48af466f616f82ff9c8f999f9c7f854f876f815f951fa23fb;
    decBuf[7108] = 256'h4afb56fa39f979f828f902fb76feb1026704eb048203a8ff00fb9ef6a2f214f1;
    decBuf[7109] = 256'h8df1d5f200f40ff5bdf472f4b6f470f5f8f629f935fb11fd45feeefe21ff4fff;
    decBuf[7110] = 256'h25ffb2fe78fdfdfb66f937f639f3f2ee1aec8cea14ea5ceb15ee8ef073f32bf6;
    decBuf[7111] = 256'h3bf7d6f84cfa28fc53fef400b902540409042d020aff31fb91f756f37df0e7ed;
    decBuf[7112] = 256'h7eec10ec3bed4aee41ef21f055ef20ee97ecfeebe6ec5eeff7f399f9e7fe5902;
    decBuf[7113] = 256'h3a04cb043502f9fdb6f78bf3c1efb0ed91ef6af200f55af7c8f7d6f512f476f2;
    decBuf[7114] = 256'h2cf2f8f2a8f4c0f559f615f5f1f250f0d7ed3cec5beb17eb4cec45eea9f032f4;
    decBuf[7115] = 256'h7df756fbedfd4700b4008affc5fde1fa61f717f4f3f102f0f2eefbedb1ede5ec;
    decBuf[7116] = 256'h2bec83eb50ebdbebffeda0f083f41af764fad2fa35fb26fae6f7dbf577f3dbf1;
    decBuf[7117] = 256'h66f022f05ff098f097f17ef251f3c4f35cf3c0f1e7ee2eecb5e9bee834eaa8ed;
    decBuf[7118] = 256'he3f103f775fa56fcc4fb3ffbc7faa3f879f71ef728f647f57bf4c2f339f2a2ef;
    decBuf[7119] = 256'h74ec75e9f6e59ce32ee392e30be639ea7cf052f6a0fb72005302c1012bffe0fb;
    decBuf[7120] = 256'h07f879f601f66ef660f8baf868f85df6f9f314f15cee4ced9fede9ed2dee74ed;
    decBuf[7121] = 256'h0bebcbe880e8d4e973ed2df498fa6e003001e001bffe2dfea9fd03000103f304;
    decBuf[7122] = 256'he30311ffdef85ef152ec92e968eaaeec1ff000f2b5f331f3a9f317f441f5bbf7;
    decBuf[7123] = 256'hfbf970fbc4fc7efd26febffe6000ca02ae0566082b0ad90938079f02fdfcaff7;
    decBuf[7124] = 256'hddf2fcf023ee96ec2cebbfea22eb9ced25f160f55cf9fcfc56ff5402d4051e09;
    decBuf[7125] = 256'hd30df410a9122512bc10980e190bce07f5034cffaaf95cf489ef68ecb3ea40ec;
    decBuf[7126] = 256'ha9eda8f060f3daf51af8bafa9efe3d02880586083f0b4e0c450d900d4c0d930c;
    decBuf[7127] = 256'h0a0bd90863070f064d068506b806d00558030bfe39f7a3f278ee32ec43eea5f2;
    decBuf[7128] = 256'hc5f797fcb9ffb5034b06a508c90a810dfb0f96114b116f0fd10b3108f603faff;
    decBuf[7129] = 256'h6cfe03fdbbfb1efce3fd7eff1f029804d8064e0882074d06540478023a027202;
    decBuf[7130] = 256'hd7031c054306030725078407db072908e207f4061905b50276006afe16fdd9fc;
    decBuf[7131] = 256'ha1fca0fd41ffaa0133057e08570cf70f51127414d81432153b14c612520f160b;
    decBuf[7132] = 256'h1a077a033fff66fcd9fa60faf3f91dfb97fd20016a044408d1093a0bcd0a300b;
    decBuf[7133] = 256'h210a730a280af40aa50c2e0e2d0fb80f8e0f810e8d0d700cb00b020be509f207;
    decBuf[7134] = 256'h1606eb030a034e038304ed068808680924096b08c207290758078207f5071808;
    decBuf[7135] = 256'h7708cd08ec09df0b430e2811191329143213bc11e00f300e170d180cd40a0409;
    decBuf[7136] = 256'h5d06e303480293025f038b0596077209220b1b0d7f0fbf1135137913c9117f0e;
    decBuf[7137] = 256'h430a6b07dd05650588077a09f30bea0c350d690c340b8c0a250bc60ca00f5812;
    decBuf[7138] = 256'hd214c815e8148412fb0ec00ae7074804cf033d0467059608940b4d0e1110ad11;
    decBuf[7139] = 256'hb8130c15bc164518de18f6177e155012760ed70a8c07690577031d03ca02ab03;
    decBuf[7140] = 256'h870537073009940bd40ddf0fcb124a1695196f1dfc1e741f511d0a19eb13180f;
    decBuf[7141] = 256'hb60a970525024400b2ff3700810311095f0ed111f2148415ff14a5128210570f;
    decBuf[7142] = 256'h480ef60dd60e2a10da11431483168e18e219a5193b17b313860e53087d02b3fe;
    decBuf[7143] = 256'h42fba1fa57fcf6ff31045109850faf13f5156719481bfd1c8b1e221d231a1615;
    decBuf[7144] = 256'he20e0d09bf03ae010d01e6038607d00aaa0e4011a9123c12830fa00bf706d603;
    decBuf[7145] = 256'h21029c01f603d007810dcf12a2178319f1184814e70f0e0d800be90ce80fa012;
    decBuf[7146] = 256'h4612bd0e9109be045d00cbff5801a3047d08130b7c0cea0cbf0b46096106a903;
    decBuf[7147] = 256'h990290035c07fb0a370fec1068100e0eea0bc00a650a5c0b3c0c700bc0095707;
    decBuf[7148] = 256'h6006ab060f09f30be40d3f0eff0bc908ef045902e0014e023f044f0546069006;
    decBuf[7149] = 256'h4c069305eb041e05a9052407ef089f0a480b150b2d0a0908fe0522047202e900;
    decBuf[7150] = 256'h1effe9fd21fe52001e04c608280ddd0e590eff0b4b07e90210007afd01fd6ffd;
    decBuf[7151] = 256'h99fe1301f703af067408c608e607fa0441027d002b00a00104044406ba07ee06;
    decBuf[7152] = 256'h47046300cdfd73fbe0fb99fe7c021c067608be09220ac709d008f00724077405;
    decBuf[7153] = 256'h9a02e2ffb3fc90fa2cfa87fa7efbc8fbfcfa4cf933f800f845f9bdfbebfeea01;
    decBuf[7154] = 256'h4d02a802fa02da032e055a07d0088c08d30769052a038900c4fe85fce4f96af7;
    decBuf[7155] = 256'hcff5eff443f6eaf883fde40104071509f60a640ad7087d067e03c60097fdbef9;
    decBuf[7156] = 256'h1ef6e3f10aef74ececec35eeedf067f3a6f587f6cbf608f7b1f7b0f8aefa12fd;
    decBuf[7157] = 256'hf6ffaf022805c3060e07420616047601b1ffbafe70feb4fefafd91fbbff6edf1;
    decBuf[7158] = 256'h4aec80e86fe650e84cecfef14cf75df93efbacfa15f8bbf598f36df2c8f2bff3;
    decBuf[7159] = 256'h34f510f7c1f84afa7bfc1bff95013003a604da0333019afcf8f6aaf138ee57ec;
    decBuf[7160] = 256'hc5eb5ceec5ef58ef2deeffea00e8d6e630e770e911ec8aee81ef36ef7aef2af1;
    decBuf[7161] = 256'h74f4a0f973fed502ad053b07b3076b067904b502d1ff18fd35f995f55af13aec;
    decBuf[7162] = 256'h67e746e491e215e37ee4a2e693e8eee89ce8bbe7efe6a9e712ea3fee5ff392f9;
    decBuf[7163] = 256'hbdfd0300b400d3fe90f8baf26cedfae99aea73ed1cf27df656f9d2f878f679f3;
    decBuf[7164] = 256'h88f12df124f22ff483f546f5bdf3c0f00beca9e7d1e431e1c8df80dee3dea8e0;
    decBuf[7165] = 256'h30e46ce88bedfdf01ff4d4f561f7daf722f986f9e0f945f83af6d6f396f120f0;
    decBuf[7166] = 256'h54ef9beef3edf4ecafeb88ea62eacaea29ebd3ea4be971e62be22fde98db20db;
    decBuf[7167] = 256'h68dce8df23e41fe8b6ea1fec43ee34f063f317f8b9fd0703180578049f01eefb;
    decBuf[7168] = 256'h1cf5dbec4fe748e488e1b3e0f1dfa1e0c0de2fdeaadd23de46e08de4d0eaa5f0;
    decBuf[7169] = 256'h6ff4e1f741f7aff622f5a9f417f57af5d5f5def4d3f2e7efa0eb81e60fe3eedf;
    decBuf[7170] = 256'h5cdff2e12ee62aeac0ec39edf0ebffe93ae8e8e75ee9c2eba6eed1efe0f08ef0;
    decBuf[7171] = 256'h43f00ff1bff209f663f887fa23faaaf721f4d6f0b3ee88ed2eeddbec66eb7ae8;
    decBuf[7172] = 256'hfae4a0e258e110e4f4e7a5edf3f265f646f8d8f84af7e1f599f4fcf457f54df6;
    decBuf[7173] = 256'h03f6bff50ef415f2c1f008f040f041efa0ed56ea2ae557e076de08df9fe1dae5;
    decBuf[7174] = 256'hfaeaccef2ef42af8dcfda6011805b805260587011e00d5fe39ff48009a00fafd;
    decBuf[7175] = 256'hacf8daf199e90de407e1f1e11ce6eeec2ff5bbfac6ff8602b1016bff5afd39fa;
    decBuf[7176] = 256'h83f8edf593f370f17eefbaed1eec69ec35ed61ef6cf1d0f310f61bf87ffabffc;
    decBuf[7177] = 256'h60ffd9011904240678073a072206f1035001d6fe97fc8bfa9ff7e7f4b8f195ef;
    decBuf[7178] = 256'hf8efbdf18ff6c2fc98026206120772069903faffa0fd57fc2dfbd2fa24fb6ffb;
    decBuf[7179] = 256'hb3fb6cfc85fdb6ff5702d004c7051206360413013afd9af940f71df5b9f414f5;
    decBuf[7180] = 256'h53f71ffbc8ff29042608bc0a440ad609730918090f0aef0abb0b020b09092d07;
    decBuf[7181] = 256'h01058b03bf0206025e01c5009600c1008001000365044d05cb0558051e04f702;
    decBuf[7182] = 256'hd102c503a0058c087d0a8d0b960a8b08af067a059206c308640b290d7b0d050c;
    decBuf[7183] = 256'hb10a8508100734050803670039fd3afad7f99bfbc8ff0c068c0d9c143219b21b;
    decBuf[7184] = 256'h741c631a41176914c9106f0e270d350b260ae607db0577038002a0016c021c04;
    decBuf[7185] = 256'h3505ce0542057004960416061309a20e6c127d14dd1304115c0c3b09a908360a;
    decBuf[7186] = 256'h810d5b11f1135a15ed14c213fe110711521196114f1217124c10a50d760a7807;
    decBuf[7187] = 256'h86057704c904140558051a055205b70612093f0d5f123117d41c1a1fca1f2a1f;
    decBuf[7188] = 256'h2e1b8516e310950b8409e308990a2f0d7a109d1201135b1352143215fe153c16;
    decBuf[7189] = 256'hb314b611270c5d084c06ec06c5095b0cb50ed81091130a169319de1cdc1f0721;
    decBuf[7190] = 256'hf71fb81dec194c161112380fa20c390ba60b0a0c190dc70ce70b1b0b580b510d;
    decBuf[7191] = 256'hc5101014ea17801ae91b7c1b511af719a4195a198e18d417bc16f11441132812;
    decBuf[7192] = 256'h8f11bd1138130315b416cc173317d814f411750e0c0dc30bee0cfd0d980f0e11;
    decBuf[7193] = 256'hea129a149316e7171c19e4187f17de1574133511940ecf0c340be90a3d0c600f;
    decBuf[7194] = 256'h1514b719051f1621f7221e20871d5b182812fd0daf08dc03fc016a01f7024206;
    decBuf[7195] = 256'h1c0ac40ee511be1455179f1a9e1dc81ed81f3c1e711ad1169612e110530fcb0f;
    decBuf[7196] = 256'h830e910cae080504a4ff12ff9f00bc063d0e51176b1d871e851d1917990f8908;
    decBuf[7197] = 256'hf3031e036405d608380d1010a71210147e14a815b816ae178f18d3189e173415;
    decBuf[7198] = 256'h5012d10e770c530af0094a0af80918093c0710059a034602090241020e028301;
    decBuf[7199] = 256'h040111021c047d08e111461b60217c227e23942214204a1c771794107e0619fd;
    decBuf[7200] = 256'hfff6abf3adf443f9c300ce058f086409260a370c580f5513f4164e19e0186115;
    decBuf[7201] = 256'h440fc407b4001efc9ef9e4fb56ff3906ce0af90ebb0faa0dc90b140a9009080a;
    decBuf[7202] = 256'h760a4b09d206a402a8fe1bfd84fe820102054c089509310922082b07e0061406;
    decBuf[7203] = 256'hd7052e0595040a04dd04d006bc09ad0bbd0c6a0cca099b069d03ab015101ec02;
    decBuf[7204] = 256'h62042e0574047b028fff9efdd9fbe2fa02fabef905f9cdf898fa36fedf028108;
    decBuf[7205] = 256'hcf0d4111e1112c10950d4b0a7106db039fffc6fc1ef8bcf3e3f056efbff0e3f2;
    decBuf[7206] = 256'hf0f7c3fc65022f064008210ab30a400ca90dcd0fbe116411240fc30ae0039ffb;
    decBuf[7207] = 256'h13f603ef43ec6eeb30ec41ee62f13bf4daf725fb49fd3aff4a00e501f003cc05;
    decBuf[7208] = 256'hf807d8089408e4060a0452018dffdfff5501b90354059f053b030effeef9bbf3;
    decBuf[7209] = 256'h90efc6eb76ec57ee77f349f86bfb43feda005201c0012302c90189ffe8fc6ffa;
    decBuf[7210] = 256'h2ff87af856fa79fd770069020e0217013700e3fea5fefdfd98fcf7fa8df84df6;
    decBuf[7211] = 256'hadf3e8f14df098f064f114f37df519f7f9f7b5f7fcf6e3f57cf6c1f7e4f91afd;
    decBuf[7212] = 256'h19000a021a03c802bc00d0fd8af98ef5f7f29df07aee4fed40ec49eb94eb70ed;
    decBuf[7213] = 256'h0ef1b7f518fa38ff49012a0398021402ab0062ff71fdf7fa13f85af577f1e0ee;
    decBuf[7214] = 256'h96eb72e948e838e78ae700e964eba4edafef8bf144f27df27cf31df567f8a2fc;
    decBuf[7215] = 256'h9e003e04c603c700f3fa1df5cfef5decbdeb72ed09f062f2d0f2a5f1e1efeaee;
    decBuf[7216] = 256'h9fee6befa0f0b9f120f122ef36ec7de9b9e754e920edd1f21ff891fb72fde0fc;
    decBuf[7217] = 256'h53fbe9f97cf918f9bef8c7f7bcf548f2fdeeffeb0deab3e905eae5eab1ebefeb;
    decBuf[7218] = 256'h27ec5aece5ec64ed8aed67ed48ed64ede7edbdeebfefb4f052f16ef1bdf104f2;
    decBuf[7219] = 256'h9bf273f33df4f3f43bf57cf505f611f7b7f840fa3ffbb4fa90f8c5f41cf0fbec;
    decBuf[7220] = 256'hffe868e6ffe491e4f5e4b9e69ee91ded59f131f4c8f64ff6e2f5b7f4a8f356f3;
    decBuf[7221] = 256'h75f221f1f6ee55ecdbe9e5e89ae866e9a4e9dce9a9e934eaafebacee86f225f6;
    decBuf[7222] = 256'h8ef7d7f801fac6fb05fea600b6011a00b9fbd6f46bee96e8d4e723e704e9b9ea;
    decBuf[7223] = 256'h3eebd5e967e9cbe9daea75ec16efdbf02df1e2f09ef057f150f3c4f60ffa0efd;
    decBuf[7224] = 256'h71fd17fdd7fa36f8bdf57df372f186ee06ebbbe798e56de47de5bde788eb1fee;
    decBuf[7225] = 256'h6af1b2f216f325f4c0f5f7f8f5fb3c001403a20439033a0066fae5f2daed6fe7;
    decBuf[7226] = 256'hefe4b1e5c2e764ed36f4ccf8f7fc3dff2cfd0afa0ef681f4f9f41cf70ef91dfa;
    decBuf[7227] = 256'h82f84cf572f1d3ed6aecfceb27ed36eed2efb2f07ef12ef397f5d7f74df919fa;
    decBuf[7228] = 256'hd2fa9afa67fa7ff9adf853f7b2f599f400f48bf45bf686f892fa6efca2fd4bfe;
    decBuf[7229] = 256'he4fe12ffe8fe75fe81fd25fce0fab9f9faf891f874f735f550f2d1ee86eb3eea;
    decBuf[7230] = 256'hdae9eaea2aed35ef11f13df348f5bcf806fc05ffbd011802c6017b0137017501;
    decBuf[7231] = 256'h1d025002680145ffa4fc2afa46f755f590f350f1dbef0fefd1eecaf0b6f335f7;
    decBuf[7232] = 256'h80faa4fccefddefe7900ef01cb037b05b305b404fc01b6fdbaf923f7baf527f6;
    decBuf[7233] = 256'hc4f51ef683f478f224f1e6f050f321f855fe2a047809ea0c8a0df90c620a1807;
    decBuf[7234] = 256'h88013afc07f6dcf112ee61ed42ef3ef3def629fa4cfcb0fc55fc5efb14fb68fc;
    decBuf[7235] = 256'h18fe8100c102cc0420065507fd07fc08410abc0b210d660e900ed00dc50bf907;
    decBuf[7236] = 256'h5103aefd60f88ef36cf0dbef5ff0c8f1ecf3ddf557f897faa2fc7efeb3ffebff;
    decBuf[7237] = 256'hb8ff430015016f02100429052806c907330a600e80135218731bbe191615330e;
    decBuf[7238] = 256'hc80747003cfb51fad1f793f844f9a3f812f88df715f782f7adf8dbfbb5ff5403;
    decBuf[7239] = 256'h9f06e70712096c09080b130d770f5b124d145c150a159413b811110f970c0f09;
    decBuf[7240] = 256'hc4050f01aefc8ef71cf43bf2aaf149f584f9c8fff3034109520b730e2810b611;
    decBuf[7241] = 256'h1f1367147612470f930a31063502b00119033d05f507ba096809f20716065d05;
    decBuf[7242] = 256'h950560071009090bd50b970bd00bcf0c700ef90f5e118c110e110110c70ef50d;
    decBuf[7243] = 256'h820dbc0b15097c04dafe10fbfff89ff99cfd4402e6072c0a3d0c5d0aa7081a07;
    decBuf[7244] = 256'ha206ea07a30a860e26127015de157a156b14cf12851241127e12b712ea12a511;
    decBuf[7245] = 256'h810fb60b0d07ab02d3ff4effc6ffea01a204670602084d08a109cd0b030fdc12;
    decBuf[7246] = 256'h7315eb157e155314441396137614421505159b12120fd70adb064404cc031405;
    decBuf[7247] = 256'h7805d2058005cb050f064407ad09ed0bf80d4c0ffc101512e01387164c18e719;
    decBuf[7248] = 256'h07191b160d11da0aaf0669041905fa06f60a8d0de70f5410b810121164114512;
    decBuf[7249] = 256'h0112cc10630e230cad0a790b200e4f114d143f16e415a5136e10950cfe09a407;
    decBuf[7250] = 256'h81058f0335033e02890255038a04f306d709570d83125617771a091b841a3917;
    decBuf[7251] = 256'h6013c00f670d1e0cbb0b150cc30be30a170a5d09060a370c6d0f6b125d140214;
    decBuf[7252] = 256'h6712310f0d0de30b3d0c7d0e8810dc11a810ce0d8809680495ff74fcbffa4cfc;
    decBuf[7253] = 256'h8800cb064b0e5b15c61bf11fb3200320e11c091a69163d116a0c09080c047601;
    decBuf[7254] = 256'hfe0046023804b1064c089708530891081a0ab10cdf0fde12cf14c0132412840f;
    decBuf[7255] = 256'hbf0d110e1d10f911b21229112c0ec2072c0301ff3ffe500031020a05a908f40b;
    decBuf[7256] = 256'ha8100a152a1a3b1c9b1b9e17ed119f0c2d09cd09a60c4510af118b0f450b2506;
    decBuf[7257] = 256'h520131fec3fe5000aa02ce04f8055306a506f006bc077508ad08e008c809430b;
    decBuf[7258] = 256'hda0d5310381362140814c811bd0fd10cdf0a6608ca06bf04f3033a0372030b04;
    decBuf[7259] = 256'h960469052906a8077309240b3c0c6f0cce0ad50871067a052f0573052c06d506;
    decBuf[7260] = 256'h0807d9065b06e805f4045604c6037803ee03dc04ba059d057d043e025affa1fc;
    decBuf[7261] = 256'hddfae6f931fa85fbb0fde700c00460089b0c740f01117a113110400e7b0c9709;
    decBuf[7262] = 256'h1706dc01e0fd40fae6f779f731fa15febd02df0594070f07a60583035802fe01;
    decBuf[7263] = 256'hf4020005dc0695075d07f8059d031400d9fbddf746f5ecf2a4f1cef2def31df6;
    decBuf[7264] = 256'hfef6caf783f89cf999fc28027607a90dd4111a14cb14ea1211107b0d3f094305;
    decBuf[7265] = 256'h92ff44fa71f550f2bef14bf396f695f94dfcc7fe6200d8012c03690331033202;
    decBuf[7266] = 256'h340048fd90facbf879f8c4f8a0fa59fb21fbf0f84ff6d5f33af21af38ef6cafa;
    decBuf[7267] = 256'ha3fd4201ab02190343049e049405df051305e7021cff73fad1f407f195edf5ec;
    decBuf[7268] = 256'h87ed26f152f625fb87ff830319067308bc09e60a8c0a4c08eb0348fefaf866f1;
    decBuf[7269] = 256'h5becc5e745e583e434e514e7ede98dedc8f1e8f65afa7bfd30ffbe003601c800;
    decBuf[7270] = 256'h10fe96fb0ef8b4f590f366f2c0f2b7f397f4ebf5a5f6ddf6aaf67bf6fdf570f6;
    decBuf[7271] = 256'haaf722fa50fd4f00400250035902b8ff8afcb0f81af6cff2f6ee4deaebe5efe1;
    decBuf[7272] = 256'h59dfe0de04e183e4bfe8bbec5af0b4f2d8f43bf596f544f563f41ff4d9f4d2f6;
    decBuf[7273] = 256'h46fa81fe7d021d0677082e07e802c8fd95f7bff179ef68ed49effef08bf204f3;
    decBuf[7274] = 256'hbbf1caef9becc2e822e5d8e1b4dfc3dd1dde14dfe0e291e863efcef5a4fb6eff;
    decBuf[7275] = 256'h1e007effc9fd3bfcd2fa65fac8fa6efad2f832f603f305f085ec2bea08e8a4e7;
    decBuf[7276] = 256'h4ae741e8f6e73ae8fce7a4e8d5eaa1ee4af3abf7a8fb35fdbdfc99fae1f767f5;
    decBuf[7277] = 256'hccf3ecf220f267f1deef79ee91edbbed14ef59f083f02aef72ec9ee673e2a9de;
    decBuf[7278] = 256'hf8ddd9dfb2e251e69ce9bfebb1ed2af06af236f6d5f911feea0077020e01c5ff;
    decBuf[7279] = 256'h0dfd93faaff7f7f413f162eb14e641e120de8edd1cdf57e377e8aaeed5f29ff6;
    decBuf[7280] = 256'hb0f850f9e2f955f8ebf6c8f448f1feedffea0ee9b3e861e841e90dea4bea83ea;
    decBuf[7281] = 256'h1ceb4beb75eb02eb99ea3aea57ea42eb1ced90f0dbf3b4f754fbaefdf6fe2100;
    decBuf[7282] = 256'h11ff76fdaaf902f5a0f0a4ec04e98ce8d4e98dec06efa2f0ecf030f177f0aff0;
    decBuf[7283] = 256'he2f011f1e7f027f0edee72ed0dec82eb57eb7eebe6ebc4ec73ee1af194f3d4f5;
    decBuf[7284] = 256'h49f78df750f737f604f68ff60af809f994f916f923f7bff424f3aef1f2f127f3;
    decBuf[7285] = 256'hcff368f4ddf362f263f135f1b0f2adf586f926fd80ffedfffcfdcdfacff74ff4;
    decBuf[7286] = 256'h04f1e1eeefece0eb8eeb43eb0fec4dec85ec84ed25ef6ff29bf7cffda403f208;
    decBuf[7287] = 256'ha30902094d07ae03540130ff3ffd10fa37f68ef12ced54eacfe938eb37ee7df2;
    decBuf[7288] = 256'h56f5edf746fab4fadefbeefc40fd8bfd47fd8efc56fceffcd6fda6ff5601df02;
    decBuf[7289] = 256'h12032a02b2ffcffb26f7c4f2c8ee3bedb3edfceeb4f1e3f4bcf85cfca6ffa502;
    decBuf[7290] = 256'h96045b06f607d6081a09dc0854075704c7fe79f9a6f4c6f257f3eef51afbedff;
    decBuf[7291] = 256'h0e03e7056b060205040284fe2afce2fa45fb0afda5fe1b00d7ffa2fea9fcddfb;
    decBuf[7292] = 256'h1bfc84fe0d024806fd078b091209ca07d805140479020301bf00fd008602b704;
    decBuf[7293] = 256'hc2069e08dc08c307f805cc0356028a01c80151031c054807e909620ca20e4311;
    decBuf[7294] = 256'h52125b11bb0e6d091f04ecfdc1f97bf72bf8cbf881fa17fd71ff7002ef052a0a;
    decBuf[7295] = 256'h030da3101b11ae10f50d7c0b97086d073109160c5c105814e6154f1706164e13;
    decBuf[7296] = 256'hd410950e890c250a41078904c402cd01ae029a05e009b90c460edd0cba0ac808;
    decBuf[7297] = 256'hb9070b08160a6a0ba80b8f0af807ca0481031e032d041207ca09440cdf0d550f;
    decBuf[7298] = 256'ha910d412e014cc17bd19cd1ad619a016eb11890db10a23099c09bf0b780e3c10;
    decBuf[7299] = 256'h8e10190fb50c750a6a081607e105380505053405af06e008160c150f0611cb12;
    decBuf[7300] = 256'h1d136813241361139a1367137f12af10ff0ee60d4d0d7c0d520ddf0cea0b4c0b;
    decBuf[7301] = 256'ha30b2a0d0410f61150121010af0b4d077504f0033b07140bc61090140218e219;
    decBuf[7302] = 256'h741af01986186316711443111f0ff50de50c930cb30be70aa90ae10a460cfe0e;
    decBuf[7303] = 256'h7d12d714fb169716d3149312c70e310ce608c306d104c2036f0350043c07bb0a;
    decBuf[7304] = 256'hf70ef3128915e3175118ed1793179c1651160d164b168316b61688160916b014;
    decBuf[7305] = 256'h0f13a510c10d080bda07db04ea0225012f00a401900410084b0c4810de123815;
    decBuf[7306] = 256'hca1467145713051350131c14d5147e157f1424129b0e600a6306cd035403e702;
    decBuf[7307] = 256'h1104d60571077c09680c210f9a11da13ba14761442132912f61181125413c713;
    decBuf[7308] = 256'h5e13c311ea0e6a0b1f084604af014600d9ff75ff3a017a03b006d308c50a1f0b;
    decBuf[7309] = 256'hcd0a820a3e0a730b6c0d58101113201417153714e312291281114e11d9115812;
    decBuf[7310] = 256'h3112f7107f0ee709450473fd32f5def1d7eec2ef98f56afcaa046e0c7e131418;
    decBuf[7311] = 256'h941a561ba61a051a2d1796142d130911180f9e0c1609cb05f2016400fbfe8dfe;
    decBuf[7312] = 256'h2afe84fe7bffc6ff92004b01f4018d021803e7040a08e30b8c10ad133f14c314;
    decBuf[7313] = 256'h4b14dd134114e6139413f3105b0cb906e7ff26fda6fae4f995fa75fc07fd8cfd;
    decBuf[7314] = 256'hf5fe18019804e207060a300b8b0bf0097a082607e80691075c090c0b440bdf09;
    decBuf[7315] = 256'h27071a02a8fe87fb3cfdd2ffff04d109f20ca80e110cb709de054703cf028601;
    decBuf[7316] = 256'h23015eff68fe87fdcbfd7cffe501c90482079108e408990855089c078306b804;
    decBuf[7317] = 256'h1102e2fe09fb69f70ff5a2f4ccf546f8cffb19fff3028905e3075108b4085a08;
    decBuf[7318] = 256'h630783063f06010639066c068405b5030d012afd93fa2af998f9c2fa87fcd9fc;
    decBuf[7319] = 256'h63fbfff8c0f6dff5abf6cef9cdfc85ffe0ff8dffadfe69fe1900f302ab052508;
    decBuf[7320] = 256'h7708970733054f0296ff1dfd38fa80f706f522f231f0d6ef28f034f298f420f8;
    decBuf[7321] = 256'h6bfb6afe2201e702dd032804e403a603fe02ff01ba003fff74fd48fba8f8e3f6;
    decBuf[7322] = 256'h48f5fdf4c9f579f773f9d7fb72fdbdfd79fdc8fbcff96bf7d0f5f0f434f568f6;
    decBuf[7323] = 256'h81f71af8ecf719f70cf6a4f542f6f1f798fa5dfc54fd09fd3dfc7bfc23fdeefe;
    decBuf[7324] = 256'h2300cb0066ff0bfd27fa6ff7aaf50ff4c4f380f3bef3f6f3c3f3f1f373f300f3;
    decBuf[7325] = 256'h97f278f2b4f3d7f50ef90cfcc5fed4ff82ff77fd13fbd3f832f66ef477f397f2;
    decBuf[7326] = 256'h53f21ef176f0ddeff5eecbeef1eee5ef41f19cf380f639f9b2fba9fc5efc82fa;
    decBuf[7327] = 256'h56f84bf6f7f4c2f3aaf2abf120f1a1f014f194f25ff40ff698f7fdf82bf956f9;
    decBuf[7328] = 256'he2f834f817f70bf65cf5bef42ff4dbf223f0a4ec68e86ce4d6e14ee24de5cce8;
    decBuf[7329] = 256'h07ed04f1a3f4eef7ecfa6cfec6000e02ab0131ffa8fb6df771f3daf071ef04ef;
    decBuf[7330] = 256'h2ef089f036f056ef7aed45ec9deb9cec3dee37f013f2ccf204f337f365f38ff3;
    decBuf[7331] = 256'hb6f393f334f36bf280f121f177f162f2fdf3f6f5d2f707f93ff9a6f862f7e7f5;
    decBuf[7332] = 256'he8f4a3f37cf289f09dede5eab6e76ee60ae6cfe7b3ea6bed30efcbf0abf1fff2;
    decBuf[7333] = 256'h2bf5ccf745fa3cfb87fbabf97ff7def41af323f26ef23af3f3f32bf492f34ef2;
    decBuf[7334] = 256'h7ef0ceee26ee59ee41ef64f16ff34bf505f6cdf5cef42cf3a3f172ef67ed03eb;
    decBuf[7335] = 256'h68e9f2e7aee767e860ea4cedccf017f4f0f77ef9e7fa79fa4ff98af7eff50ff5;
    decBuf[7336] = 256'hcbf48df4e5f380f225f0e5ed6feca3eb65eb7eec7dedc2ee3df0a2f1a0f304f6;
    decBuf[7337] = 256'h44f8b9f9fdf944f92cf82df745f672f5fff40bf470f277f09bee66edbdec24ec;
    decBuf[7338] = 256'hf6ebccebf2ebe6ecc1ee35f270f66cfa0cfe75ffbe005a0096fefafceffa03f8;
    decBuf[7339] = 256'h4bf5d1f236f156f012f058ef40ee75ec40eb98ea31eb2feda3f0def4daf87afc;
    decBuf[7340] = 256'hc4ff0d01fe0259036202ec0010ff69fcf0f954f874f730f7e9f772f971fafcfa;
    decBuf[7341] = 256'h7efad8f86ff68af399f13ef191f19cf388f679f889f937f92bf7d7f51ef537f6;
    decBuf[7342] = 256'h68f808fb37fe5a004c02a60254020902b50081ff88fd24fb88f913f857f810f9;
    decBuf[7343] = 256'h99fa98fb23fca1fc14fd4efe1e00ce01c7031b05500668070108d30704066502;
    decBuf[7344] = 256'hb4fce2f577efa1e95be76ce9ceed11f4e7f9b1fd2301c3015502e2034b054a08;
    decBuf[7345] = 256'hc90b140f371162125211130f720c43094506fe0102fe5af9f8f41ff2a4f2fdf4;
    decBuf[7346] = 256'hb2f914fe100294022b0108ff16fd71fdb1ffe702e5059e08ad09b708d6070a07;
    decBuf[7347] = 256'hcd06750774085c0986091309640848073b061806770607072107da069505f403;
    decBuf[7348] = 256'hdb0242022a03a5040a06f206c806bc053c043d03b2028802ae025c0379041f06;
    decBuf[7349] = 256'h1808040bbd0d810f7810c310f70fc20e390d6e0b4209cd07f105bc04a303a402;
    decBuf[7350] = 256'h6001e100080187021e054d084b0b3d0d970dea0d9f0d5b0d990d410e740e460e;
    decBuf[7351] = 256'h1f0d790bf0095709cc08f608cf08ac084e0831087f08b4092f0bfa0c2f0e470f;
    decBuf[7352] = 256'h7a0f4c0fce0e5b0e660d4a0c3d0bd50a330b700c970d560ea80dce0b6a092a07;
    decBuf[7353] = 256'hb405e804aa04e3044a0478044b058a076e0a270da00f9710b70f630e2e0dd70d;
    decBuf[7354] = 256'h08103e131717ae19081c9a1b701aab186b1660140c135c11d30fa20d010bd307;
    decBuf[7355] = 256'hf903630109ffc0fd5dfd6cfeac004d03c6050608110a750c6c0d4c0e080ecb0d;
    decBuf[7356] = 256'h730e720fcd11b1146a172e19251ada198618cd1725178c165d1636154313cf0f;
    decBuf[7357] = 256'h850cd007af04fa026c01e5012d039103a00497057706cb07f7092d0d2c10e412;
    decBuf[7358] = 256'ha91444168f164b169115e91484138611120ec70a1306f20219009d0006020505;
    decBuf[7359] = 256'h4b096b0edd11be137315ef1476140914de12841231125111750fc50dcc0b6809;
    decBuf[7360] = 256'h2807b205e6042d04d504d405190794085f0a0f0c090e6d105113421507175917;
    decBuf[7361] = 256'h0e17ba1586148c123811880f8f0d2b0beb08e0060405cf03460247016000e1ff;
    decBuf[7362] = 256'h54008e0109033a054607320ab10dfc10d5147518de194b1a5a187614ce0f6c0b;
    decBuf[7363] = 256'h7007e2056a05b206dd07a109980a780b340bf70abf0a8c0a5d0a330a73093908;
    decBuf[7364] = 256'hbe06590571049f0378039b03bb03d80326046d0430051b06f8068807a2072b07;
    decBuf[7365] = 256'h940659068f0683074809f80a810c1a0dec0cc50b1f0a2608d206210598033302;
    decBuf[7366] = 256'ha8017e018b020a046f05fb052805cf032d02a4000b009600690176026a030804;
    decBuf[7367] = 256'h5e0478043104f003b5035c030b03a30210028701e600a500e000810144022f03;
    decBuf[7368] = 256'hcd0396044d05f3058b069e06da058604e5025c012901b4018602ad0273014fff;
    decBuf[7369] = 256'haffc35fa3ef9f4f8d0fa80fce9fe29019f02f3033004f803f902b5018e001b00;
    decBuf[7370] = 256'hf8ff96005f01e20159026e020c026b017d0021ffddfd0afd31fd25fe41ff4e00;
    decBuf[7371] = 256'he5ff4afee1fbfdf8d2f72df811fb90fecc02810405059c03790187ffc3fdccfc;
    decBuf[7372] = 256'h81fc2dfb7df9f4f7f5f6c7f6eef7e1f9bdfb6dfd15fe48fe77fef5feb5ffef00;
    decBuf[7373] = 256'hc1013402cc01af0009ff10fd34fbfff957f98af9b8f98ef91bf96df88ff7fff6;
    decBuf[7374] = 256'h49f6d2f591f57df5faf5eef6f9f830fc53fe45005401a601c600faffc5fe1dfe;
    decBuf[7375] = 256'h1efdd9fbb2faa6f9f7f817f934f94ef9a8f863f765f589f34bf3d4f405f73cfa;
    decBuf[7376] = 256'h3afd65febffec8fd53fc77fa42f90af93df925faa0fb9ffc2afd00fd5afbf0f8;
    decBuf[7377] = 256'h0cf61af456f24df3c2f436f881fb80fe710062ffc6fd90fa92f7a0f5fbf53af8;
    decBuf[7378] = 256'h46faaafcfcfc1cfc40fa0bf962f861f960fb4cfe3d004d0156004bfed7fa8cf7;
    decBuf[7379] = 256'h8df49cf2d7f02af174f140f275f36ef5d2f7b7fa6ffde9ff3b00c5fee9fc42fa;
    decBuf[7380] = 256'h7df8d0f8b0f914fcaffdfafda6fc7afa44f720f5f6f350f447f552f71ef8d8f8;
    decBuf[7381] = 256'h10f977f848f8c7f83af9a2f983f92df976f8fff715f8ecf829faa4fb3dfc6bfc;
    decBuf[7382] = 256'h99fb3ffa57f9d9f8fff868f988f931f912f86cf6e3f47ef3f3f21df3ddf3d1f4;
    decBuf[7383] = 256'h30f54df532f54af58bf58af60af8d5f985fb0efd0dfe98fec2fe9cfe79fedbfd;
    decBuf[7384] = 256'h12fd8afb20f93cf684f3bff16df1e3f247f52bf81cfa77fa80f9a0f8d4f796f7;
    decBuf[7385] = 256'hcef7cdf8b5f933fac0f986f8b4f7f4f617f7f4f730f957fa17fbaffa53f9b1f7;
    decBuf[7386] = 256'h48f5adf3ccf288f242f35af459f541f668f70ef907fb6bfdabff2101ed013401;
    decBuf[7387] = 256'habffe0fd2ffca7fa42f9fdf72af704f76df789f8e3f96efa98fad8f9e4f8c7f7;
    decBuf[7388] = 256'hbbf6f5f4c9f229f0afedb8ec99ed85f092f565fac7fe7c00000197ff74fd49fc;
    decBuf[7389] = 256'h3afb8cfbd7fba3fc5cfd24fd25fc83fa8af836f77df625f7bef74af874f801f8;
    decBuf[7390] = 256'h98f7f7f7c0f8dff9ecfa0ffb32fa2ff93bf85af85df997fa6afb43fb09fa3af8;
    decBuf[7391] = 256'h05f75df6f6f6def705f978f99bf93cf91ff905f91df907f9a5f828f854f7c5f6;
    decBuf[7392] = 256'h42f62af66bf6f5f6ddf739f97dfa4dfc82fd0aff09004e01c9022e0473054905;
    decBuf[7393] = 256'hef0338012afc58f7b5f16fef5eedfeed90ee15ef7ef0a1f221f66bf96afc22ff;
    decBuf[7394] = 256'h3200e0ff6afe8efcd5fb9dfb36fc1dfdf0fd7dfd89fceefa65f966f894f8bef8;
    decBuf[7395] = 256'h7ef92dfacbfae7fa36fbadfb44fca6fcdcfc8afc06fc65fb24fbc2fa68fab6f9;
    decBuf[7396] = 256'hb0f8bcf71ef73bf75af800fafafbd6fd0aff930092017a02f802d202980120ff;
    decBuf[7397] = 256'hf2fb18f879f43df065edd7eb50ec98ed18f153f573fa45ffa70380060d089507;
    decBuf[7398] = 256'h4c06cd0282ff84fc59fbb4fbf4fd69ffadff79fe9ffb1ff8c6f558f54af778fa;
    decBuf[7399] = 256'h77fd2f008a0093ffb3fe5ffd21fd59fd8cfdbafd3cfd2ffcb0fae5f8b0f708f7;
    decBuf[7400] = 256'h6ff640f66af691f685f75ff9d3fcff01d206f309a80b1b0ae005c0004efd6dfb;
    decBuf[7401] = 256'h22fdb9ff220190019effbbfb1bf8c1f52ff620f804fca3ffee023604d303c302;
    decBuf[7402] = 256'hcd01ec00a800efffd6fe71fd73fb1ffae2f96afb01fe300153034505ea049804;
    decBuf[7403] = 256'h220356029402cc0299020e0293002eff46fe70fe16008002c0040a05b6038b01;
    decBuf[7404] = 256'h54fe56fb2bfad1f96cfbe2fc46ffe100ec025005ec06f708c3098509dd08de07;
    decBuf[7405] = 256'hf606230663056f045303600184ff58fd78fc34fce4fdbe003d048807ab090f0a;
    decBuf[7406] = 256'hff08bf061f04f000cdfea2fdfdfd4ffe5a003602e6036f05d406bc07e6070d08;
    decBuf[7407] = 256'h3008d107b4073107ea06d4063707d70744080908fd06bd047d0207013b007001;
    decBuf[7408] = 256'h690345057a06b206e506b706e10607077007900700071506f80438041504b304;
    decBuf[7409] = 256'hb60536070109b10a3a0c9f0d870eb10e8b0edc0dff0cfc0bc20af308c7062604;
    decBuf[7410] = 256'h6202c70051ff95ff4e006701cc026d04f6055b07430815098909f1098f0a590b;
    decBuf[7411] = 256'h440c210db10dcb0d840d180d670c910bc80a450a5d0af40a1b0ced0c610df80c;
    decBuf[7412] = 256'h5d0b64098807d705bf04c0033503b6024302660204034004bc05ed07f8095c0c;
    decBuf[7413] = 256'h9c0ea710fb11391290112b102d0e510c1c0be40a4b0a6309e807b70516039d00;
    decBuf[7414] = 256'h02ff21feedfe9e000703a204ae068a083a0ac30b8e0d3e0f37111313cc139413;
    decBuf[7415] = 256'h2f123110450d8d0a1308d3055e040a03d5019d019c029a040e08580ba10c040d;
    decBuf[7416] = 256'h400ba509990755070f08b708500968089906e904600393031e04f00464058605;
    decBuf[7417] = 256'he8040505f005cb07b70a6f0de90f841139116d10bd0e340dcf0b2e0a15091608;
    decBuf[7418] = 256'h7506ec04bb024501010136029f042808820aa50c090dae0c5c0c7c0b380bfa0a;
    decBuf[7419] = 256'h520aed08ee068a044b026a012601e001f802c304f8058107e6082b0aa60b0b0d;
    decBuf[7420] = 256'hf30d1d0e5d0d230cff098a08ae0670063806d1065c078607c606d205f5046504;
    decBuf[7421] = 256'h16042e04ed0364030b03fa027f038b047e06d2070709af09e2096d0a970a570b;
    decBuf[7422] = 256'h060c650c480cc50bef0aed09f908dc0783063e05c3035e0219019b007400dd00;
    decBuf[7423] = 256'h3c015901a701bf012b0203037904440678072108ee07a906da04200459045805;
    decBuf[7424] = 256'h5607aa086309bb085607b4059c04690497046a05dd054506a406c106db06f306;
    decBuf[7425] = 256'h0807ce0650065d05dd03780233016100d4009902c504d006ac086f08e6064f04;
    decBuf[7426] = 256'h200122fef7fc9dfc93fd74fec8fffc0015027a03d505b908ab0a6f0cc10cb60a;
    decBuf[7427] = 256'h5208c90470024c00e9fff800ef01650331046e04c6036102c00037ff9efe6ffe;
    decBuf[7428] = 256'heefeaeff5c0039013c0230038c04d105a3061607f4065506c6050f056904fc03;
    decBuf[7429] = 256'h4c0347020d01e6ff8cfea5fd26fd99fd48fee3ff6c016b023c02c10090feeffb;
    decBuf[7430] = 256'h76f924f96ef9d2fb12fe48016c035d056d061b06a50441020100f6fd2afde3fd;
    decBuf[7431] = 256'hdcff4002dc0326045a03aa01b1ff5dfe28fd80fce7fb5cfbddfab7fa65fbc1fc;
    decBuf[7432] = 256'h63fe5c00b001ed0126028d01a5002600b3ff4bff6dfebefc92fa5cf75df4a5f1;
    decBuf[7433] = 256'h4af19df112f3fef5b7f830fbccfc41fe95ffca00e30148038c040b053105c904;
    decBuf[7434] = 256'heb037502aa0003fe8afb4af93ff773f635f6ddf6dcf77ef996fa95fb20fc9ffc;
    decBuf[7435] = 256'h2cfcc3fb28fa2ff853f6a3f48af357f3e2f309f562f604f88df9f2fa36fc5dfd;
    decBuf[7436] = 256'h1dfe86fea5fefbfe4afff0ffb300cd002700e2fe2bfce4f70bf57ef305f34ef4;
    decBuf[7437] = 256'h78f588f6daf68ff6c3f50af5d2f46bf553f67af786f87bf919fa6ffabdfa34fb;
    decBuf[7438] = 256'ha0fbb4fba2fb10fb5ffab9f94df912f947f999f91dfa53fa84fa1dfa54f9def7;
    decBuf[7439] = 256'h79f6d8f44ff31cf3eef218f38bf3aef38ef338f31ef365f3fcf3adf453f516f6;
    decBuf[7440] = 256'h01f7def71bf996fa61fc95fdaefe47ff75fff7fe84fed6fd7afc35fb66f9b5f7;
    decBuf[7441] = 256'hbcf5e0f330f2a7f0dcee23ee7bed48ed76ed49eea2efa0f104f4e8f6a1f965fb;
    decBuf[7442] = 256'h5cfca7fcdbfb22fb09fa70f9e5f8bbf8e1f84af9a9f9fff9e5f93ef925f8ccf6;
    decBuf[7443] = 256'h87f560f43af45df4fbf48bf571f59bf45ff3e4f14bf1d6f1a5f34cf630fac6fc;
    decBuf[7444] = 256'h20ff8eff2affb1fcccf914f74ff5b4f3d4f290f2cef296f2c9f29af219f3d8f3;
    decBuf[7445] = 256'h12f539f693f7d7f856f9c9f931fa51faa7fac1fad9faeffadbfac9fa98fa14fa;
    decBuf[7446] = 256'h2bf9cff72ef6a5f440f3fcf1d1f1f8f160f2fff201f4f5f4d3f50ff78af8eff9;
    decBuf[7447] = 256'h91fba9fc42fd14fdeafc77fcc8fb69fbdafa23fa4df911f8eaf644f52bf42cf3;
    decBuf[7448] = 256'ha1f223f296f2fef29cf39ff4d9f554f71ff94bfbc1fc9dfe56ff8efff5feb0fd;
    decBuf[7449] = 256'h35fcd0fa2ff9a6f7a7f6bff5edf42df47ef35ff328f4b0f589f842fbbbfdb2fe;
    decBuf[7450] = 256'h67fe13fde8fadcf800f747f60ff642f6cdf6a0f7acf8e6f961fbc6fc52fdd0fd;
    decBuf[7451] = 256'h5dfd69fc8bfbc2fa3ffa57fac3fa25fb37fbc6fae8f94df8c4f6c5f597f56df5;
    decBuf[7452] = 256'he0f549f6e7f6b0f7cff875fa6ffc4bfe7fff2800f5ff6aff97fe71fe93feb3fe;
    decBuf[7453] = 256'h09ff87fe22fdf1fae6f882f6e7f432f576f526f73ff83ef96cf942f968f9d1f9;
    decBuf[7454] = 256'haefa24fc89fd2aff4300dc00c401eb025e038103a302f400c8fe28fcaef96ef7;
    decBuf[7455] = 256'hf9f5b5f577f51ff61ef763f88af996fafffa1ffb75fb2cfc60fddcfe41008501;
    decBuf[7456] = 256'h58027e021602f900a0ff5bfe88fdaffda3fe3e00c7016002d5010500dafd64fc;
    decBuf[7457] = 256'h20fcd9fcf2fd25fe3dfd19fb78f869f7bbf731f91dfcd5fee5ffeefe0efe42fd;
    decBuf[7458] = 256'h80fd79ffdd011d0492054e0595040c0341010c00f4fe5bfe89feb3fec0fffa00;
    decBuf[7459] = 256'hcc018c02af025002c1013e0198002c00a2ff49ff18ffcefe71fed3fde5fc47fc;
    decBuf[7460] = 256'hf1fba8fc0cfe3d0048022404d4057d06b006de066006ed053e05610498037e03;
    decBuf[7461] = 256'hf403b7043a05f204ae03530113ff08fd3cfc7afc73fed7007202e8031c03e701;
    decBuf[7462] = 256'h5e00f9fecbfef2ff31021605ce079309890ad40a900a520a1a0ae7095c098d07;
    decBuf[7463] = 256'h610556037a01c100d901d8021d049b042804ee02c70107012a014702ed03e605;
    decBuf[7464] = 256'h3a07f307bb078807fd06d605ca04d603f802db025e03c2048d063e08c6095f0a;
    decBuf[7465] = 256'h8e0abb09fb089308340851086b08530812088907e8065006c7054a05f904ea04;
    decBuf[7466] = 256'h4805fd0585070e090d0a520b7c0b560b1c0aa108d606aa043403f002b202cb03;
    decBuf[7467] = 256'hca04b205300657067906d80668078708e109250b4c0c0c0dbb0dda0dbd0d3b0d;
    decBuf[7468] = 256'h950cfd0b4d0ba60ab8095d085e068204d2022a025d02a1031d058206c607f007;
    decBuf[7469] = 256'h1708f4079507b2079807df0776087509f50ac00c700e890f2210f30fcd0e260d;
    decBuf[7470] = 256'h2d0bd909a5088c07590771069e05f8036f0270014201bd0254058308810b730d;
    decBuf[7471] = 256'h180d210cac0ae009a2094a0ae30a6e0b440bd10a9709c508b807c4062606d005;
    decBuf[7472] = 256'hb505fd05bf06df07eb08df097e0ad40a220b3a0ba60b080c3e0c6f0c250c920b;
    decBuf[7473] = 256'hba0ab709c308a607e6063806d905830535055f045c03dc01dd005200d1002a02;
    decBuf[7474] = 256'h28048c06cc08420a1e0c490e551031126e125611bf0e900b9208a00646069806;
    decBuf[7475] = 256'he3069f06e605cd04ce0343036d032d04db043a05900576055e059f052906ed06;
    decBuf[7476] = 256'hd80777089308ad083708f607e207f407040831082308ce075507e4067c066f06;
    decBuf[7477] = 256'hac063b07eb07c10851096b09f408db078206e0045703f20167013d01fd01f102;
    decBuf[7478] = 256'h0e04670508072108ba08e80813093909a209000a1d0a030a5d09180877067e04;
    decBuf[7479] = 256'h2a03f5014d011a014801c7013a02e802c5038f0446058d05ce053006d106ea07;
    decBuf[7480] = 256'hf608300aaf0a880a4e097f07cf0546044703bc02e901c3015a01fb0018013201;
    decBuf[7481] = 256'ha90115029e02f802ab03b004ea0565076408ef08710817077605ed035403c902;
    decBuf[7482] = 256'hf3021903f60258025601a70009005f007f0125031e0572062b0783061e052003;
    decBuf[7483] = 256'h44018a00c300c201a902280301035302b50125010b01b10174025f03be031404;
    decBuf[7484] = 256'h2e041704aa0321035c023d01300082ff23ff06ffbdff9300cf01f602b6031f04;
    decBuf[7485] = 256'hff03a903f202ab023f020402aa01f800c3ff48fe7dfc48fba0fad3fa17fc3bfe;
    decBuf[7486] = 256'hdc000a040907fa080a0ab70942086606b5042c03c701e000b9ffacfee7fc36fb;
    decBuf[7487] = 256'h3df9e9f730f7d8f7a3f9cffb70fee9008502fa033e0401045803590215019600;
    decBuf[7488] = 256'h2300bbffdaffbdff6ffff8fe36fe7ffdd9fcc3fc4cfd58feb2ff9a001801a500;
    decBuf[7489] = 256'h6bfff0fdf1fc66fc90fc03fdb1fd10fef4fd71fd9bfcd2fb84fbcbfb8dfc44fd;
    decBuf[7490] = 256'h1afe70fe8afe14fe7cfdf3fcbdfcadfc9efc41fc8bfb6bfa5ff925f8a7f71af8;
    decBuf[7491] = 256'h0ef9a9fa32fc97fd22fea0fec7fe2fffcdffd0007f015f015c0051feb0fb37f9;
    decBuf[7492] = 256'hf7f617f65bf699f641f7daf7c2f840f94dfa41fb5efcd1fcf4fc95fccbfbe0fa;
    decBuf[7493] = 256'h42faecf9d2f949fa89fac4fad6faa5fa3efae1f9bcf9c7f90dfa84faf6fa5dfb;
    decBuf[7494] = 256'hbafb0ffc72fcb5fcc1fc74fcdefbc5fab9f97ff8acf739f7d0f6f0f60df727f7;
    decBuf[7495] = 256'h6ef731f884f926fb1ffd73fe2cfff4fe8ffdeefbf4f9a0f8e7f7aff7e2f710f8;
    decBuf[7496] = 256'h3bf8c7f719f7baf69df6ecf6c2f7c4f8b8f957fa73fac2fa09fb75fbfefb58fc;
    decBuf[7497] = 256'h27fc67fb48faa2f819f780f652f67cf6eff69df77ef727f7a5f62ef618f6a2f6;
    decBuf[7498] = 256'haef7a1f97dfbb1fccafd97fdaffc88fbe2f959f85af772f6f4f5cef565f585f5;
    decBuf[7499] = 256'ha1f524f6faf6fdf7abf849f966f94cf934f94af984f902fa53fa44faccf9d8f8;
    decBuf[7500] = 256'h9ef777f6b7f54ff56ef5fef5e9f606f812f9c1f95ffa7cfa62faebf9aaf96ff9;
    decBuf[7501] = 256'h81f9b2f936fad7fa43fb57fbdafae6f921f871f658f525f553f526f67ff767f8;
    decBuf[7502] = 256'h3af9faf91dfa3cfa1ffa3afa22fa0cfaf9f9e7f975f9d3f867f82cf885f858f9;
    decBuf[7503] = 256'h22fad8faf0fa84fafbf9a1f991f982f95af9d5f8ecf70ff77ff699f66ff772f8;
    decBuf[7504] = 256'hacf97efa3efb32fcd1fc60fdaffd67fd23fc82faf9f894f7acf62ef654f6bdf6;
    decBuf[7505] = 256'h1bf7abf762f867f916faf3fa83fbd1fb18fc59fc46fcc9fbd5fa9bf920f887f7;
    decBuf[7506] = 256'hfcf626f799f7bcf7dbf732f8b4f88af98dfa81fb1ffc3cfcb9fb13fb7cfaf2f9;
    decBuf[7507] = 256'hbdf9edf9fcf9eff982f9c2f8d7f7f9f66af684f689f74ef97afb85fdd9fe93ff;
    decBuf[7508] = 256'h3b00080036000c0099ff5ffe90fce9f96ff78bf460f306f358f338f48cf5c1f6;
    decBuf[7509] = 256'h4af8aff9f4fa6ffc6efd56fe28ff02ff99fe7dfd70fcc2fb63fb2cfcb4fd3dff;
    decBuf[7510] = 256'hd6ffa7ff80fedafc51fbb8fa44fb16fc89fc21fc04fb5ef945f846f775f747f8;
    decBuf[7511] = 256'h54f98efa60fbd4fbf6fb16fc33fc4dfc65fcd1fc81fd57fe93ffba00c7017502;
    decBuf[7512] = 256'hd402b702cc013100c8fde4fa2bf8b2f5bbf4dbf31ff4d8f461f62cf857faf8fc;
    decBuf[7513] = 256'hbdfefc00dd01a9026b02c301c400dcff09ff96fe2dfe0efef1fdd7fdbffd7efd;
    decBuf[7514] = 256'h1cfdc3fc30fccefb51fb20fb2ffb8dfb2afc18fdf6fd85fe08ff20ff35ff49ff;
    decBuf[7515] = 256'h5bff2affe0fe18fe15fddbfbb4fa8efa3cfb98fc96fe7200a701c0028d025e02;
    decBuf[7516] = 256'h8c01cc00630044009a00e8000001690042ffc7fd62fc7afba4fbb1fcebfd66ff;
    decBuf[7517] = 256'hffff2d00030090ff6dffccff95004c0122027802c7023d037e032f04a6041205;
    decBuf[7518] = 256'h250584046b03c5013c00d7fe93fd14fd3bfda3fd02fe92fe15ff8bfff7ffcf00;
    decBuf[7519] = 256'hd201c602a4036d04bb04d304bd04820471044004d90345039502ef01d9011402;
    decBuf[7520] = 256'hb502a3034104970414043f033c0202012f0009002c0009014502c103c0044b05;
    decBuf[7521] = 256'h210514044f022300adfe69fe9eff9701fb03df0698095c0bae0bce0a7a09ca07;
    decBuf[7522] = 256'hd105f50345022c01c7ffdffe61fe3afe5dfefbfe3800b3017e032e05b7061c08;
    decBuf[7523] = 256'hbd09d60a6f0be40a690938072c05600423043b050607b608cf09020a7709fc07;
    decBuf[7524] = 256'h31060504fa01a6006800100175027404c805fc06a5073e086c08ea08aa09130a;
    decBuf[7525] = 256'h330adc09f108950751062a05b7041f05fd05ac075c09550b210c5f0cb70bb80a;
    decBuf[7526] = 256'h73094c08f306ae053304ce0243026d027a038505bb08ba0bab0d700fc20fe20e;
    decBuf[7527] = 256'h160e650cdc0aab08a0064c0593045b045a05fb0684088309b1093309da079506;
    decBuf[7528] = 256'h6e05ae04d104ee0547078c08070a060bee0bc00c800d2f0ed00d070db30b120a;
    decBuf[7529] = 256'hf908600832085c08820819083c077306f00508062107c708500ab50b400cc20b;
    decBuf[7530] = 256'hb50a3609d107e906bf06e50693073108c10844098b09a109030a5c0a6c0a990a;
    decBuf[7531] = 256'h8b0a970afa0a8e0b650cf50c0f0dc80cda0b7e0add08c4075f06d40556052f05;
    decBuf[7532] = 256'h5205f005f3062d085409ad0a950b680cdb0c440da20dbf0dd90df10db00dd80c;
    decBuf[7533] = 256'h630b9809f0062c0535048004d40500087509c90a070bcf0a9c0a270ba50bb20c;
    decBuf[7534] = 256'h600d020dc50ba2099607ba058604dd031004f804cb05d706cc07e808f509740b;
    decBuf[7535] = 256'hd90c1e0ef10e640ffb0edf0d850ce40aeb08970762064905b004c8034a037003;
    decBuf[7536] = 256'h93033104fb04e605c306c607ba089709610ae30a2b0b150b010ba80a360a9409;
    decBuf[7537] = 256'ha6084a0706063604010359022602b102d8033105d306eb07ea081909ef08c808;
    decBuf[7538] = 256'h600840085d0877085f081e089507f4065d06220610060006d305400568049f03;
    decBuf[7539] = 256'he802d10268038e04b505c206700790073a078306dc051a05cb0484049a04fc04;
    decBuf[7540] = 256'h9d055f06e2065907430793068d05530481035a03090425057f060a07e006d305;
    decBuf[7541] = 256'h99047203b3024a02a902390387039f0389032703f10202032e037103ad03a203;
    decBuf[7542] = 256'h5c030a03e9021b0392034504bb04fc04e9048f041d04b60373031e03d1024f02;
    decBuf[7543] = 256'h8b01a000c2ff33ff18ff8fff7d009a015a02c2022402ae00e3fe33fd8bfcbefc;
    decBuf[7544] = 256'h49fdc4fe29006e019402a1030a0429044604f803b003ee02ce0128009ffed4fc;
    decBuf[7545] = 256'h24fb7cfa49fa31fbacfcabfdeffe1afff3fe45fee6fd90fdaafdf1fd5dfebffe;
    decBuf[7546] = 256'hf5fe05ff14ffecfee0fea9fe77fe12fe9afd08fd57fcb1fb9bfbfdfbe6fc42fe;
    decBuf[7547] = 256'h86ff050091ff58fe34fc29fad5f81bf8e3f77cf864f937faf7faa5fb04fc5afc;
    decBuf[7548] = 256'ha9fc1ffde2fd99fe3fff55fff3fee6fd40fcb7fa52f96bf840f867f88af8e9f8;
    decBuf[7549] = 256'h3ff959f971f95bf9f9f834f849f76cf616f664f6c8f793f9bffb35fd79fd3bfd;
    decBuf[7550] = 256'h22fc57fa23f90af871f79ff71ef891f8f9f8daf811f8bdf61cf503f404f3d6f2;
    decBuf[7551] = 256'habf21ff387f325f428f5a8f673f8a7f9c0faf3fa68fa95f93cf8f7f625f6b2f5;
    decBuf[7552] = 256'h8ff530f513f5c5f41ef45cf3a5f2fff1bef1f9f1e1f2bef3c1f470f58ff5acf5;
    decBuf[7553] = 256'h92f57af539f5d7f412f45cf3e5f279f265f2e2f274f325f4cbf40cf56ef5a4f5;
    decBuf[7554] = 256'hd5f5c6f5b9f533f592f4d0f3e5f207f277f1f5f07ef012f0feef34f0c6f077f1;
    decBuf[7555] = 256'hacf2d2f32cf570f697f7a4f8c7f8e9f73af60ef46ef1a9ef57ef0cefd8ef91f0;
    decBuf[7556] = 256'h3af16df13ef169f18ff13df29cf2b9f29ff2b7f2f7f281f345f4fcf414f5fef4;
    decBuf[7557] = 256'h4ef4d7f396f383f3b8f309f4ddf365f3b2f27df156f04aef9beebbeef7efc7f1;
    decBuf[7558] = 256'hf2f368f534f6f6f5def479f334f262f13bf118f138f1a8f026f0afef6eefa9ef;
    decBuf[7559] = 256'h4af038f193f2d8f3fff40cf600f75ff742f728f781f6eaf539f564f461f36df2;
    decBuf[7560] = 256'h50f1f7ef0fefe8ed28ed4bed28eed8ef03f279f355f50ef6d6f509f638f662f6;
    decBuf[7561] = 256'hd5f6f8f699f696f517f418f38cf20bf317f451f524f64af6e2f544f5b4f49af4;
    decBuf[7562] = 256'hb1f4c7f4b3f45af4c8f317f3d0f2baf21cf3e1f3ccf4aaf539f6f0f637f7a4f7;
    decBuf[7563] = 256'hb7f711f862f8acf8d4f8f8f8c1f87bf829f8f2f7e8f7dff7b6f754f7c1f610f6;
    decBuf[7564] = 256'h9af559f56cf57ef58ef59df5c5f563f651f76df8c7f9affad9fab2fa04fa66f9;
    decBuf[7565] = 256'h49f998f90efa7afa8efa7cfa4bfa1ffa12fa1efa29fa33faf3f977f98ff8b2f7;
    decBuf[7566] = 256'h22f73cf712f8c1f9edfbf8fdc4fe86fedefd79fcd7fabff926f954f9d3f992fa;
    decBuf[7567] = 256'h87fba3fc63fdccfdacfd1cfdfdfbf0fafcf99df9f4f9aafa0ffc74fdb8fe37ff;
    decBuf[7568] = 256'h5dff3aff1bfffefe18ff5fff4affc0fefcfddcfc1cfcb4fbd3fb63fc4efd6bfe;
    decBuf[7569] = 256'h77ff6c008801950243036303d3027f01deff55fef0fc65fc8ffc4ffdfdfd5cfe;
    decBuf[7570] = 256'hb3fecdfe14ffabffaa00e4015f03c404ac057f06a506c8066906da052305ee03;
    decBuf[7571] = 256'hc702210198ff33fe4bfd21fd94fd88fe2300ac017703ac0454058705b6058c05;
    decBuf[7572] = 256'hb2056006ff068e07dd07f407b4077907d806400641050704e102d40126010601;
    decBuf[7573] = 256'h96014d0252038c045e056b065f07fd07c608490990097b0940097b085c070206;
    decBuf[7574] = 256'hbe04eb037803e103fd04f006cc08f80a6e0c3a0dfc0c540cef0aaa0983087607;
    decBuf[7575] = 256'h0e07af06cc06e606fe06e8065f0676055a049a037703d6034b057c071d0a970c;
    decBuf[7576] = 256'hd60ee21036126a1332133312ef10cb0ec00c6c0bb30a0a0a71092d0809066803;
    decBuf[7577] = 256'ha4010800beff9a0141042408c40b0f0f321124137e13d013f01224126b11c210;
    decBuf[7578] = 256'hc30fdc0eb50d0f0c860a210939080f083508e3084209d209550a2a0bf40b130d;
    decBuf[7579] = 256'hd30d3c0e5b0e780e920e090f4a0f850f2b0f780e730d7f0ca20b4b0b9a0b400c;
    decBuf[7580] = 256'h590db30ef70f1e119111b411551119109e0e390d970b7f0ae609b7098d09000a;
    decBuf[7581] = 256'haf0a4d0b160ccd0c730ddf0d690e0a0f23107c11c112931307145813bd11c40f;
    decBuf[7582] = 256'he80dbc0b460a7a093d09e509180a000b7e0bf10b140cb20c7c0d9b0ea80f5610;
    decBuf[7583] = 256'h76101f109d0f560f150f280f160f470f380ff60eb90e560ec30dc40c8a0b0f0a;
    decBuf[7584] = 256'h10098508af086f09630afe0b870d520f86109f11d2114711c910bc0f0e0f6f0e;
    decBuf[7585] = 256'he00df50c990b540a2d0907096f098c0ae50b2a0d540d7b0d120df20c0f0d5d0d;
    decBuf[7586] = 256'h750d600dd60c590cc70b8c0b7a0b6a0b3e0bc50a530acf099909ca094f0aef0a;
    decBuf[7587] = 256'hdd0bbb0cbd0d6c0ecb0eae0ef70d930cc80a1809ff076607940713088608ee08;
    decBuf[7588] = 256'h0e09b808d208ba082609b009740a2b0b010c570c710cfb0be10a8809e707ce06;
    decBuf[7589] = 256'h350663063607f607ea088809a50922091d08e306bc0549056c050a0646076d08;
    decBuf[7590] = 256'h2d0996093709e1085e081708d607c2076907180793061606e505d605e4050806;
    decBuf[7591] = 256'h1306cd057b05ec048a047804c9046b052e06e506cd068c068d059904fb03de03;
    decBuf[7592] = 256'h2d04d3046a05a505930562051905f104e404ad0453049e03e702110281019b01;
    decBuf[7593] = 256'he3014f02ff027603e20344047a048a047b0439049b03d8022102ab016a017d01;
    decBuf[7594] = 256'hd7014902b002a2027e021b02d801b401d501df01b10135012900d0fe8bfdb9fc;
    decBuf[7595] = 256'h46fcf4fc11fe6affaf00d50149026b024c02f601a70160011f01e400af003d00;
    decBuf[7596] = 256'hb8fff3fe3dfe67fd9efc1bfc03fc19fc54fc89fc79fc6afc78fccdfc5cfd0cfe;
    decBuf[7597] = 256'h83fe6dfe0bfe47fd90fc48fc5efce7fc65fdd6fd03fedafd9efd25fd93fce2fb;
    decBuf[7598] = 256'h3cfbd0fa95fa83fab4faa5fa97fa5bfa24faf2f9c4f9abf995f973f979f9b7f9;
    decBuf[7599] = 256'h11fa97faf0fa21fb12fb05fbe0fad5fadffad6fa8cfa1efa5ef9a7f831f846f8;
    decBuf[7600] = 256'h81f8fef82ff903f970f898f708f7eef635f7cdf77df8c4f8aff84df8d0f75ef7;
    decBuf[7601] = 256'h4ff792f7e7f71ef828f81ff816f8f1f7cff771f7a8f6a5f56cf445f3d2f23af3;
    decBuf[7602] = 256'h57f4fdf586f785f810f992f8d2f723f785f668f6b7f62ef718f7ddf63cf67af5;
    decBuf[7603] = 256'hf7f4dff49ef463f4e6f3f3f273f174f0e9ef67f027f11bf2b9f210f35ef3a5f3;
    decBuf[7604] = 256'h68f4bbf55df7e6f87ff9f4f8cdf7daf586f451f319f3b2f3e0f35ff4ecf3b2f2;
    decBuf[7605] = 256'h37f1d2ef46ef1cefdcefd0f0aef104f2eaf144f1d7f0ebf021f1b3f164f2daf2;
    decBuf[7606] = 256'h46f3d0f329f49bf4c7f4d5f4b0f48ff449f41cf4d1f363f3c1f2d3f1f6f0f3ef;
    decBuf[7607] = 256'h8aef6befc1ef78f04ef117f265f24ef2b6f12df18cf076f0b1f0e7f038f147f1;
    decBuf[7608] = 256'h1ff1faf047f1ddf122f366f4e5f40bf517f4faf23af2d2f131f2faf2b1f399f3;
    decBuf[7609] = 256'h02f3dbf1b4f0a8ef85efa5ef34f0b7f02ef16ff182f1b8f1e9f132f25af27ff2;
    decBuf[7610] = 256'h8af26cf263f25af244f22ff229f23af27df2f3f265f3ccf30ff4ebf3b4f382f3;
    decBuf[7611] = 256'h66f36ff376f354f3f6f263f2b2f10cf1cbf0dff014f1a7f130f2f5f277f3eef3;
    decBuf[7612] = 256'h2ff46af47cf46bf45df4fff392f3d2f2e7f149f1f3f00df1b3f1a1f27ef381f4;
    decBuf[7613] = 256'heaf448f59ff521f669f6d5f637f725f7f4f66ff6f2f581f537f50ff5d2f46ff4;
    decBuf[7614] = 256'hc1f31bf358f20af222f2b9f26af310f47cf490f4a2f4d2f457f563f6bdf701f9;
    decBuf[7615] = 256'h28fa9bfa33fa94f9cbf8acf7ecf63ef69ff583f59df5b5f521f6aaf64bf739f8;
    decBuf[7616] = 256'h55f915fac4fae3fa54fa9df997f8a3f705f7aff661f619f6d8f576f541f5b2f5;
    decBuf[7617] = 256'h90f6ecf78df916fb7bfc06fd30fd0afd5bfcbdfb2dfb13fb5bfbf2fb7bfcf8fc;
    decBuf[7618] = 256'h09fda1fcd9fb9dfa21f922f897f7c1f735f8e3f881f911fa5ffad6fa6dfb1efc;
    decBuf[7619] = 256'hc4fc5cfdbefd17fe48fe92febafec6fe8ffe21fe7ffd12fdfffc11fd82fdeafd;
    decBuf[7620] = 256'h62feb3fefdfe40ff7dff88ff2eff78fe58fd4cfc9dfb3efb95fb4cfc21fd5efe;
    decBuf[7621] = 256'h84ff4400f3009101ae015f011801ac0071005f00d10091014702ee022f031b03;
    decBuf[7622] = 256'hc2020f020a015b00bdff67ff81ff27001501b30143025d02e6017a013f012d01;
    decBuf[7623] = 256'h7f012102e4029a037004c60415052d051705b504a3049304bf043705a9051006;
    decBuf[7624] = 256'h03069605b9049c038f029b013c01930149024f03fd03da0431057f05f6058d06;
    decBuf[7625] = 256'h3e071408a30826093e0928091409df086d08cb0708071d064005760428044004;
    decBuf[7626] = 256'h8104e304600513068906ca06de0685063306070665061b07a2080c0ba70c870d;
    decBuf[7627] = 256'hcb0d120df90bfa0a130a400980088c07ee062506d605be05d4050f0621065206;
    decBuf[7628] = 256'h9b062e07df07b508b809660a430bd30b210c390c240c100cfe0b0e0c580c9b0c;
    decBuf[7629] = 256'ha70c440c7b0bb20ac709ea08930879083208f107b6078107b107540842099d0a;
    decBuf[7630] = 256'he20b600cd40cf60c980c410c270c0f0c250c110cdc0bab0b9c0b8f0bb30b000c;
    decBuf[7631] = 256'h460c860c7e0c490ce20b400b7d0a9209f40864087f08f508b8096f0a450b9b0b;
    decBuf[7632] = 256'h1d0c650ca60c2f0dac0d1e0ea30efc0e0c0fe00e820efd0da40d320dad0c300c;
    decBuf[7633] = 256'h5d0b200aa5084007fc057d05f005e5068008790acd0b020daa0ddd0d680e3e0e;
    decBuf[7634] = 256'h640ecd0eed0ed00eb60e0f0e4d0d960cf00b580b1d0be80a760af10974090209;
    decBuf[7635] = 256'hf40837098b09ee09fc09d709b609c009250ad30aa80b380cbb0ca30c8d0c530c;
    decBuf[7636] = 256'h1d0cec0bc00bb30b8e0b990bb70b090c400c4a0ce60b380b620a6009b108d407;
    decBuf[7637] = 256'h4407f606de064a07d307bc0899099c0a4a0ba90bff0b4e0c950cd60cc20c690c;
    decBuf[7638] = 256'hd70bff0a360a7f09a908e0075d07160700076207df075108b808c608d2081f09;
    decBuf[7639] = 256'h7909fe099f0ae00acc0a730a010a7d0947091609cc083908610798064a066206;
    decBuf[7640] = 256'hf906d1079a08b4086d08aa07f3067d0692061c070408e10871095709e008f207;
    decBuf[7641] = 256'h150785063706ae061a0755076707f5065306bb0580059205e3052d0655064906;
    decBuf[7642] = 256'h28060a06ef05e705c1059f057f056f059205c50503061c062306010607062f06;
    decBuf[7643] = 256'h67068d065c06ff053605c003c10236020c0232029b02780308048b04a3048d04;
    decBuf[7644] = 256'h2b04d103c1030b048304f5042105f9048c0442043504590490048604fd03d702;
    decBuf[7645] = 256'hb0015700ccffa2ff15000901e601af0266030d044d043a04040492034903eb02;
    decBuf[7646] = 256'hae02770209028501e400a3008f00c5005701b90113020202b9015b010601cf00;
    decBuf[7647] = 256'h89003700eaff90ff6cff77ffbdff3300a500ef001701f300d2008c003900d6ff;
    decBuf[7648] = 256'h94ff6fff90ffeaff70001001510165012f019d001400baff69ff3dff15ffc0fe;
    decBuf[7649] = 256'h47feb5fd04fd8dfc4cfc39fc6efcc0fc27fdd5fdaafe74ff5f00fd0053016d01;
    decBuf[7650] = 256'hf70009002bff29fe34fdd6fc7ffc31fc19fcd8fbc5fbd7fb07fc8cfc09fd7bfd;
    decBuf[7651] = 256'ha7fd9afd75fd3efd48fd76fdd1fd26fe47fe3dfe21fed7fda5fd65fd1bfdadfc;
    decBuf[7652] = 256'h0bfc48fb91fa1afa05fa18fab9fa7cfb33fcd9fc45fd59fd47fdd5fc8bfc63fc;
    decBuf[7653] = 256'h3ffc4afc68fc5ffc46fc12fcb8fb63fb16fbd0faa3fa9afac0fa0cfb66fba2fb;
    decBuf[7654] = 256'hc3fba5fb53fb1cfbfefa2cfb76fbbcfbd7fbbffb8afb3efb0cfb03fbfbfad6fa;
    decBuf[7655] = 256'hb3fa6efa2ffa16fafff9f8f90bfa06fa1ffa5bfab6fa23fba8fbdefbcdfb66fb;
    decBuf[7656] = 256'hb8fa12fa7bf940f952f982f907fa84fa37fbaefbeffb02fca9fb17fb3ffa75f9;
    decBuf[7657] = 256'h8af8ecf75cf742f75af7c6f750f8f0f888f911fa8efae0fa29fb51fb5efb53fb;
    decBuf[7658] = 256'h21fbcefa81fa4ffa10fae6f9d0f992f948f9eef899f84cf81af8ecf7d3f7bdf7;
    decBuf[7659] = 256'hb6f7d5f72af8aff850f913fa95fadcfaf2fab7fa3afaa8f9f7f880f840f853f8;
    decBuf[7660] = 256'h65f8b6f800f90df91af90ff919f946f980f9b4f9d7f9b8f963f9def861f8eff7;
    decBuf[7661] = 256'hc3f7b5f7c1f7ccf7c2f7b9f7d2f707f86ef810f9a7f931fa8afabbfaacfa69fa;
    decBuf[7662] = 256'hfcf977f9faf888f83ff8fcf7bff75cf719f7ddf6d2f618f78ef721f8aaf8e0f8;
    decBuf[7663] = 256'hf0f8e1f8b9f8c5f812f96cf9d9f940fa69fa2cfab3f9bff8cbf7eef697f67df6;
    decBuf[7664] = 256'hc5f65cf7e5f73ff84ff840f84ef872f8a9f803f940f935f92bf9ebf8a0f882f8;
    decBuf[7665] = 256'h67f83ef827f813f819f84cf8a5f82af9a7f9d8f9acf969f9e4f867f815f8aef7;
    decBuf[7666] = 256'h86f749f7fcf6a2f67ef65df67bf6cdf630f7a8f73bf8c4f81df9b0f912fa6bfa;
    decBuf[7667] = 256'hfdfa38fb6efb1dfb7afa8df9aff8e6f798f750f73bf700f7a6f655f646f6a4f6;
    decBuf[7668] = 256'h42f730f8cef824f93ef926f911f94cf9c9f95bfae4fa3efb0dfb88fac4f9d8f8;
    decBuf[7669] = 256'hfbf732f7aff668f67ef6b8f659f747f825f9b4f937fa4ffa0efad3f97af969f9;
    decBuf[7670] = 256'hb3f92bfabefa20fb32fbc0fa3bfa77f9c0f878f838f824f836f846f855f898f8;
    decBuf[7671] = 256'h05f98af907fa58fa84fa92fa85fa90faaefaa5fa7cfa1bfa87f925f9ccf8dcf8;
    decBuf[7672] = 256'h26f99ef910fa5afa9dfad9fafafa2cfb35fb2dfb26fb1ffb19fb1efb05fbbffa;
    decBuf[7673] = 256'h65fae0f986f956f947f954f960f955f94bf979f9b3f923fad6fa4dfbe4fb95fc;
    decBuf[7674] = 256'h0cfd78fddafd0ffefffdb5fd22fd72fccbfbdefa3ffab0f92df915f92bf966f9;
    decBuf[7675] = 256'h07fa9efa76fb79fc27fd04fe21fe07fe90fdf9fc70fcf2fbc2fb95fb6dfb31fb;
    decBuf[7676] = 256'hfafadcfa09fb85fb4afc35fdd3fd63fe7dfec4feaefec2fed4fee4fe9afe3dfe;
    decBuf[7677] = 256'hd0fd4bfdf2fca0fc74fc4cfcf7fbaafb64fb36fb60fbd0fba3fca6fd9afe78ff;
    decBuf[7678] = 256'h07008a00a20061002600f0ff9fff55ff13ffd6fe89fe43fedffd81fd2cfd21fd;
    decBuf[7679] = 256'h3ffd7ffdeafd51feaffe04ff51ffbfff4400e5007c01b701a501130114001fff;
    decBuf[7680] = 256'h03fe90fd6dfdccfd95fe4cfff2ff5e009900f2004401e6017d02df02ce027c02;
    decBuf[7681] = 256'hda01ec004e00beff70ff29ff13fffffeeefeddfe0aff9dff4d00530147022403;
    decBuf[7682] = 256'hb40336044e040d04d2039d030b0381029901bb00b9ff50fff1fe0eff91ff0700;
    decBuf[7683] = 256'h7300fd00c10178027e032c04ca045a0574058c05760562052d05dc0439047703;
    decBuf[7684] = 256'hc0021a02ad0173013d010c01e000ed0012018b013d021303dc0393040a057605;
    decBuf[7685] = 256'hb1050a063b064a063d06e8055905a804d203090386026f02db028b0361042a05;
    decBuf[7686] = 256'had05f4050a06f605e405b40587055f052305c0044704d6036e0346036b03b803;
    decBuf[7687] = 256'h4e04e50496056b06fb06b207f9073a084e081808c7077d07050793062c06ce05;
    decBuf[7688] = 256'h790558052605f904ae04680428041004260480040505ca05800686077a081809;
    decBuf[7689] = 256'ha809f609af094309b908f5077207cc066006fe05c805b80501067a06ec067007;
    decBuf[7690] = 256'h820772076307560762079907df071f0869089b0880084608d5074307ba066006;
    decBuf[7691] = 256'h7106d8066b07f4077208a208ec084a099f09ec091e0a140aba097d0946091409;
    decBuf[7692] = 256'hd4085808700753069405e5040505ce05ed0647088b095e0ad10af40a140bbd0a;
    decBuf[7693] = 256'h6f0af8098c0951093f092f090309c00883083608dc07d007f1070f086108ae08;
    decBuf[7694] = 256'hf4085909b609f309140af60992093409c708600838082b084c08a60814097b09;
    decBuf[7695] = 256'hd809e509ae095409ff08de08fc084e099b09b909b009760932090509fd080409;
    decBuf[7696] = 256'h0b09ec08c4088c086608600872089a08dc081c0945097a099c09a309a809ad09;
    decBuf[7697] = 256'hb209d009db09ca099b093409af083208c0077607690775076a0774079007c907;
    decBuf[7698] = 256'h3a08ed086309cf090a0ad50983091c09bf08820877086d089b08e5082b095809;
    decBuf[7699] = 256'h5009ef085c08ab07050799068506de065007b70715086a088b08810865081b08;
    decBuf[7700] = 256'had0746071e07120749077b07bb07d307ea07f107030814080508d20779072407;
    decBuf[7701] = 256'hed06e306fe0627073e072907f106ae066e0665065e0665067806720677067206;
    decBuf[7702] = 256'h660643061006d20588056a05610569058e05bf0503066806c5061a0751073307;
    decBuf[7703] = 256'he1065206c9056f053f056b0578059d057c053605bf044d04e603a3037f037403;
    decBuf[7704] = 256'h7e03be0308044e048e04a604900452041804110441048604fc046e05b805e005;
    decBuf[7705] = 256'hd405870519057704b403fd02860245023202200210020102d901cd01d801f601;
    decBuf[7706] = 256'h11025b02b5023b03dc037304d504c304310459039002d9019201510164015301;
    decBuf[7707] = 256'h4201340126013201530171019f01c801df01f3011302230233021c02e4018301;
    decBuf[7708] = 256'h0b017800160099ff68ff5aff9cff2200c3005a01bc01ce019d0119019b002a00;
    decBuf[7709] = 256'hc2ff80ff73ff68ff72ff8eff96ff9eff7bff36ffe4fe97fe79fe95fedffe61ff;
    decBuf[7710] = 256'hdeff50009a00c2009d005000ceff2dff96fe0dfed7fdc7fdf3fd1bfe27fe06fe;
    decBuf[7711] = 256'hacfd27fdaafc59fc0ffc01fc56fcfbfc01fef5fed2ff280042009cffdafeeefd;
    decBuf[7712] = 256'h50fdc1fc72fc5afc70fc84fcb9fceafcf9fcebfcaffc62fc08fccbfb94fb9efb;
    decBuf[7713] = 256'hbafbe3fbeafbe3fbc4fbbffbb9fbd1fbfffb38fc6cfcaafcd3fceafcf1fcd1fc;
    decBuf[7714] = 256'h9ffc61fc06fc99fb32fb9ffa15fa98f967f976f9b9f9f6f92dfa23fad0f983f9;
    decBuf[7715] = 256'h51f97ff9fbf9bffa76fb1dfcb4fcc8fcb6fc64fcc2fb00fb49fa73f9e3f895f8;
    decBuf[7716] = 256'h4ef838f824f836f826f852f860f89cf8d3f819f96bf9cef92cfa69fa8afa6cfa;
    decBuf[7717] = 256'h19fab6f959f934f913f909f9eef8e6f8b1f881f849f805f8c6f77bf735f7f5f6;
    decBuf[7718] = 256'hedf613f76cf7f1f76ff8c0f80af9e1f8bdf886f840f800f8e7f7c2f7adf7c0f7;
    decBuf[7719] = 256'hc6f7eaf713f824f81ff811f8daf796f756f7fcf6bff688f656f65ff678f69df6;
    decBuf[7720] = 256'hb2f6d1f6ccf6dbf60ef75af7b4f721f82ff822f8e5f782f725f7e8f6b1f693f6;
    decBuf[7721] = 256'h78f63ef6fbf5dff5c6f5ecf545f6b2f637f7b4f7c5f7d3f790f70bf78ef63df6;
    decBuf[7722] = 256'hf3f5e6f50af641f687f6c7f6cff6c8f6a5f654f607f6d5f5baf5d2f525f69ef6;
    decBuf[7723] = 256'h10f777f79ff793f788f742f714f7fbf6d6f6c1f6c8f6b7f6bcf6caf69bf64af6;
    decBuf[7724] = 256'hd1f53ef5dcf4a7f4d7f47af53cf6f3f699f706f819f82bf81bf8d1f7a9f785f7;
    decBuf[7725] = 256'h7af784f79ff786f761f731f7d3f690f653f61cf6d6f5a9f590f5a6f50ef6b0f6;
    decBuf[7726] = 256'h72f729f8a0f8b6f8c9f894f842f816f8d3f797f74af718f7fcf605f71bf730f7;
    decBuf[7727] = 256'h5bf761f785f7c1f70bf879f8e1f823f948f953f921f9e1f8b8f874f834f8fbf7;
    decBuf[7728] = 256'ha8f75bf729f7fbf604f747f799f712f884f8cef8f6f81af951f997f9fcf974fa;
    decBuf[7729] = 256'hc5faf2fae4faa8fa45fae7f97af930f9edf898f861f807f8b2f77bf75df78bf7;
    decBuf[7730] = 256'h07f8a8f896f9b2fa72fb20fcbffcdbfc8dfc46fcdafb50fbd3fa41fab7f95ef9;
    decBuf[7731] = 256'h0df9e1f8eef812f975f9eef95ffac7fa24fb61fb82fb8cfba7fbd1fb23fc70fc;
    decBuf[7732] = 256'hb6fce4fcbafc59fce1fb4efbecfab7fac7fad6fa18fb55fba2fbe8fb4cfcaafc;
    decBuf[7733] = 256'hfffc4cfd56fd3bfd01fdbdfc7dfc65fc5dfc72fc78fc89fc8efc93fc9ffccafc;
    decBuf[7734] = 256'h08fd52fdacfde9fd0afe14fe0bfee1fdcbfdc4fdd7fdf3fd17fe2efe32fe17fe;
    decBuf[7735] = 256'hf8fdd1fdadfd84fd68fd4efd53fd8afdfafd8dfe3dff85ff9aff87ff2dffdcfe;
    decBuf[7736] = 256'hb0fea2fedffe2cff72ffb2ffdbff010007000100cfff83ff3dffebfecafee8fe;
    decBuf[7737] = 256'h3aff9dff30009200a40094004a00d2ff80ff72ff9affefff3c006e0077007f00;
    decBuf[7738] = 256'h78008c00b800f60040017201a001c901fd0120023f0239020b02ae011a019100;
    decBuf[7739] = 256'h380007003300ac003e01c701fd012e023c0214020802130245028502cf020103;
    decBuf[7740] = 256'h1d031403fe02ce02950261023f022c02260240027302b102ea02100332034503;
    decBuf[7741] = 256'h61038503ca0310043e0446041204c603940366036f039403b703bd03b7039e03;
    decBuf[7742] = 256'h90039c03bf03f20330045904700477047d048304a604d904fc04270538052905;
    decBuf[7743] = 256'h1b050605fa040c0534055c058a059d05800552050e05ce04a404bb04d0040805;
    decBuf[7744] = 256'h3c05510570059805bb05f805310648065c06630668068206ac06bc06cc06be06;
    decBuf[7745] = 256'h8f06570631060106d605b905aa05c10501066506de064f077c07890765072e07;
    decBuf[7746] = 256'h1007f406dc06d406bf06b906ca06ee0621075f078807ad07c207e107dc07d707;
    decBuf[7747] = 256'hb6077f074a07280722073e07620779079707b207c307ec0713082d0844084808;
    decBuf[7748] = 256'h3d0840084a084708490839081908ef07de07d907f0070e082908500869086e08;
    decBuf[7749] = 256'h6a084f081a08f507d207d80722086808ba08f108fb08cd08a4088d086b087108;
    decBuf[7750] = 256'h82087d08a708d90817097209960975092f09b9082608eb07b607a607d207c407;
    decBuf[7751] = 256'hb807d9070b083908a408ee08160922092d09370953096b0973097a0967091e09;
    decBuf[7752] = 256'hd8087308fb07aa0760076d07aa0723089508df082109fd08c608940854083b08;
    decBuf[7753] = 256'h34081f08260836085a088d08cb08e408eb08c9089d08760852083b082e081b08;
    decBuf[7754] = 256'h0908fa07eb07d407ca07c207b407c507e50705083d08710886088c0870083708;
    decBuf[7755] = 256'h0308b7075d0721070007f60623074d079007d0070a0820083508480864087d08;
    decBuf[7756] = 256'h82085308f5077d07eb0661062c06fb050a0617063c067306b9060b0758077607;
    decBuf[7757] = 256'h7f07770760074b076b079207b607cd07b8077e0723079e062006af0547050505;
    decBuf[7758] = 256'h11054805a205f7055a068206be06c906d306dc06d406a00670062b06eb05b105;
    decBuf[7759] = 256'h8c054e051405d104a304ab04d1042a059705e105090615060a06ec05d105a805;
    decBuf[7760] = 256'h64051205c50493048a049204a904bd04b704900461044204260421040a04ec03;
    decBuf[7761] = 256'hd903d503e503100448047d049104a4049e048f046f042f04ef0394033f031e03;
    decBuf[7762] = 256'h14031e0326031e03fc02d0029e027b028e02aa02d8021003450367036e035103;
    decBuf[7763] = 256'h0503a2024402ef01e401ee01090222022a0231022a0225021502fe01cf018b01;
    decBuf[7764] = 256'h4b012201290159019101b701be019f0161011601d000a300690053004c006b00;
    decBuf[7765] = 256'h9e00db0005011b011401f500e400d500c700a1005400dbff49ffbffe66fe56fe;
    decBuf[7766] = 256'h82fec5fe01ff22ff40ff5cff74ffa9ffd9ff050016000600efffc9ff9bff56ff;
    decBuf[7767] = 256'h16ffbbfe7ffe32fe00fed2fd98fd64fd42fd22fd28fd42fd62fd77fd73fd69fd;
    decBuf[7768] = 256'h5ffd6efd90fdbafde1fdf0fdf5fdf1fdd6fdb6fd90fd57fd14fdd4fc8afc58fc;
    decBuf[7769] = 256'h3cfc24fc0dfcf9fbf2fbf8fb1cfc45fc6dfc7cfc6efc51fc2efcfbfbcbfb9ffb;
    decBuf[7770] = 256'h61fb27fb02fbedfae7faf8fafdfaf8faf4fae8faecfa1bfb4bfb90fbbdfbd6fb;
    decBuf[7771] = 256'hdefbd7fbb7fb90fb4dfbe9fa71fafff998f93af92ef90df9dbf8c0f8b7f8cef8;
    decBuf[7772] = 256'h27f9adf94dfae5fa6efba4fbd5fba8fb80fb13fb71faaef9f7f851f8e5f7d1f7;
    decBuf[7773] = 256'hbff7d0f7def707f85bf8a8f802f957f98ef9acf9b5f9cef9d6f9f8f917fa1dfa;
    decBuf[7774] = 256'h03fadaf991f937f9e2f869f8d6f774f71bf7eaf6dbf604f728f75ff791f7d1f7;
    decBuf[7775] = 256'h3cf8a3f801f956f961f96bf974f96cf964f96bf93ff9ebf87ef8f9f7a0f72ef7;
    decBuf[7776] = 256'h02f7bff6b3f6a8f6c6f62af7a2f735f8bef8f4f8e3f8b7f874f838f817f8f9f7;
    decBuf[7777] = 256'hddf7e6f7cff7baf79bf769f72bf701f7ebf600f738f78af7d7f731f86ef8a5f8;
    decBuf[7778] = 256'hebf819f931f91bf9cff839f8a2f740f7e6f6f7f605f72df76af775f793f7aef7;
    decBuf[7779] = 256'hb7f7bef7c5f7bff7c4f7def7ecf701f81cf819f80ff807f8f4f7f2f701f807f8;
    decBuf[7780] = 256'h1af837f85af884f8c1f8ebf8f2f8def899f859f80ff8ddf7c1f7caf7c2f7c9f7;
    decBuf[7781] = 256'hdcf7d6f7dbf7e9f7e5f7e9f7faf710f83bf873f8b7f8e5f80ef915f901f9faf8;
    decBuf[7782] = 256'hf5f80ef926f93bf93ff93bf919f9f8f8dbf8b8f897f87af84ff83ef839f850f8;
    decBuf[7783] = 256'h7ff8c4f804f94ef994f9aff9c8f9c0f990f965f948f939f947f965f969f96cf9;
    decBuf[7784] = 256'h63f94ff951f970f996f9baf9d1f9d6f9d2f9dcf9ecf90bfa3afa4dfa5efa59fa;
    decBuf[7785] = 256'h4bfa36fa2afa18fa0ffa01faeef9e2f9dcf9d2f9dbf9f0f915fa58faaafa0dfb;
    decBuf[7786] = 256'h6bfba7fbb2fba8fb9ffb76fb50fb20fbe8faa5fa65fa2bfa14fa29fa48fa86fa;
    decBuf[7787] = 256'hd0fa2afb67fbb4fbe6fb01fc2bfc32fc55fc80fca8fcd6fce9fcd8fc9ffc5cfc;
    decBuf[7788] = 256'hf7fbb5fb78fb6dfb63fb6cfb74fb7cfb83fb89fb8ffbb2fbdcfb30fc85fcfefc;
    decBuf[7789] = 256'h70fdd7fd1afe6ffe90fe9afe91fe57fe14fec2fd75fd2ffd01fdf9fc00fd07fd;
    decBuf[7790] = 256'h0dfdfcfce3fcc2fcadfca2fcbafce9fc50fdd5fd52fea3fe0aff33ff26ff1bff;
    decBuf[7791] = 256'h11ff1bff33ff59ff7bff81ff7cff58ff2efff0fec7feb1feaafeb0fec1fee5fe;
    decBuf[7792] = 256'h0eff36ff4fff5dff59ff36ff0dffdafec5feccfefefe4affb8ff1f009700e900;
    decBuf[7793] = 256'h32015b0167015c013e0122010a01f300ec00d900c900b900990073004f002e00;
    decBuf[7794] = 256'h19002c006100a400f700440162017d0185016f016801620172019601c9010702;
    decBuf[7795] = 256'h41028402b202cb02d202cb02a0026d022f020602ef01f60115023d026b028a02;
    decBuf[7796] = 256'h90028b0286027902750287029702bc02e002130343036f039603b003b403b003;
    decBuf[7797] = 256'hac03a903ac03b403c103c403c203c003b303b203b303af03b303b403b903c603;
    decBuf[7798] = 256'he40313043f04660480048e0489046e0464045a0463048004aa04d204f6040d05;
    decBuf[7799] = 256'h09050505fa04f7040005170521052f052c0521051e0524053805550570057305;
    decBuf[7800] = 256'h640544051e050e051305310563059305b205cf05de05ec051b0653068706d306;
    decBuf[7801] = 256'h05070e07f506c10675062f06dd05a605740546051d0507050e052d058105d605;
    decBuf[7802] = 256'h39069706ec062307550782079b07cf07e407ea07e507d507b507970765071907;
    decBuf[7803] = 256'hd306810634060206e705de05e605fb050d0640067006c10624078207d7070e08;
    decBuf[7804] = 256'h18080f080608e107cc07c607d707f10708080308f007d107aa07860779077d07;
    decBuf[7805] = 256'h810792078f078107790772076b077507770765075007360724072e0753078c07;
    decBuf[7806] = 256'hde072b0871089f08b708a1088c086d0851084c0850085d0880088e0881086608;
    decBuf[7807] = 256'h3908f407b4078b075607420748074d0771079b07b707db07f207ff071a082b08;
    decBuf[7808] = 256'h41085b086d0876089008a108be08e008f808eb08d0089b0849081208e007c407;
    decBuf[7809] = 256'hcd07d407cd07c707b6079c0798079c079807b107c707db07fd07140832085508;
    decBuf[7810] = 256'h75089308ae08b1089b087c084d081508ef07db07e107e707ec07d507b7078407;
    decBuf[7811] = 256'h47072e07170710072307340758078207b407e4071d08420857085d084c083208;
    decBuf[7812] = 256'h1208ec07b3078e076c0733070e07d006960662063f06390655068306af06ed06;
    decBuf[7813] = 256'h16071e07400746074c075b0760075c0758074d0737071e07f006b80683065306;
    decBuf[7814] = 256'h34062306280624061f060c06ec05e005d405ca05cd05ca05b705ac059d058f05;
    decBuf[7815] = 256'h8d058b058a058e058d0585058405810586059305b105ce05ea05ed05e405c405;
    decBuf[7816] = 256'h8d0549050905bf048d044d042404f003cd03ba03aa039a038303760372037603;
    decBuf[7817] = 256'h9203bd03ef0312043d045a04690477047b0468044f042004d5037b033e03f102;
    decBuf[7818] = 256'hbf029102790253023f0213020202f301ee01fb010e022e024b025f0269026602;
    decBuf[7819] = 256'h4c022d020602ce01a901860173015701480131011301f800d800c300b800ad00;
    decBuf[7820] = 256'haa00a10099009c00a200ac00bf00c700b70097005100f7ffa3ff56ff38ff2eff;
    decBuf[7821] = 256'h47ff5eff72ff60ff2dffeffeb5fe81fe6cfe66fe6cfe7bfe9bfeb9feccfedefe;
    decBuf[7822] = 256'hdbfed2feb5fe92fe69fe41fe13fee8fdc0fd9cfd8efd82fd76fd65fd36fdeafc;
    decBuf[7823] = 256'ha4fc64fc3bfc42fc65fc91fcc3fcd8fcd2fcb5fc87fc5cfc29fc07fc00fc06fc;
    decBuf[7824] = 256'h0bfc10fc14fc01fce1fbbbfb8dfb61fb3afb0bfbecfad0facbfad0fae5faf8fa;
    decBuf[7825] = 256'hfcfaf9fad9faaafa7efa57fa33fa25fa19fa1cfa27fa1efa04faebf9bcf98cf9;
    decBuf[7826] = 256'h6df946f92cf91ef909f9fdf801f910f930f95ff97ef98ff97ff956f923f9f3f8;
    decBuf[7827] = 256'hbbf8a4f8abf8a5f89ff89af871f83ef80ef8c9f789f770f75af761f774f784f7;
    decBuf[7828] = 256'h94f7b4f7c1f7d4f7edf7f6f7eef7d6f7a7f769f72ff7fbf6e6f6edf6f2f60cf7;
    decBuf[7829] = 256'h2cf730f725f713f7f1f6daf6cdf6c1f6c5f6cef6c0f6b3f6a7f687f667f65af6;
    decBuf[7830] = 256'h3ff626f61df609f6fcf5f5f5ddf5d4f5d7f5dff5f4f514f620f61cf619f6f7f5;
    decBuf[7831] = 256'hdff5dbf5d7f5f7f51df637f64ef652f637f617f6faf5c0f596f571f533f51af5;
    decBuf[7832] = 256'h04f5fdf403f52af544f564f57af566f54ef538f51ef51bf543f576f5a6f5def5;
    decBuf[7833] = 256'hf5f5eef5e8f5c0f592f573f540f510f5fdf4e1f4f1f41af542f565f58ff595f5;
    decBuf[7834] = 256'h85f56ef548f52ef520f51cf537f565f591f5adf5c6f5b8f592f56ef53bf519f5;
    decBuf[7835] = 256'h1ff525f549f57cf590f5b0f5ccf5d1f5d5f5daf5cef5cbf5d4f5d7f5e9f50df6;
    decBuf[7836] = 256'h26f647f65cf650f638f61cf6f1f5caf5baf5adf5b9f5d4f5edf509f624f62ff6;
    decBuf[7837] = 256'h38f64cf654f66ef695f6aef6d8f60bf72df74cf774f76ef761f74bf728f708f7;
    decBuf[7838] = 256'hfbf6f0f601f71df731f750f76ef77af784f787f773f766f76df77cf79af7daf7;
    decBuf[7839] = 256'h1af843f859f852f859f85ef863f87bf898f8acf8cbf8e9f8fcf815f92bf92ef9;
    decBuf[7840] = 256'h26f91ff910f90ef916f928f947f976f995f9bdf9d6f9d2f9cdf9c9f9bff9cff9;
    decBuf[7841] = 256'hfaf932fa75fab5fadffae6faedfadafad5fadafad5fae2faedfaf8fa14fb3ffb;
    decBuf[7842] = 256'h66fb9efbd3fbf5fb08fc0efcfefbf0fbecfbe8fb01fc29fc51fc7ffc9efcaffc;
    decBuf[7843] = 256'hb4fcb0fcb4fccffcf5fc24fd5cfd81fda4fdb6fdc7fdccfddafddffde2fdedfd;
    decBuf[7844] = 256'hfdfd0bfe23fe32fe46fe5efe7afe95feb5fecafeddfeeffe05ff24ff53ff8bff;
    decBuf[7845] = 256'hcffffcff15001d000800f5ffe4ffeafff7ff0d0028004700540067006b006800;
    decBuf[7846] = 256'h6b0073009100c000f8003c017c01b601db01fd011d022e0233022e022a022602;
    decBuf[7847] = 256'h22021f0228022b022d022b02250223022b02390253028d02c702190350039603;
    decBuf[7848] = 256'hc403ed03f503ee03e803e203dd03eb03ef03fb03050408041704190417041904;
    decBuf[7849] = 256'h1f0421042f044d047404b604f6041f05540568056f056905640556055a056605;
    decBuf[7850] = 256'h70059305aa05b705c205c605b005ad05a5059e05b105d305f40522065b068006;
    decBuf[7851] = 256'hb006d006e006f006fe06f106e506e206cc06d506e206f2060a07190711071307;
    decBuf[7852] = 256'h0707fd0607071e0733075f078a07a607c007d707db07ef07f907f607ff070708;
    decBuf[7853] = 256'h00081308250831084d08580855085208490837083e084408420852085c085608;
    decBuf[7854] = 256'h63086b086f0884089e08af08cb08e708f1080d0921092b093b09490941094809;
    decBuf[7855] = 256'h3e092809250918090709120914090b0916091b091709270936093c0956097109;
    decBuf[7856] = 256'h7c099809a309a709bd09c009b809ba09b4099e099b09930987099609a409ad09;
    decBuf[7857] = 256'hbb09bd09ae09a709a1099509a709b809c209dc09f509fe09120a1a0a0e0a100a;
    decBuf[7858] = 256'hfe09db09d609c809bb09c709d809db09ef09f709f009ee09e009c909c609c909;
    decBuf[7859] = 256'hc109d609e509ed09070a180a1b0a240a1c0afd09f109d509b609b209b609b909;
    decBuf[7860] = 256'hcf09e309e609f609f809ee09ed09de09c809c509bd09b109b809b2099f099709;
    decBuf[7861] = 256'h86096a0967096309530962096a096c0988099b09a609b509be09ab09a9099609;
    decBuf[7862] = 256'h79096d094e0930091d090b09fc080a090d090a090c09fa08dc08cf08bb08aa08;
    decBuf[7863] = 256'hba08c208c508da08e308db08dd08ce08b408aa089408740868084d083b083808;
    decBuf[7864] = 256'h3b083d0853085b085408480830080808ec07c807b107b507b107ad07b707b407;
    decBuf[7865] = 256'ha707a9079607790766074d07310726071b071207150712070b070907ff06eb06;
    decBuf[7866] = 256'hde06bf06a2068e067d0673067c067f067c067a066c065506460626060806ed05;
    decBuf[7867] = 256'hce05b005ac05a20598059b0593057e056a054d05320520050405f104e604d704;
    decBuf[7868] = 256'hce04d104ce04cc04ca04be04ac049b04800465044c0436041c0412040204fa03;
    decBuf[7869] = 256'hf203dc03bd03970368033d031503fc02ee02e102e502e802f202f502f202eb02;
    decBuf[7870] = 256'hcf02ac028c02660242023402300224021a020a02fc01e901cf01b00192017701;
    decBuf[7871] = 256'h5e01480134012c011c010d01ff00ef00dc00c400af008f0071004e0037002200;
    decBuf[7872] = 256'h16000500fbffe7ffd5ffc9ffb2ff9cff88ff70ff54ff41ff2fff19ff11ff09ff;
    decBuf[7873] = 256'hfdfef6fee4fed4fec5feaffe9bfe83fe61fe40fe2bfe08fee8fdd3fdb8fd9ffd;
    decBuf[7874] = 256'h8ffd7bfd64fd54fd40fd2efd26fd18fd0efd0ffd07fdf7fce8fccefcaefc99fc;
    decBuf[7875] = 256'h76fc5ffc52fc37fc26fc1cfc08fcfbfbf4fbe1fbc9fbbafb94fb7bfb6dfb57fb;
    decBuf[7876] = 256'h4cfb3afb1efb03fbf2fad5fabafab0fa9afa86fa83fa77fa6dfa6ffa62fa5efa;
    decBuf[7877] = 256'h59fa47fa3bfa35fa23fa09faf7f9d5f9b5f99ff97cf95cf94ff93cf92af92ef9;
    decBuf[7878] = 256'h1ff912f910f9f8f8dcf8d1f8b8f8a2f8a5f89df89bf8a1f897f88bf886f870f8;
    decBuf[7879] = 256'h53f840f821f80bf8f8f7dff7d6f7d3f7c6f7baf7bcf7aaf79af793f77df775f7;
    decBuf[7880] = 256'h72f766f764f766f756f747f73df723f708f705f7f5f6ecf6eff6def6cff6c5f6;
    decBuf[7881] = 256'habf690f68df677f66ef676f66ff671f67ff67af67bf686f679f66ef667f652f6;
    decBuf[7882] = 256'h44f641f630f626f62cf61ff617f616f601f6e7f5ddf5baf5a3f5a8f59cf5a6f5;
    decBuf[7883] = 256'hbcf5bff5c7f5d3f5c8f5c2f5c1f5b2f5acf5b1f5acf5aef5baf5b2f5aef5b4f5;
    decBuf[7884] = 256'ha4f59ef5a0f590f58af588f578f56df573f572f57af58af588f586f581f568f5;
    decBuf[7885] = 256'h5ef561f55ef566f57bf584f591f5a2f5a4f5aef5bef5b7f5b5f5b7f5a8f5a6f5;
    decBuf[7886] = 256'hacf5a4f5a5f5aff5abf5aef5bbf5b3f5aaf5aff5a3f5a4f5b2f5baf5d0f5e9f5;
    decBuf[7887] = 256'hedf5fdf511f619f624f633f631f630f638f62df631f642f644f64ef65af655f6;
    decBuf[7888] = 256'h57f663f665f66ff681f683f68ef69cf6a1f6adf6c3f6ccf6e1f6fdf609f71bf7;
    decBuf[7889] = 256'h30f72ef730f73cf736f73cf748f74df75af76ef775f786f799f79cf7a8f7b7f7;
    decBuf[7890] = 256'hb9f7c5f7d7f7e7f703f826f83df85bf876f879f87cf88bf888f894f8a7f8aff8;
    decBuf[7891] = 256'hc0f8d7f8e7f8fbf812f916f924f931f92ff935f943f94cf95ef978f990f9acf9;
    decBuf[7892] = 256'hcff9e6f9fcf907fa0bfa1afa2ffa3cfa5bfa81fa9afabbfad9fae4faf6fafffa;
    decBuf[7893] = 256'hfcfafafaf7faedfaf3fa02fb15fb32fb5dfb79fb9dfbbdfbd3fbeefbfffb09fc;
    decBuf[7894] = 256'h17fc29fc3ffc59fc7ffc99fca7fcbcfcc0fcc3fcc6fcc9fcd6fce7fcfafc17fd;
    decBuf[7895] = 256'h3afd5afd78fd93fdacfdb5fdbefdcbfde0fdf4fd07fe21fe39fe43fe57fe64fe;
    decBuf[7896] = 256'h70fe7ffe8dfe99fea7febdfed2feeefe0aff29ff47ff5aff6cff82ff90ff9dff;
    decBuf[7897] = 256'haeffc1ffd3fff2ff07001b00330036003f00420049005800660079009000a600;
    decBuf[7898] = 256'hc000d900ef00030115012a013f0151016201750187019801a201b001c701d701;
    decBuf[7899] = 256'heb01fd01090218022602320241024f025b026a02780280028c029c02ab02bd02;
    decBuf[7900] = 256'hce02dd02ef02ff02120325033a034303550366036c037e038f039903ab03bc03;
    decBuf[7901] = 256'hc203cc03d903da03e203ee03f303fe030a04120426043804440457046f047804;
    decBuf[7902] = 256'h8c049904a004af04b904be04c704d104d004d804e304e404ea04f204fb040b05;
    decBuf[7903] = 256'h1605200530053f0545055405630565057505800582058e0599059b05a705af05;
    decBuf[7904] = 256'hae05b705bb05ba05c705d705dd05ef05fb05fd05070610060e06190620061e06;
    decBuf[7905] = 256'h2806320636064706530655065b06590654065c06620664067006780677068606;
    decBuf[7906] = 256'h90069506a406aa06a406a906ae06ac06b506bb06ba06c206ca06cb06d806e606;
    decBuf[7907] = 256'he406e906e706d806da06df06de06eb06f806f90604070807ff060207ff06f206;
    decBuf[7908] = 256'hf406fa06fb06090715071a0727072d0728073207310728072907220717071c07;
    decBuf[7909] = 256'h2607280735073b07320734072d071d071b07150708070a070f07100723073507;
    decBuf[7910] = 256'h33073d073b072f072a0726071f0723071f071407190717071107140715070e07;
    decBuf[7911] = 256'h0c070707000707070a07080710071107040702070007f906f806ef06e006e206;
    decBuf[7912] = 256'he006d806dd06de06d506d906d606cc06d006cf06c506c106bd06b106b606b406;
    decBuf[7913] = 256'hb006b406a70695068e0684067a067b0680067c067d067c0676067b0679066f06;
    decBuf[7914] = 256'h70066806570650064e06480646064106360632062c062406230616060006f205;
    decBuf[7915] = 256'he505d905df05e505e705ec05ed05e605e305dd05d205d005c405b505b705b605;
    decBuf[7916] = 256'hb105b205ae059b05890574055a054f054005310529052705210527052c052e05;
    decBuf[7917] = 256'h3505310523051e0516050e050d050705fd04f804f004df04d304bc0499048204;
    decBuf[7918] = 256'h6d0459045d0460045d04600462046004620464045f045a04460432041f041804;
    decBuf[7919] = 256'h0e0410040a04ff03f103db03bf03ab039a0384037b036e03670369036b036903;
    decBuf[7920] = 256'h6803600354034f034a03440345033f0334032a031d030f030903fc02eb02da02;
    decBuf[7921] = 256'hc302ad0299028b02800279026b025b0255024b02490248024902450246024502;
    decBuf[7922] = 256'h42023e02340228021c020f02fc01ef01e301d801c601b1019d018f0184017501;
    decBuf[7923] = 256'h6f0166015b0156014f014e014d01480143013c01310128011f0113010b010001;
    decBuf[7924] = 256'hf100e700e200dd00d500c900b700a2008e0080007000690063005b0059005800;
    decBuf[7925] = 256'h5900550052004d0041003300250015000a0008000300fbfff4ffeaffdfffd1ff;
    decBuf[7926] = 256'hc1ffaeff9cff87ff72ff6bff63ff66ff70ff75ff73ff72ff6eff62ff55ff45ff;
    decBuf[7927] = 256'h36ff28ff1cff17ff19ff14ff11ff0bff00ffedfedffecafebcfeb9feb2feb0fe;
    decBuf[7928] = 256'haefeacfea4fe9ffe93fe84fe76fe67fe5cfe56fe54fe53fe54fe50fe4afe4bfe;
    decBuf[7929] = 256'h4afe46fe43fe38fe29fe1ffe16fe0bfe09fe05fefafdeffddefdc8fdbafdadfd;
    decBuf[7930] = 256'ha6fda3fd9dfd9ffda7fda9fdaafdaefdabfda4fd9dfd92fd8afd88fd84fd7efd;
    decBuf[7931] = 256'h78fd71fd6afd64fd5bfd50fd48fd39fd27fd25fd1afd1cfd21fd23fd24fd20fd;
    decBuf[7932] = 256'h15fd0efd0cfd03fdfefcfdfcf8fcf6fcfcfcfdfcfefcfdfcf3fce7fcdbfccefc;
    decBuf[7933] = 256'hc2fcbafcacfca7fca8fca4fca0fca6fca3fca0fc9ffc99fc94fc97fc98fc9efc;
    decBuf[7934] = 256'ha9fcabfcacfcb3fcadfca3fc99fc87fc6ffc5ffc4bfc49fc46fc48fc46fc4cfc;
    decBuf[7935] = 256'h47fc45fc49fc4dfc55fc5efc5dfc5efc65fc66fc6efc78fc79fc6efc66fc57fc;
    decBuf[7936] = 256'h49fc3dfc2efc20fc18fc0ffc0bfc12fc18fc22fc2cfc2dfc2cfc2ffc30fc36fc;
    decBuf[7937] = 256'h40fc3efc3dfc3cfc37fc39fc43fc44fc43fc3efc2ffc20fc16fc10fc0cfc0dfc;
    decBuf[7938] = 256'h06fc07fc0ffc14fc20fc2bfc2dfc28fc27fc22fc23fc29fc2bfc2efc2ffc2efc;
    decBuf[7939] = 256'h31fc38fc3afc3bfc38fc2bfc1dfc14fc0cfc0dfc17fc1bfc20fc2bfc33fc3afc;
    decBuf[7940] = 256'h43fc3ffc38fc2ffc22fc1dfc22fc29fc36fc43fc48fc49fc53fc54fc55fc54fc;
    decBuf[7941] = 256'h47fc35fc29fc23fc2dfc40fc52fc63fc72fc70fc6bfc62fc52fc3ffc32fc26fc;
    decBuf[7942] = 256'h2cfc3afc4dfc65fc81fc85fc89fc7ffc77fc6ffc6cfc66fc60fc62fc6afc7afc;
    decBuf[7943] = 256'h8dfc9bfca2fca4fc96fc83fc75fc73fc75fc7bfc80fc8cfc99fc9ffcaafcb4fc;
    decBuf[7944] = 256'hb0fca8fca2fc99fc95fc99fca2fcb4fcc7fccefcddfcebfce9fce4fcdafcc5fc;
    decBuf[7945] = 256'hb1fca9fca2fcacfcbefccafcd9fce3fce8fceafceffceafce9fce8fce5fcedfc;
    decBuf[7946] = 256'hfefc0efd22fd2ffd31fd22fd18fd05fdf8fcf1fce6fce4fce9fcf1fc02fd19fd;
    decBuf[7947] = 256'h29fd37fd3afd33fd2cfd2efd30fd35fd3dfd41fd47fd4dfd4efd4dfd4cfd42fd;
    decBuf[7948] = 256'h39fd32fd2ffd32fd3afd3ffd48fd51fd55fd5afd63fd67fd69fd6afd67fd64fd;
    decBuf[7949] = 256'h67fd69fd75fd83fd85fd84fd85fd81fd7ffd81fd7dfd7cfd7ffd7afd7afd7efd;
    decBuf[7950] = 256'h81fd87fd8ffd90fd93fd9bfda2fdabfdb7fdbbfdbffdc8fdcbfdd0fdd5fdd2fd;
    decBuf[7951] = 256'hccfdc2fdb6fdaefdaffdb6fdbffdcbfdd0fdd2fdd6fddafdddfde4fde8fdeffd;
    decBuf[7952] = 256'hf5fdfbfd06fe12fe19fe1afe19fe14fe11fe10fe11fe15fe1ffe23fe24fe2afe;
    decBuf[7953] = 256'h2ffe35fe3dfe40fe41fe42fe41fe45fe4bfe50fe54fe5afe5ffe61fe66fe67fe;
    decBuf[7954] = 256'h6dfe75fe7afe81fe8dfe98fe9ffea4fea5fea1fe9cfe9afe9bfea4feaefeb7fe;
    decBuf[7955] = 256'hbffec2fec6fecafecdfed1fed4fed5fed6fedefee8fef4fefffe07ff08ff0aff;
    decBuf[7956] = 256'h06ff05ff0bff11ff18ff1eff26ff36ff47ff52ff54ff52ff47ff36ff34ff36ff;
    decBuf[7957] = 256'h3fff4dff5fff70ff7fff89ff92ff96ff95ff8eff88ff82ff85ff92ffa4ffbeff;
    decBuf[7958] = 256'hd0ffd9ffe2ffe5ffddffd3ffc5ffb9ffb0ffafffbbffd0fff0ff0e0021002500;
    decBuf[7959] = 256'h28001f00170010000e0014001d002f00490061007700860088007c006d005f00;
    decBuf[7960] = 256'h57004f0053005d006d0080009200a800b600be00b700a800960094009e00b000;
    decBuf[7961] = 256'hcf00ed0000011201210124011c010c01fd00eb00e400e200ec00ff0017012c01;
    decBuf[7962] = 256'h3b0143014a014c01460141013901370143015c017b019901ac01b701b401ab01;
    decBuf[7963] = 256'h9901880175016d01660171017f019901b401cd01dc01e501e201db01d501d301;
    decBuf[7964] = 256'hd401dd01e401f00102021302260233023102260218020502f801fa01fc010602;
    decBuf[7965] = 256'h1602250237024c025b0263026a025f025102480247024b025502650274028202;
    decBuf[7966] = 256'h8e0296029e029c029402870279027302740280028d02a102ae02b502bf02c902;
    decBuf[7967] = 256'hcb02ca02c502b902b102af02b602c602d502e702f302f502ef02f102e902de02;
    decBuf[7968] = 256'hdd02de02df02e802f8020703190325032703290324031c03170313030b030903;
    decBuf[7969] = 256'h08030d031a032803340340033e03370331032b0326032b0333033a0347035703;
    decBuf[7970] = 256'h620370036e036303580349033b033d033e0343034f0357035c036b0375037703;
    decBuf[7971] = 256'h75036e036103590358035c036a0376037b03820381037d037c0379036f036e03;
    decBuf[7972] = 256'h6d036c03710377037903810382037d037c037c037703760374036e0370037303;
    decBuf[7973] = 256'h75038303910399039e03a0039903900388038103820385038403860387038303;
    decBuf[7974] = 256'h80037a036f036703620364036f037903830393039e03a003a203a30399038f03;
    decBuf[7975] = 256'h8403760371036f0371037d038503870386037d0370036c036403600361036903;
    decBuf[7976] = 256'h72038203950398039a0390037e03720367035d03630367036903700374037203;
    decBuf[7977] = 256'h730371036703600355034b034c034d034e035703600366036d036f036d036803;
    decBuf[7978] = 256'h620359034f0346033c033d033f033e03430345033f033b0335032b0324031e03;
    decBuf[7979] = 256'h160319031f03270333033b0340034403430336032b031b0307030003f402ed02;
    decBuf[7980] = 256'hf302000308030c030b030203fc02f502ec02e802e402dc02e102e502e802ee02;
    decBuf[7981] = 256'hed02e402dd02d402c302b702b102a702a502a702ab02b202bd02c202c602c002;
    decBuf[7982] = 256'haf029e02940286027d027b0277027e02810285028c028d028102760268025202;
    decBuf[7983] = 256'h4202390237023902440252025b025f025b025a024c02350225021d0210021202;
    decBuf[7984] = 256'h18021e0224022902210217020702f001e001cc01ba01b301b501bf01d201e401;
    decBuf[7985] = 256'heb01ee01e801d401c201b1019e0196018f0191019701a0019e0197018b017501;
    decBuf[7986] = 256'h67015501440139012f012e0133013d01470154015a0152014401310119010a01;
    decBuf[7987] = 256'hfb00f300f100f300f500fa00f900f100ea00da00c300ad0099008c0080007e00;
    decBuf[7988] = 256'h80008c009400980097008e0080006e005d004e00480043004100430044004000;
    decBuf[7989] = 256'h3d00300020000d00fbffeaffdbffd1ffc9ffc7ffc8ffcdffd3ffd6ffd5ffd1ff;
    decBuf[7990] = 256'hc5ffb7ffa9ff9dff94ff8dff86ff82ff7dff74ff68ff5eff4fff45ff39ff30ff;
    decBuf[7991] = 256'h2cff25ff21ff1eff1fff1cff1dff1cff1aff14ff0afffbfeedfee1fed2fec8fe;
    decBuf[7992] = 256'hbcfebafeb6feb4feb0feadfea4fe99fe8bfe7ffe74fe6cfe68fe6cfe6ffe6cfe;
    decBuf[7993] = 256'h68fe62fe5afe50fe49fe3efe33fe29fe21fe1bfe16fe12fe0cfe07fefefdf1fd;
    decBuf[7994] = 256'he9fde2fdd8fdcdfdc2fdbbfdb8fdb4fdb5fdb8fdb5fdb1fdabfd9ffd97fd90fd;
    decBuf[7995] = 256'h86fd80fd78fd71fd67fd66fd5dfd55fd4efd46fd3ffd38fd2afd20fd1ffd1dfd;
    decBuf[7996] = 256'h1ffd23fd24fd25fd22fd17fd0bfdfefceefcdffcd9fcd0fcccfccdfcccfcc8fc;
    decBuf[7997] = 256'hcbfcc6fcc4fcbffcb7fcb6fcb7fcb1fcadfcacfca6fca1fca1fc95fc8afc7ffc;
    decBuf[7998] = 256'h73fc68fc60fc56fc55fc59fc5cfc60fc68fc67fc62fc5dfc52fc4dfc4ffc4dfc;
    decBuf[7999] = 256'h4efc54fc51fc4dfc4cfc42fc36fc31fc23fc17fc12fc0efc0ffc18fc19fc1afc;
    decBuf[8000] = 256'h20fc1ffc20fc21fc17fc11fc0ffc05fc01fc07fc0bfc10fc18fc16fc13fc11fc;
    decBuf[8001] = 256'h04fcfafbf4fbe9fbe5fbebfbeafbf2fbfdfbfffb03fc06fcfffbfafbfafbf3fb;
    decBuf[8002] = 256'heffbf4fbf5fbf9fb00fcfffbfefbfbfbf2fbe8fbe4fbd8fbd9fbe1fbe0fbe3fb;
    decBuf[8003] = 256'hebfbeefbf4fbfcfbfbfbfcfbfdfbf3fbeffbf0fbedfbeefbf2fbf3fbf9fb01fc;
    decBuf[8004] = 256'h02fc05fc05fcfbfbf4fbf3fbebfbeefbf9fb01fc09fc0dfc0efc0ffc14fc12fc;
    decBuf[8005] = 256'h13fc17fc14fc15fc1afc19fc1bfc25fc29fc2ffc37fc36fc35fc3afc34fc2ffc;
    decBuf[8006] = 256'h30fc2ffc34fc3cfc3ffc46fc51fc56fc5bfc67fc69fc6dfc71fc70fc71fc78fc;
    decBuf[8007] = 256'h79fc7ffc89fc8dfc93fc9dfc9cfc98fc97fc90fc91fc97fc9ffcaefcc0fccbfc;
    decBuf[8008] = 256'hdafce4fce6fce8fce9fce8fcecfcf1fcf2fcf8fcfefc03fd09fd14fd19fd21fd;
    decBuf[8009] = 256'h28fd29fd2cfd31fd34fd3afd44fd4afd58fd64fd70fd7dfd86fd84fd80fd81fd;
    decBuf[8010] = 256'h80fd86fd91fd9bfda5fdb0fdbbfdc4fdcdfdd3fdd8fddcfdd8fdd7fdd8fdd8fd;
    decBuf[8011] = 256'he0fdeffdfdfd10fe23fe2efe35fe37fe32fe33fe35fe3cfe49fe5dfe6afe71fe;
    decBuf[8012] = 256'h77fe79fe7efe7dfe7efe80fe86fe8cfe95fea2feaffebdfecbfed7fee3feeafe;
    decBuf[8013] = 256'heefef2fef1feeefef1fef9fe00ff09ff15ff1fff26ff2fff34ff3bff43ff4bff;
    decBuf[8014] = 256'h56ff5eff67ff70ff78ff81ff8cff97ffa3ffa8ffa9ffa8ffa9ffaaffb1ffb9ff;
    decBuf[8015] = 256'hc6ffd4ffe2fff2ff0100070010001100130017001d0023002a00300038003b00;
    decBuf[8016] = 256'h42004c005300590063006a00730078007f008b0093009a00a400af00b400bb00;
    decBuf[8017] = 256'hc100c200c500cb00d500e100ec00f400fb00ff000001030105010b0113011b01;
    decBuf[8018] = 256'h24012d012e01310139013f0146014f0156015c0164016b01710177017c018001;
    decBuf[8019] = 256'h86018b018d019301980199019f01a101a801b301bb01c001c601c501c901d201;
    decBuf[8020] = 256'hda01e401f101f601f701fb01fd01fb010002030206020e021102120216021902;
    decBuf[8021] = 256'h1c022302290230023d0247024c0251025002510257025d0264026e0272027302;
    decBuf[8022] = 256'h7902780277027902790278027e02820285028b028c028b02910294029802a202;
    decBuf[8023] = 256'ha902ac02b602bb02be02c802cd02d302db02dc02d702da02db02da02de02df02;
    decBuf[8024] = 256'hde02e302e202df02e402e402e502ed02ee02ed02f502fb0202030d0315031703;
    decBuf[8025] = 256'h1b031c031d0322032303210321031f0319031b031a0318031c031f0320032803;
    decBuf[8026] = 256'h2d03300338033b033a033d033c033b033e033d0339033b033e033f0348034a03;
    decBuf[8027] = 256'h4b034c0345034103420341034203460349034a034e03510351035b035f035e03;
    decBuf[8028] = 256'h5f03580350034d034603410348034e03540361036703650364035f0355035403;
    decBuf[8029] = 256'h5303520356035703550359035a0357035c035d0358035703560354035a035d03;
    decBuf[8030] = 256'h5d03620363035e035d035d0358035b03560350034f034f034e03500353035003;
    decBuf[8031] = 256'h510350034f0352035303500353034f03480346034003360332032e032d033203;
    decBuf[8032] = 256'h36033b033d033d033603340331032d032e032d032803260323031f031c031a03;
    decBuf[8033] = 256'h150313030c030103fc02f802f602fa020003030305030303fd02f802f402ec02;
    decBuf[8034] = 256'he902e202da02d402cf02cb02c602c402be02bb02b802b202b302b002a902a302;
    decBuf[8035] = 256'h9e029a029c029f029e029b02930287027c0271026a0267026502620262026202;
    decBuf[8036] = 256'h5c025a02520245023a02300223021e021d0219021a021d021a02190219021102;
    decBuf[8037] = 256'h0b020202f701ec01e501dd01d701d201ca01c501be01b401aa01a4019a019601;
    decBuf[8038] = 256'h92018c018901870182017e017b0174016e0169015e01520148013b0130012801;
    decBuf[8039] = 256'h1f01190113010c0106010001fa00f300ef00e900e300dd00d700d000d000c900;
    decBuf[8040] = 256'hc200b700a8009a00920086007f007b0072006a006300590052004f0049004400;
    decBuf[8041] = 256'h400038002b00200016000f000d000c000b0007000100f5ffeaffddffd0ffc8ff;
    decBuf[8042] = 256'hbeffb1ffa9ff9fff98ff92ff8aff7fff77ff70ff68ff62ff5fff57ff54ff51ff;
    decBuf[8043] = 256'h4eff4dff4bff44ff37ff29ff16ff09fff8feeefee4fedbfed0fec8fec4fec3fe;
    decBuf[8044] = 256'hc4fec7fec6fec3febdfeb4feaafea1fe95fe89fe82fe78fe6dfe66fe5cfe53fe;
    decBuf[8045] = 256'h4bfe42fe3cfe36fe2ffe2dfe2afe26fe23fe21fe1afe13fe0bfefefdf5fdeafd;
    decBuf[8046] = 256'he2fddbfdd5fdcffdcafdc9fdc3fdbffdbbfdb4fdaefdacfda4fd9cfd99fd8ffd;
    decBuf[8047] = 256'h88fd85fd7dfd76fd70fd64fd5cfd5bfd59fd58fd5efd5dfd58fd57fd51fd4bfd;
    decBuf[8048] = 256'h49fd41fd3bfd36fd2bfd1ffd15fd0bfd05fd04fd01fd00fd03fd02fd03fd07fd;
    decBuf[8049] = 256'h06fd07fd08fd05fd01fd00fdfafceefce6fcd6fcc7fcc1fcbcfcbdfcc5fcc9fc;
    decBuf[8050] = 256'hcdfcd0fccffccefcd3fcd3fcd4fcd7fcd1fccbfcc6fcbdfcb3fcaffca7fca2fc;
    decBuf[8051] = 256'ha2fc9dfc9bfc9ffca0fca4fcb0fcb4fcb6fcbafcb4fcaefcabfca5fca1fca3fc;
    decBuf[8052] = 256'h9ffc9cfca1fc9cfc9bfc9cfc9afc97fc9afc9bfca1fcaafcaefcb2fcb8fcb7fc;
    decBuf[8053] = 256'hb4fcb7fcb1fca9fca3fc9afc94fc95fc94fc97fca4fcaafcb3fcc1fcc7fcc9fc;
    decBuf[8054] = 256'hd1fccdfccefcd2fccefccffcd4fcd3fcd0fcd5fcd4fcd3fcd7fcd6fcdbfce4fc;
    decBuf[8055] = 256'hebfcf4fc00fd05fd07fd0efd11fd15fd1cfd1dfd18fd17fd11fd0ffd16fd1efd;
    decBuf[8056] = 256'h29fd3afd40fd4afd53fd55fd59fd60fd61fd65fd6afd69fd68fd70fd75fd7efd;
    decBuf[8057] = 256'h8cfd91fd96fd9bfd99fd9dfda5fdaafdaefdb8fdb9fdc0fdcafdd1fddcfde9fd;
    decBuf[8058] = 256'hf2fdfafd02fe06fe0afe0dfe08fe05fe08fe0bfe12fe21fe2ffe3bfe47fe51fe;
    decBuf[8059] = 256'h58fe5efe62fe63fe65fe64fe64fe68fe69fe71fe7ffe8dfea1feb3febffecefe;
    decBuf[8060] = 256'hd4fed2fed0feccfec5fec1fec5fec6fecdfed8fedefee7fef1fefbfe09ff1cff;
    decBuf[8061] = 256'h29ff3aff40ff42ff44ff45ff44ff45ff44ff41ff3cff3dff3dff45ff56ff67ff;
    decBuf[8062] = 256'h76ff88ff98ffa3ffa9ffaeffadffaeffadffaeffafffb0ffb1ffb0ffb1ffb5ff;
    decBuf[8063] = 256'hbfffc9ffd6ffe3ffebfff5ffffff0a00180024002c003300350039003a003700;
    decBuf[8064] = 256'h32002c00260022001f001e002100290035004a005e007b008f00a000a900ac00;
    decBuf[8065] = 256'haf00ad00aa00a000940089007e00750076007e008d00a000b200c300d200dc00;
    decBuf[8066] = 256'he100e300e100dd00d700cf00ca00c700ca00cd00d400da00e300ee00fc000801;
    decBuf[8067] = 256'h170121012601280126011c0114010701f900ef00e900eb00f9000c011e012f01;
    decBuf[8068] = 256'h3e014401490147013d01330125011d0118011c012601360145014b0150014b01;
    decBuf[8069] = 256'h4101350129011f012301290131013e014a01560163016c0171016f0168015801;
    decBuf[8070] = 256'h49013b0132012e012c012b013101370140014d015d01680176017b017d017e01;
    decBuf[8071] = 256'h74016401550143012e012501230120012b013d0152016c0185018e0197018f01;
    decBuf[8072] = 256'h790165014e013e0130012d012b012d01370140014e015c0165016d0175017901;
    decBuf[8073] = 256'h7a017b0174016c0160014e013d012e011c0115011301150128013b0150016401;
    decBuf[8074] = 256'h710174017a0178017601750173016a01610159014a0144013a012d0122011201;
    decBuf[8075] = 256'hfe00f700ef00f60008011d013701570174018f01a101aa01a2018f0170014a01;
    decBuf[8076] = 256'h26010601e000c600b800ab00b700d000ec0016013e01620179018e019a019601;
    decBuf[8077] = 256'h8601610133010701e000c600b800b400c000d800ee000e012301360148014b01;
    decBuf[8078] = 256'h42013501290116010e010c01060108010901040106010a010e0116011d011a01;
    decBuf[8079] = 256'h1701100108010301fe00f600ef00e800e100e900fa0010012401310133013101;
    decBuf[8080] = 256'h270117010801f200de00d100d400e700090132014f015e0150013b011001e900;
    decBuf[8081] = 256'hbb009b008b0085009d00c300fb00300160017f0185018001680142011e01eb00;
    decBuf[8082] = 256'hc900b600a500ab00c200d700f2000b011a0123012b012d012b01290124011f01;
    decBuf[8083] = 256'h1a0113010d010a0103010001ff000501130129013d0154015e015b014e013801;
    decBuf[8084] = 256'h1901fb00d800c100ac00b000ba00dc0006012d0151016801750181017d017401;
    decBuf[8085] = 256'h6b015e014e014301350122010a01f400e000ce00c700c900d300e600f8001201;
    decBuf[8086] = 256'h320150016b018a019701aa01b501b201af01a7019201720143010b01d700a600;
    decBuf[8087] = 256'h870082008700a700de0022016201ac01f2010d0226022e020b02df01ad016f01;
    decBuf[8088] = 256'h3501f200c400ab00a400b800e4000c0144017801a901c801ef01ff01f101d301;
    decBuf[8089] = 256'h99015f012b010801020108012101420170019c01c301dd01d801c30199017101;
    decBuf[8090] = 256'h4d01360129012d0138014701610181019f01b201b501a601970190018d019401;
    decBuf[8091] = 256'h9a0198018c017c017101670169016b01690168016401630168016b0166016201;
    decBuf[8092] = 256'h55014b014c015e017d01a301c701de01f401f001de01bc0180013601f000c200;
    decBuf[8093] = 256'h9900af00df0018016a01b701e90104020d02f601c6018e013b010401d200c900;
    decBuf[8094] = 256'he20007012a0149015a0169016e017b017f017b0178016f01670165015a014401;
    decBuf[8095] = 256'h1901e100ad008a009000b800f00034018601bd01db01e401dc01a7015c01ee00;
    decBuf[8096] = 256'h86005e003a0045007700b700e000140129012f012a011001e600bf00a500b300;
    decBuf[8097] = 256'he20027016701a001a80193015b01fa009c001700bdff4bff1fff2dff69ffccff;
    decBuf[8098] = 256'h5f00c1003f019001bc01e401c0019f014501f0008d002f00daff8dff5bff40ff;
    decBuf[8099] = 256'h38ff3fff6fffc1ff24006700a300da00e400ed00e500cf009e005a001a00d0ff;
    decBuf[8100] = 256'hb2ff84ff7cff74ff6dff74ff84ff9effb5ffdbfff5ff03000700fcfff1ffe8ff;
    decBuf[8101] = 256'hd4ffbcffa0ff85ff6cff69ff6cff69ff6cff61ff57ff4eff46ff45ff49ff4fff;
    decBuf[8102] = 256'h59ff68ff76ff83ff8bff7dff63ff29ffdffeadfe7ffe77fe7efea1feccfefffe;
    decBuf[8103] = 256'h3dff77ff9cffa3ff84ff46ffebfe96fe49fe2bfe22fe3bfe51fe74fe93fea4fe;
    decBuf[8104] = 256'hb3feaffea2fe87fe75fe72fe75fe87fe98fe9afe8cfe75fe59fe46fe34fe25fe;
    decBuf[8105] = 256'h16fe09fe02fe0dfe27fe3ffe55fe58fe40fe1efef4fdcdfd9ffd73fd4cfd32fd;
    decBuf[8106] = 256'h37fd5dfda0fdf2fd55feb2feeffe10ff06ffd8fe8efe0cfe6bfdd4fc4afcf1fb;
    decBuf[8107] = 256'hc0fbcffb12fc67fccafc5dfde6fd63fed5fe1fff2cfff0fe77fe05fe80fd03fd;
    decBuf[8108] = 256'hb2fc86fc78fc84fca5fcc3fcccfca3fc6ffc23fcf1fbe8fb32fca0fc42fd05fe;
    decBuf[8109] = 256'h88fefefe6bff57fffefe4bfe75fd72fc7efbe0fa8afaa4faebfa2cfbb5fb56fc;
    decBuf[8110] = 256'hc2fc4cfda5fdf6fd23fe15fef1fdd0fd9efd5efd14fdcefc7cfc2ffcfdfbcffb;
    decBuf[8111] = 256'hb6fba0fb99fbacfbdefb2afc98fcfffc42fd66fd71fd53fd38fdfefcd9fcb6fc;
    decBuf[8112] = 256'h97fc86fc77fc69fc65fc61fc4ffc3afc20fc07fcf8fb00fc13fc36fc5afc8dfc;
    decBuf[8113] = 256'hbdfce9fc10fd20fd1bfdf5fcb2fc72fc28fcf6fbdbfbe3fbf9fb29fc7bfcc8fc;
    decBuf[8114] = 256'h22fd46fd3bfdf5fc7efc0dfca5fb63fb3efb75fbbbfb44fccdfc4bfdbcfdcbfd;
    decBuf[8115] = 256'ha3fd4efdd5fc63fcfcfbb9fb95fba0fbd2fbfffb4afc90fcbdfce7fceefcd9fc;
    decBuf[8116] = 256'hbafca9fc9afc95fca2fcaefcbffcd5fcd8fcd5fcbbfc8efc55fc21fcfffb05fc;
    decBuf[8117] = 256'h37fc91fcfefc65fda8fdb4fd93fd39fdccfc47fccafb79fb6afb92fbfffba2fc;
    decBuf[8118] = 256'h39fdeafd60fea1fe8efe58fee6fd62fdc1fc29fcc7fb92fb81fb90fbeefb5bfc;
    decBuf[8119] = 256'he0fc5dfdcefd18fe26fe19feccfd5efdf7fc9afc75fc96fcdcfc53fde5fd47fe;
    decBuf[8120] = 256'ha1feb1fe67feeffd3cfd66fc9dfbe6facefae4fa95fb9afcd4fdfbfe07007000;
    decBuf[8121] = 256'hcf007800c2ffbcfe82fd5cfc4ffbe6fac7fa1dfbd4fbaafcacfd5bfebafe10ff;
    decBuf[8122] = 256'h2affe3fecdfeb9fea8feb8fec7feb9fe95fe32feb9fd27fdc5fc6cfc3bfc67fc;
    decBuf[8123] = 256'hc5fc4afdebfdaefefcfe73ff88ff9cffaeff9eff71ff49ff25ffd8fe7efe11fe;
    decBuf[8124] = 256'haafd4cfdf7fcc0fcb6fcd1fc1cfd8afd0efeaffe72ff2900cf006601c901b701;
    decBuf[8125] = 256'h650188006cff5ffe25fdfefb8bfb68fb06fc09fd43fe6affc300ab01d501af01;
    decBuf[8126] = 256'h46016900a0ffe9fe72fe5cfe97fef1fe83ffe5ff3e004f004000c7ff56ffd1fe;
    decBuf[8127] = 256'h54fe03fe11fe54fef2feb4ffa0007d010d025b024302d701ff0036004bffadfe;
    decBuf[8128] = 256'h57fe71fee7feaaff6100d800190105018800d5ff2fff97fe5dfeb6fe69ff6e00;
    decBuf[8129] = 256'ha801cf028f033d041d04540369020d01c8fff6fe36fe13fe72fe02ffb9ff8e00;
    decBuf[8130] = 256'h1e016c01b40173015f012a01190146018801f6017a02d402e402d5027802da01;
    decBuf[8131] = 256'h17019500eeffaeffc1ff1b008c0011018e0100024a0272027e02730269026002;
    decBuf[8132] = 256'h37022002fe01de01e401f301260264029e02c302bd02840214028201d1002b00;
    decBuf[8133] = 256'hbfffd2ff2c00ff003b026203bb04a3052206fb054d05f103ac02850179001000;
    decBuf[8134] = 256'h6f00ff00ea01c7029103df03c7035b03d20231029901370149019a015a024503;
    decBuf[8135] = 256'h2304ec04a305ea05a905470582049703ba02f101a2018b01a00102027f02d102;
    decBuf[8136] = 256'hfd02f002cb0294028a02ca0246032e040c0548061a0741071e0780064405c803;
    decBuf[8137] = 256'h6302c2001a0081ff0c00de00eb0125034c045805c10520060306b5059d058705;
    decBuf[8138] = 256'h7405860596056a050c056e04810364025701a9008900a6009101ed028e041706;
    decBuf[8139] = 256'h7c076408e308bc08c8076c062805ac034702bc013e0164011302b102b403a804;
    decBuf[8140] = 256'hc4058406ed060c07b606ff05fa040604e90276025302f102f4037405d9061d08;
    decBuf[8141] = 256'h44096b09bc08210728054c039c018300500038010703b804b1060508be081608;
    decBuf[8142] = 256'h17077505ec038702fc017b023b03ba041f06c107d9080c093b09bc08b0073006;
    decBuf[8143] = 256'hcb048603b4024102630202033e046505be0603088108f408d10833083007f705;
    decBuf[8144] = 256'hd004c3031503f5024b030204d804db05cf066d07c307dd07c607b0074e071807;
    decBuf[8145] = 256'he706d906b106a4066d064f0634062c06330663068f0695067b063606b4051305;
    decBuf[8146] = 256'ha7046c04a20434050c06d506c0075e08b4089a0853081208b0077a074a073b07;
    decBuf[8147] = 256'hf806bb066e060006b7058f058205b905ff056406dc064e07b507f807d4078707;
    decBuf[8148] = 256'h05076406f805e4053d06d006a8077108f3080b099f08a0076606eb04ec036103;
    decBuf[8149] = 256'h8b034b048505540704091d0ab60ae40a660a0d096b07e2057d049503c0037f04;
    decBuf[8150] = 256'h740590065007fe07df07c2073f07c9065d0649065b068c06f30636075a076507;
    decBuf[8151] = 256'h3307e1067e062006cb05aa05a005ce05f7052c062506e0057c051e05c904d404;
    decBuf[8152] = 256'h2e05e405cf06ad077608c408dc089b08c307c106870560045303a5028502a202;
    decBuf[8153] = 256'hf002970359041005b605220636062406d3054e05d1048004540461048504a604;
    decBuf[8154] = 256'hc404e004d704df04d804d204c1047e041a048703d6023002c401620174010602;
    decBuf[8155] = 256'hde021a04ed04f9051c06bd05f404d5032e02a600a7ffbffe40fe67fecffeadff;
    decBuf[8156] = 256'he90010021c0311046f04530404048e03cb0214026e010201ee000001f000e100;
    decBuf[8157] = 256'h6900b6ffe0fe17fe94fd4dfd8efd3efe14ffa4ffbeffa6ff0fff5efe89fdf9fc;
    decBuf[8158] = 256'hdffc55fd43fe9fffe4000b027e02a10203028d00c2fe96fc8bfa37f97ef8b6f8;
    decBuf[8159] = 256'hb5f9f9fa20fc93fcfcfcdcfcf9fc13fd8afdf6fd7ffe6efefcfd1ffd44fb68f9;
    decBuf[8160] = 256'hb8f79ff606f691f664f70af993faf8fbe0fc5efd38fdcffc31fc68fbb1fa0bfa;
    decBuf[8161] = 256'h73f939f9dff86df8e9f700f723f693f511f558f51af606f722f8e2f890f971f9;
    decBuf[8162] = 256'h54f969f88cf789f6daf53cf520f5a2f578f641f72cf88bf835f8b2f7adf673f5;
    decBuf[8163] = 256'hf8f3f9f26ef244f2b7f2abf3c8f4d4f5c8f667f710f725f6c9f428f39ff1a0f0;
    decBuf[8164] = 256'h72f044f19ef2f9f438f7aef87af9c1f8c8f664f4dbf090ed6deb09eb64eba4ed;
    decBuf[8165] = 256'h44f073f396f588f72df737f62bf4c7f12cf0b6eefaeeb4ef3cf107f3b8f460f5;
    decBuf[8166] = 256'h2df545f476f24af03feeebec32ec6aeccfed13ef8ef0f3f1dbf25af3e7f27ef2;
    decBuf[8167] = 256'ha1f1d7f020f0aaef3eefdbee82ee51ee08eedfed34eed9eedfef5ef1c3f2abf3;
    decBuf[8168] = 256'h29f403f40ff3f2f199f054ef82ee5bee7eeeddee33ef82ef6aeffeee9ceefbed;
    decBuf[8169] = 256'h8fed54ed42ed52edb9ed82ee85efbff0e6f13ff327f451f4def3eaf2cdf174f0;
    decBuf[8170] = 256'h8cef0defe7ee0aef69efbfefd9ef20f036f04af038f0e7ef62efe5ee93eea2ee;
    decBuf[8171] = 256'h35ef34f06ef195f255f3bef39ef3d5f2eaf1cdf00df0eaef0af09af051f1f7f1;
    decBuf[8172] = 256'h0cf2f9f19ff14ef13ff182f108f2ccf2b7f395f45ef5e1f5c9f55df536f4bbf2;
    decBuf[8173] = 256'hbcf1d4f0aaf01df1ccf1ebf108f222f2dbf11cf2a5f26af355f472f57ef6b8f7;
    decBuf[8174] = 256'h8bf84bf96ef90ff9d2f757f68cf4dcf2c3f12af1fcf07af187f292f49df601f9;
    decBuf[8175] = 256'h41fb21fc65fcacfb23fa58f8a8f68ff590f405f4dbf39bf4d5f550f7b5f8faf9;
    decBuf[8176] = 256'h24fa4afae2f983f99ff9eef965fafcfa5efbb7fba7fb40fb77fa02f99df711f7;
    decBuf[8177] = 256'he7f6f4f7b9f9e5fb5bfdaffeedfe25fff2fec3fe99fed9fd9ffc24fbbff9d7f8;
    decBuf[8178] = 256'h59f8ccf87bf9d6fa1bfc42fd9bfee0ffb30026010301e300c60078006000f4ff;
    decBuf[8179] = 256'h6bff82fea5fddcfc59fc12fc53fcdcfce8fd8efff8013804ad0579063c064204;
    decBuf[8180] = 256'h66023b002ffe63fda1fd4afeaffff3006e02d303bb043a057a0440031c0111ff;
    decBuf[8181] = 256'h45fe07feb0fe7b0022039b05db07e609b20a750a5c0991076505ef0313025a01;
    decBuf[8182] = 256'h22015501e0010703ad04a606fa07380890079106ef04d7033e030f033903ad03;
    decBuf[8183] = 256'h1504f3042f06fe07ae09370b9c0ccb0c4c0c400b060a8b0826078405fb036203;
    decBuf[8184] = 256'h91036304560632085e0a3e0b0a0c510ba90a4409ff07d8061806b0050f064b07;
    decBuf[8185] = 256'h7208cb09b30a310b580b350bd60a800a310a1a0ad909ec09690afc0a850b970b;
    decBuf[8186] = 256'h050bde09b708ab0788076508db09a60bdb0cf30d260e9b0d200cbb0a1a099107;
    decBuf[8187] = 256'hf80626074d08f3097c0b7b0c060d300d710c080ce80bcc0bb10bc90bb40bee0b;
    decBuf[8188] = 256'h480c990c000d0e0dd10c420c910bbc0a2c0ade099609ac09350afa0ae50b020d;
    decBuf[8189] = 256'hc20d700e900e730e240edd0d710d0f0d6e0cab0b290be20af70a320bfc0a8b0a;
    decBuf[8190] = 256'he80951096509710a640cc80e07117d1239128011f70f2c0e7c0cf30a5a0a880a;
    decBuf[8191] = 256'h070b600ca50dcc0e3f0fd60eb90dc70b730a3e090609050a030cdf0d0b108011;
    decBuf[8192] = 256'h3c1183108a0eae0c790bd10a040b480c6f0d7c0ee50e430f270f410f590f6e0f;
    decBuf[8193] = 256'h0c0f8f0edc0d950dab0d340ef90e7b0f340f1b0ec10c200b780a450a2d0bfc0c;
    decBuf[8194] = 256'hac0e351034116211381178103f0fc30dc40c390c0f0c820c760dd20e17109211;
    decBuf[8195] = 256'h9112bf124112e810ea0e0e0d5d0bb50ae80a730b9a0c5a0d4e0e2b0ff50fe010;
    decBuf[8196] = 256'hfc11bc129912fb11bf10440fdf0df70c790c520c2f0c4f0c6c0cee0c950dae0e;
    decBuf[8197] = 256'h0710ef101612d6123e135e1308131d123f11c90f640e200df90b390b5c0bbb0b;
    decBuf[8198] = 256'hf70c720e3d10ed110613d3128e11bf0f930d1e0cda0b170ca00d6b0f1b11c411;
    decBuf[8199] = 256'h5d122e12b0113d118f10f00f270f3c0e5f0d5c0cae0b8e0b1e0c090da40e2d10;
    decBuf[8200] = 256'h9211d61255137b13cd12b0110a10110e350c090a2909e5081a0a130c770eb710;
    decBuf[8201] = 256'h9711db112211990f340eef0c710ce40cd80db50eb80f21100110380f180ebf0c;
    decBuf[8202] = 256'hd70b050b2b0b940b710c740d220e810ef10d060d2c0b50091b087307a607ea08;
    decBuf[8203] = 256'hba0ae50c5b0eaf0f681081111a12ec116d117a0f160d320ab306590435020b01;
    decBuf[8204] = 256'hb000020178025404fb062a0a4d0c060fca101d11fd11b9110011770f120eb70b;
    decBuf[8205] = 256'hd3081a06ec02edfffcfd37fce5fbc5fc29ffb202fd05fb08b40bc30c150d350c;
    decBuf[8206] = 256'hf10bbc0ac308e706bb0446037a023c02e4027d03ac032d036d02bf0160014301;
    decBuf[8207] = 256'h5e0175010901ce00e000720199021404130541051705be037902aa00fafee1fd;
    decBuf[8208] = 256'h48fd1afd98fd58fe4cffeaff4000beff17ff80fef7fdc1fd90fd82fd74fd80fd;
    decBuf[8209] = 256'hb7fd39feb6fe08fff9fe66fe67fd73fc56fb49fa9bf9fdf8a7f88cf8d4f815f9;
    decBuf[8210] = 256'h77f989f958f90ef91bf989f948fa33fb92fb76fbbffab9f9c5f866f883f89df8;
    decBuf[8211] = 256'h56f893f7a8f68cf57ff416f4f7f3daf3f4f30cf422f484f401f593f544f619f7;
    decBuf[8212] = 256'h1cf8cbf869f912f927f84df671f4c1f238f19ff0b7ef90ee83ed4aec1fec79ed;
    decBuf[8213] = 256'hd4efb8f270f535f787f73cf770f6b7f50ff510f4cbf2fcf0d0ee5aed8eecccec;
    decBuf[8214] = 256'he5ede4ee6fef45ef85ee91ed74ec01ec6aec08ed44ee13f048f1d1f26af398f3;
    decBuf[8215] = 256'h6ef3aef274f1f9ef2eee87eb0ee972e792e65ee70ee9e8ebd9ede9ee3bef5bee;
    decBuf[8216] = 256'h9feeddeef5eff4f023f1a4f0feee05ed29eb79e9d0e837e8ace7d6e7fde7f1e8;
    decBuf[8217] = 256'h4dea91eb0ded0cee97ee15efa2ee39ee9bedd2ece7eb49ebb9ea6bea53ea12ea;
    decBuf[8218] = 256'hd7e97ee94de95ce99fe9c3e9e4e9eee9d3e9ebe95cea50ebcfec34eebfee41ee;
    decBuf[8219] = 256'h81ed47ec20eb14ea20e981e8f2e76fe728e769e719e81fe958ea7feb8cec80ed;
    decBuf[8220] = 256'hdfed35ee4fee08ee1aed3decc7ea62e97ae8a8e734e757e7b6e746e831e9cfe9;
    decBuf[8221] = 256'h98ea84eb22ec24ed19ee35efa8efcbef2deff1ed76ec11eb6fe9e6e781e6f6e5;
    decBuf[8222] = 256'hcce5d9e658e889ea2aedefee8af06af1aef170f1c8f0c9efcbed67eb27e9b1e7;
    decBuf[8223] = 256'he5e623e7ace8ddeae8ecc4ee7eef96f02ff101f1d7f064f0b5efd8ee0feeefec;
    decBuf[8224] = 256'he3ebeeea11eaf4e977ea7cebfcec61eeeceebfef32f09af0b7f110f3f8f3cbf4;
    decBuf[8225] = 256'ha4f4b0f315f21cf0b8ed78ebd8e8c8e7d1e6b2e716ea9eede9f0c2f459f7c2f8;
    decBuf[8226] = 256'h30f9ccf872f8d6f6cbf4eff248f083eee8ec72eb2eebe8eb70ed3befecf075f2;
    decBuf[8227] = 256'h74f3fff3d5f3aef3d1f36ff472f5acf67ef7a5f782f765f659f51ff4a4f2a5f1;
    decBuf[8228] = 256'h1af19bf0c2f0b6f112f310f564f698f760f7c7f6dff50df5e6f4c4f422f579f5;
    decBuf[8229] = 256'h5ff576f561f574f586f5f8f57df641f7f8f79ef8dff8a4f84bf8d9f7cbf70df8;
    decBuf[8230] = 256'hc3f8e3f956fa79fadbf9d8f89ef723f624f5dff361f33af3e9f3c3f5aff868fb;
    decBuf[8231] = 256'h96feba00e4018a01eeffe3fd7ffb3ff99ff6daf4e3f399f3ddf396f48ff6f3f8;
    decBuf[8232] = 256'hd7fb90fe0901a502ef02ab0277017dff29fe70fdc8fc2ffceafa6ff9a4f76ff6;
    decBuf[8233] = 256'hc7f5faf59bf724f955fb60fd3cff68017303c7048105d8040d036600edfdadfb;
    decBuf[8234] = 256'h37fa7bfa34fbbdfc22fe0affddffb6ff4effb0fe20fe06fedbfe18003f014b02;
    decBuf[8235] = 256'hb4025502c5010e016800d1ff6fffcefe62fe27fe5cfe30ff6c00e7014c033404;
    decBuf[8236] = 256'hb2042505480529055f040c036a0171ff1dfe64fd9cfd01ffff00db0207057d06;
    decBuf[8237] = 256'hc106fe0637079e066f06f1057e051505f803ec02b201df006c00d500b201b502;
    decBuf[8238] = 256'ha90347046404b20429051706730714092d0a2c0bb70b390bc50a8c09bc070c06;
    decBuf[8239] = 256'ha30307022701e3001802110475061008f008bc09fa09c209290957098209f509;
    decBuf[8240] = 256'ha30a410bd10beb0bd30be50ac9096f08ce0645054604bb03e503f204b706e308;
    decBuf[8241] = 256'h840bfd0d3d10b3117f12bc128412eb114a10510eed0b090917075305b7036d03;
    decBuf[8242] = 256'h29035d047605a707480a760d75102d13f214e8153316ef15ba14321367113b0f;
    decBuf[8243] = 256'h9a0cd60a3a09c507f9063607df074409420ba60de60ff111451383134a13b112;
    decBuf[8244] = 256'h2612a811e8107f10e10f520f030fbc0e7b0eb60e330fa50f65101b1192112a12;
    decBuf[8245] = 256'h3d1208129611f4105c1049107e10af10be107b10dd0f1b0fcc0e130f5810b312;
    decBuf[8246] = 256'hf21493175819aa195f1993186716c7134d11690e770cb30abc099c0af00b1c0e;
    decBuf[8247] = 256'hbd103613761581175d19921aca1a971aaf193418031663139e110310230fdf0e;
    decBuf[8248] = 256'h1c0f35109a11821200137313dc13fc138b144215e815ab162e1745175b172017;
    decBuf[8249] = 256'hc71655167815dd1354128910540fac0e790e040f2b1037117112ec13b7156817;
    decBuf[8250] = 256'hd1196c1b4c1c081c581aef170b155212d90f3d0ec80c840cc10c6a0dcf0e7010;
    decBuf[8251] = 256'h69124514f515ef17bb1874193c19a3180117781547133c11600fb00d970c640c;
    decBuf[8252] = 256'h4c0d1c0f4711bd12991452158a155715cc144e142814bf13e212df11eb10ce0f;
    decBuf[8253] = 256'h5b0f380fd60f9f105611cd11e3118111e0104810bf0f420f110f200f7d0f3310;
    decBuf[8254] = 256'h1e11bd114c1232122d11f30f240e730c5b0b280bb30b820d330f2c1180123913;
    decBuf[8255] = 256'h011368128011ad10ed0ff90edd0dd00c500b510ac6099c090f0abe0a9b0b640c;
    decBuf[8256] = 256'h1b0d920dd30d0e0efc0dab0d260d850cee0b8b0b7a0b8a0b0f0c8c0cdd0cec0c;
    decBuf[8257] = 256'hc40c3e0cc10b0e0b390aa9092609af086f085b08b4088809510a080b7e0b690b;
    decBuf[8258] = 256'h910a5509da0775068d050e05e8040b05a905ac062b08f6092b0b440c770c8f0b;
    decBuf[8259] = 256'h680a75082107ec05d404a1042c055605c905ec05cc053d05ee04a7046604a104;
    decBuf[8260] = 256'h1e059005f7051f061306c60530056d04b7031003790265029b020d0374039c03;
    decBuf[8261] = 256'h78032b03d1027c029d02f702ad036404da041b0508058a04f803480372026f01;
    decBuf[8262] = 256'h7b001fffdafdb4fc40fc1efcfbfcaafe5a005402a80361042904f6030e033b02;
    decBuf[8263] = 256'h2f013a005dff5afe66fdc8fc38fceafba3fbb8fb1afc74fc27fd2cfeabff1001;
    decBuf[8264] = 256'h550228034e03a0024401a2ffa9fd55fc21fb08fad5f94af9cbf858f87bf8daf8;
    decBuf[8265] = 256'hddf95cfbc1fca9fd28feb5fd4cfd6ffcdffb90fb49fb34fb20fb0efb3ffb6bfb;
    decBuf[8266] = 256'hc9fb05fc10fccafb41fb6afaa0f9e9f873f8dbf7a0f747f7f6f6e7f6daf616f7;
    decBuf[8267] = 256'h79f7d7f75cf8fdf869f97df98ff93ef9b9f818f881f71ef7e9f6d9f605f748f7;
    decBuf[8268] = 256'h9df7eaf744f868f831f89bf7adf6d0f506f584f4cbf462f5ecf569f679f612f6;
    decBuf[8269] = 256'h9af507f5a5f470f45ff451f428f4ecf3b5f383f39ef3c7f329f4a1f4d2f4e1f4;
    decBuf[8270] = 256'heef4caf4a9f49ff483f48cf493f4a8f4c7f410f52ef501f585f479f339f19eef;
    decBuf[8271] = 256'h28ee5ced15ee9eefcff1daf3b6f570f6c7f5c8f484f309f20af1dbf05af1cdf1;
    decBuf[8272] = 256'h35f294f277f2f5f11ff11cf028ef4beebbeda1ede8edabeefeefa0f129f38ef4;
    decBuf[8273] = 256'h76f5a0f579f585f469f30ff2cbf04fefeaed03ed30ecbdeb25ecc4ecc6edbaee;
    decBuf[8274] = 256'h98ef61f0aff068f027f0c5ef6cef5cefc3ef56f007f1adf1eef101f2ccf119f1;
    decBuf[8275] = 256'h43f040ef4ceeaeed1eed9cece3ec7aed2bee60ef87f047f169f189f133f17cf0;
    decBuf[8276] = 256'ha6ef6aee97ed8becdcebbdeb4cec03ed38ee5fef1ff042f022f0ccef15efceee;
    decBuf[8277] = 256'hb8eef3ee70ef02f0b3f059f1f1f153f241f28ef159f0deee79ed35ecb6ebddeb;
    decBuf[8278] = 256'h8beca8edb4ee63efc1efdeeff8ef10f07cf0def05bf16cf122f18ff0b7efeeee;
    decBuf[8279] = 256'h6bee83eeefeec7ef90f013f15af144f109f1d4f0a3f094f087f04af0fdefcbef;
    decBuf[8280] = 256'hb0ef0bf0c1f0acf189f219f333f3ecf280f2f6f1c1f190f146f1cef03bf08bef;
    decBuf[8281] = 256'h14effeee39efdaefc8f0a5f16ff2f1f209f31ff381f3daf38df433f59ff5b3f5;
    decBuf[8282] = 256'h5af5a7f401f494f332f320f310f301f30ff34bf36cf3c6f31bf43cf41ef4ccf3;
    decBuf[8283] = 256'h27f3b0f244f231f28af23df3e3f3d1f46ff538f6bbf602f718f704f7cff69ef6;
    decBuf[8284] = 256'h8ff6b7f63df725f802f9ccf94efa07fa19f9bdf71cf693f494f3acf282f2f5f2;
    decBuf[8285] = 256'ha3f3fff4a1f60af94afbc0fc8cfdd2fc49fb18f978f6b3f461f4acf400f62bf8;
    decBuf[8286] = 256'h37fa13fc3efe1fffebff280080ff1bfe7afc81faa5f8f4f64cf67ff60af731f8;
    decBuf[8287] = 256'h8af9cffaa2fb15fc38fc96fc60fd4bfe28ff7eff99ffc3fe87fd60fca0fb7dfb;
    decBuf[8288] = 256'h9dfb2cfc7bfc92fca8fce3fc84fd72fe8eff9b000401e4005400d2ff5bff70ff;
    decBuf[8289] = 256'hd3ff97001a0191017b01f20009002cff63fee0fdf8fd39fe9bfed0fee1fe0dff;
    decBuf[8290] = 256'ha0ffc60041020c044105790546055e048c03cc02a9028902fa0143016d00ddff;
    decBuf[8291] = 256'h2c00600130035c05d106250863084a074b06aa042103220297016d01e0014902;
    decBuf[8292] = 256'ha8023703ba0390041f05d6051e065e064b065d068d06f5066d07be07cd078a07;
    decBuf[8293] = 256'hed06800646069f061107d00753086b082a08ef07960765073907f60689062106;
    decBuf[8294] = 256'ha9057805c20570067507af088209f509180af809db09c109080a1e0a320afc09;
    decBuf[8295] = 256'h6a09e008870897083a09270a050b5b0b410b9b0a030a7a098c09dd09440a870a;
    decBuf[8296] = 256'h630a000a87093609270985090a0a640ad60a3d0bb50b680c3e0d070e550edf0d;
    decBuf[8297] = 256'h9a0cf90a0009ac076e0716081509b70acf0b680cf30c1e0df70c1a0d790d960d;
    decBuf[8298] = 256'he40dcc0d8b0d020d850cd20b5b0bc40a620a2c0a1c0a830a4c0b4f0c430de10d;
    decBuf[8299] = 256'hfe0d7b0dd50c690c2e0c870cf90c250dfd0c470c5c0b7f0ab509d009460a5f0b;
    decBuf[8300] = 256'h6c0ca60dcd0e400fa90fc80f720f240f7d0e8f0df10c280ca50b2f0bee0ada0a;
    decBuf[8301] = 256'hec0adc0ab00abd0ae10a180b860bee0b300c3d0c1c0cd60bdf0b180c7a0c0d0d;
    decBuf[8302] = 256'h960df00d620e8e0eb60ef30ee80e8e0ef00dd70cca0b900a6909aa088708e608;
    decBuf[8303] = 256'h7509950aa10b500caf0c920c430cfc0bbb0b800b920b820b910b9e0baa0be10b;
    decBuf[8304] = 256'h3b0ca80c100d380d130d840cd40bcf0ada09be08fe07db07fb07fd08370ab20b;
    decBuf[8305] = 256'h170dff0d290e030e9a0dbd0cf40bd40a7b093608bb062206f4057206cc076d09;
    decBuf[8306] = 256'h860a1f0b4d0b230bb00a8d0aad0a030b1d0b350b1f0be40aaf0a7e0a520ad909;
    decBuf[8307] = 256'h47096f08a60723070b072107aa074b08e3086c09c509d609e409d709cb09aa09;
    decBuf[8308] = 256'h7809ef083e083907450668054b0565053b0677074a085609bf09df09fb09ad09;
    decBuf[8309] = 256'h07094408c1077a07900740081609a6098c0987084d07d205d304470472049804;
    decBuf[8310] = 256'h01055f05430591050806ca06b607d208450922098408820748067505b5049204;
    decBuf[8311] = 256'h7304020585055b065e075208f008d30850081c07a1053c04f70224024b02f902;
    decBuf[8312] = 256'h970360047b0463044d046104de04d205c606a307c0073d079706a9050b05ee04;
    decBuf[8313] = 256'hd4045d0470035302fa001200e8fff4007402d9031d05f00563068606e5063b07;
    decBuf[8314] = 256'h8a07420754067a0416027b0070fe2cfe69fe82ffe7002c02fe027103da03fa03;
    decBuf[8315] = 256'h160430044804070457038102f101d7011e02b60218032a03970298015e008cff;
    decBuf[8316] = 256'h65ff88ff26007d00ff00170183010d02d1028803ff03e903ea026a010500c1fe;
    decBuf[8317] = 256'heefdc8fdebfd0afe27fe41fe88fef5feccffcf0009028702ae02450268016500;
    decBuf[8318] = 256'h71ffd3fe7dfe97feaefe99fe5efe28fef8fdcbfdd9fdcdfd96fd3cfdcefc85fc;
    decBuf[8319] = 256'h92fcfffcdcfdbafebdff6b00ca00ad005f00e8ff25ff06fef9fc7afb7bfa93f9;
    decBuf[8320] = 256'h14f93bf9e9f9c7fac9fbbdfc9bfd64feb2fecafe89fed9fdd3fc9afbc7fa07fa;
    decBuf[8321] = 256'h9ef9bef914fafffaddfb6dfc23fd3bfdfafc71fcf4fb62fbd8fa5bfae9f965f9;
    decBuf[8322] = 256'h0bf9baf8c9f8d6f8faf805f9bff849f8d7f7abf7d3f789f8a8f9b5faeffbc1fc;
    decBuf[8323] = 256'h81fda4fd45fdb5fccafb6efa2af903f8aaf665f53ef47ef35bf3f9f3fcf47cf6;
    decBuf[8324] = 256'h47f8f7f910fba9fbd7fb59fb99faa5f949f804f789f58af4a2f378f3ebf325f5;
    decBuf[8325] = 256'hf4f6a5f82efa93fb1efc48fc88fb4efad3f86ef770f594f35ff2b7f184f10ff2;
    decBuf[8326] = 256'he1f288f410f60ff7f7f776f89cf879f8dbf785f702f7eaf6d5f610f722f752f7;
    decBuf[8327] = 256'h61f71ef7c9f650f67df5b4f4fdf357f316f378f319f407f5e4f5adf664f7abf7;
    decBuf[8328] = 256'h96f782f74df7dbf639f6a1f518f5bef4aef4f8f48bf53cf6b2f6c8f6b4f614f6;
    decBuf[8329] = 256'h7cf5f3f476f445f454f47cf4d1f476f51cf6dff661f7a8f768f705f765f6f8f5;
    decBuf[8330] = 256'he5f5d3f5e3f5f2f5aff572f567f585f5eaf57df606f760f74ff7cbf64ef6bbf5;
    decBuf[8331] = 256'h59f524f534f560f5bef513f676f6eef680f70af887f8b7f86ef8dbf703f700f6;
    decBuf[8332] = 256'h52f532f54ff506f6dbf6def78cf8ebf842f95cf973f907f9a5f8bdf7a0f694f5;
    decBuf[8333] = 256'h9ff401f41ef4d5f40af631f78af8cff9a1fa61fbcafbaafb54fb9dfac7f9fef8;
    decBuf[8334] = 256'h47f8a1f760f7fef6ecf6fcf646f7d9f7b1f8b4f962fac1faa4fa56fab0f943f9;
    decBuf[8335] = 256'he1f8cff800f985f926fabdfa6efbe5fbcffb94fbf3fa31fa7af9d3f8bef8f9f8;
    decBuf[8336] = 256'h76f96afa5efb7afc3afda3fd83fdbafc66fb22fafbf8d4f8f7f8d5f911fb38fc;
    decBuf[8337] = 256'hf8fc60fdbffda2fdbdfd75fd34fdd2fc79fc69fc77fcbafc0ffd88fdb9fdaafd;
    decBuf[8338] = 256'h32fd5ffc5cfb68fa09fa26fadcfae2fb1cfd42fe9cff84000201750198013901;
    decBuf[8339] = 256'ha900beffa2fe95fd5bfc89fbc9faecfa0bfbd4fbf4fc00fe3aff610021018a01;
    decBuf[8340] = 256'h6a014d01ff005900c1ff38ffdffe8dfe7ffe8cfeb0fed1fedbfed2fecafee0fe;
    decBuf[8341] = 256'h3affd7ff9a005101c801dd01a2014901d700700012008dffecfe80fe1efee8fd;
    decBuf[8342] = 256'h3afedcfecaffe600f301a1023f035c034203cb025f02af013801cc004200c5ff;
    decBuf[8343] = 256'h33ffaafe98fea8fe2dffceff6500ee0048017801a501cd0109025602b002ed02;
    decBuf[8344] = 256'h240342032703dc026e02cc010a018700e1ffa0ff65ff53ff22ff14ff21ff8eff;
    decBuf[8345] = 256'h6b008801e1022604a404cb04620485034802220162006eff0fff2bff7aff5000;
    decBuf[8346] = 256'h520146022403b403ce0386031a039102f00184012201ec009b005100f4ff9fff;
    decBuf[8347] = 256'h52ff34ff74ffefffb4006b0141020a0358039f03b503c903fe032f043e04fb03;
    decBuf[8348] = 256'h4503f101500037ffd2fd47fd71fde5fd93feb0ff0901f1011803d8038604a604;
    decBuf[8349] = 256'h8904d203fc02f90105012800d2ffecff6300fa00830100025202430236021102;
    decBuf[8350] = 256'hda0194014201f50087003d0015003a009d003001b90136026702760283025f02;
    decBuf[8351] = 256'h6a02600244020b02a9014b0127014801a2010f02760284024702e4016c01da00;
    decBuf[8352] = 256'h77001e00edffdfffecff2900b80068013e020703f203900420050605bf04fc03;
    decBuf[8353] = 256'ha9020701efff8afe5bfe31fef1fee5ff02010e020203a103f7031104ca033203;
    decBuf[8354] = 256'ha902080271010f01fd000d0139019701ec01230255025e0256023f0238023e02;
    decBuf[8355] = 256'h66029402c002d102ad026702f90192014f017401c1011b026f02900286025902;
    decBuf[8356] = 256'h510258028802c002f5020a0310032c036f03c103f803ee03650366022c015900;
    decBuf[8357] = 256'he6ff4f002c0168028f0302046b044b04f503db03c303d903ec03fe03ce03a103;
    decBuf[8358] = 256'h790355037603a803c303bb037703130380021e020c023d02c10262032504a804;
    decBuf[8359] = 256'h1e055f05730585055405ed045a04a903d30243022902a00263034e046a052a06;
    decBuf[8360] = 256'hd906f8061507fb068406c205a20496035c02890116013901d701da025904be05;
    decBuf[8361] = 256'h6007780877094909cb08be073e06d904f10373034d037003ce0398044f05c505;
    decBuf[8362] = 256'h5d0670065e064e060406dc05a0057f0561056a058305d5056406ed066b07bc07;
    decBuf[8363] = 256'had076a07fd065b06ef05650530051f054c057405e1054806c10632077c07a407;
    decBuf[8364] = 256'hb0077907e3064c069b0525050f0571051206d5068b070208430857082108d007;
    decBuf[8365] = 256'h2e076b06b4053d05fc045f052306da06b00740082508af07ec0635068f054e05;
    decBuf[8366] = 256'h6205df055106d5065207a407b207a50781074a071807d8068e062006b8055b05;
    decBuf[8367] = 256'h4f058605f4057806d206e206b60673064e066f06b506f506fe06ba064306d205;
    decBuf[8368] = 256'h6a055d0569055e052c05ec04a2048404c4044005e10578062907700785072307;
    decBuf[8369] = 256'ha606f3051e058e040b04f403de03f203e003f0031c047a04ff047c05ee05fd05;
    decBuf[8370] = 256'hba054d05c8046f041d04f103c903bd03c8032204a704240576052c059904c103;
    decBuf[8371] = 256'hf802410229026a02a502fe022f035b03b9032604ab04e004f1048904db030603;
    decBuf[8372] = 256'h7602f301dc01f1017b02f802490358034a030e03ab0268021302f201c0018001;
    decBuf[8373] = 256'h57014f017201cf017d02f40235032103a40212028901530163018f019d01a901;
    decBuf[8374] = 256'h72011801f400e900f3000e0116010001dd00e4000b014301690170013701d600;
    decBuf[8375] = 256'h930056004b0055005f0056002200f2ffd2ffb6ffc6ffe6ff1d00520082008800;
    decBuf[8376] = 256'h6c002900c5ff82ff5eff53ff85ffa0ffb9ffb1ff9dffa3ffbfffd9ffd4ff94ff;
    decBuf[8377] = 256'h0cff5bfeb5fd74fd60fd96fdc7fd10fe53fea8fe21ffb3ff15004b003b00f1ff;
    decBuf[8378] = 256'h5effd5fe7bfe09fea2fd2afdb8fc33fcdafba9fbd5fb33fce9fc3dfe81ff5400;
    decBuf[8379] = 256'hc700ea004c0049ff0ffe3cfd7dfc14fc76fbe6fa63fa4cfab8fab7fbf1fc18fe;
    decBuf[8380] = 256'hd8fe40ffa2fe12fe27fd89fc33fc19fcd1fbbcfba8fbdefb0ffc93fc10fd82fd;
    decBuf[8381] = 256'hccfdbffd6afd07fd8efc1dfcb5fb58fb03fbe2fac4faa8fa90fa88fa9dfafbfa;
    decBuf[8382] = 256'h8efb3efce5fc25fd39fde0fc2dfcb6fb4afb36fb6cfbdefb28fc50fc44fcf7fb;
    decBuf[8383] = 256'h89fb04fb63faccf991f97ff9d0f955fad2fa64fbeefb47fc98fcc4fc9cfc2ffc;
    decBuf[8384] = 256'h6ffb84faa7f951f937f97ef915fa9ffaf8fa6afb96fbbefbcafbbffb8dfb3bfb;
    decBuf[8385] = 256'hc2fa71fa27fa1afa26fa47fa79fab9faf2fa09fb1efb0bfbd8fa7ffa12fac8f9;
    decBuf[8386] = 256'h85f991f9c8f922fa8ffaf7fa54fb91fb9cfb7efb3efbc2fa21fab5f92cf9f6f8;
    decBuf[8387] = 256'he6f830f98df92bfac2fa4cfbc9fbfafbebfba8fb3bfbd4fa5bfae9f982f925f9;
    decBuf[8388] = 256'hd0f8aff8e1f845f9d8f989fa00fb6cfb58fb22fbb1fa67fa24fae7f9c6f9a8f9;
    decBuf[8389] = 256'h7bf962f96af99af9f7f970fae2fa2bfb39fbfcfa99fa3bfacef9a2f9aff9bcf9;
    decBuf[8390] = 256'hddf9e7f9cbf9b2f99cf9bef903fa55faa2fa98fa58faedf986f978f99df9eaf9;
    decBuf[8391] = 256'h44fa68fa73fa2dfa00fad6f9c0f9abf998f97cf96df97bf990f9bbf9e2f9f1f9;
    decBuf[8392] = 256'hf6f9faf906fa25fa43fa47fa36fa2cfa29fa36fa55fa51fa17faacf927f9aaf8;
    decBuf[8393] = 256'h79f8a5f81ef9b0f912fa24fa34faeaf9a8f983f978f982f9d4f937fab0fa21fb;
    decBuf[8394] = 256'h30fb08fb83fabef9d3f835f8dff7f9f740f8d7f861f902fac4fa7bfbf2fb33fc;
    decBuf[8395] = 256'h1ffc5afb6ffa53f946f898f778f795f7e3f789f84cf903fad9faa2fbf0fb08fc;
    decBuf[8396] = 256'h9cfb13fb4efacbf955f93ff953f988f9faf97ffafcfa2dfb3bfbc3fa31fa80f9;
    decBuf[8397] = 256'h09f9c8f8dcf835f9c8f978faeffa5bfb96fba8fb98fb89fb46fb3afb19fbe7fa;
    decBuf[8398] = 256'ha7fa5dfa03fac6f9bbf9edf952faaffaecfa0dfb17fb32fb7cfbeafb52fc95fc;
    decBuf[8399] = 256'ha1fc6afcfcfb77fb1efb0dfb1cfb44fb99fbbafbb0fb95fb6bfb46fb68fbadfb;
    decBuf[8400] = 256'h11fc6ffcacfca1fc5bfc09fcd2fbf0fb2ffc8afcdffc16fd20fd29fd42fd58fd;
    decBuf[8401] = 256'h7bfd75fd2bfdd1fc64fc1bfc28fc7dfc0cfd95fd12fe43fe34fe27feeafdc9fd;
    decBuf[8402] = 256'hbffdc8fdf2fd17fe1efe18fef0fdaefd80fd78fd9dfdf7fd64feaefed6feb1fe;
    decBuf[8403] = 256'h90fe86fea2fefdfe6affd1ff14002000ffffe1ffb3ff8aff47ff07ffbcfe76fe;
    decBuf[8404] = 256'h80fea9fe0aff68ffa5ffb0ffbaffc3ffdbff2e009100ef00430164016e014101;
    decBuf[8405] = 256'he6007900f4ff77ff46ff73ffebff9e007301ca01e401cc018b01290117012701;
    decBuf[8406] = 256'h54019701eb0138027e029a0281022f02a001ef004900b1ff9effd3ff4500e700;
    decBuf[8407] = 256'haa01950272033c04be040605f0043f046a036702b8011a01fe004c01c3012f02;
    decBuf[8408] = 256'hb8023503c803020438040704a003280395023302fe010e025802d0026203ec03;
    decBuf[8409] = 256'h6904ba04e604d904cd04960478044a042104ec0393032603bf027c027002bd02;
    decBuf[8410] = 256'h3f030304ee048d051c066b06b2067106e8056b05b8044104aa036f038103b103;
    decBuf[8411] = 256'hfb0359049504b604e80428056205a605e5050f0616060f06f005df05c605ae05;
    decBuf[8412] = 256'h990576054d053105210538057805ef056006e5063f076f077e0771071c07a306;
    decBuf[8413] = 256'h11066005e904a80495041205a4055506fb066707a207d807c707b907c607ea07;
    decBuf[8414] = 256'hf50713080a08c0073e079d060606a40592050306e106fd07bd086c094c09f608;
    decBuf[8415] = 256'h7308fc0765072a07f406050713073c076007ad07f30721086b089d08b808e108;
    decBuf[8416] = 256'h07090e092d09330919091409ff08e408be087b081708b907640743077507d907;
    decBuf[8417] = 256'h5208c4082b098809dd09400a9e0ac20a8b0af50907096908da07f4076a080209;
    decBuf[8418] = 256'h8b099d096c092309c508700865085b0840085808600867089308dc083609bb09;
    decBuf[8419] = 256'h5c0af30aa40b1b0c050c7c0b930a3709f307cc060c06e90548069e065507fb07;
    decBuf[8420] = 256'he908c709900a470b8e0b780bef0a2a0a3f096208d20750070807f306df06f106;
    decBuf[8421] = 256'h4207c7074408f7089d09340a970acc0a9b0a170a52093308260778061906fc05;
    decBuf[8422] = 256'h16062e069a06fc065607e8074a08a308d408c5086808fb0793076b079007b107;
    decBuf[8423] = 256'hcf07b3075807d3065606e4059a05a805e40531068b06c806ff0631075f076707;
    decBuf[8424] = 256'h5f074b070607b4063b06a9051f05a204510460048804c40427058505f2053c06;
    decBuf[8425] = 256'h9a06d606f706ed06ad0632069105ce041704a003340348035a03ab033004ad04;
    decBuf[8426] = 256'h3f05c90522063206e8053b059404d2034f0308031d03310367039703a603b403;
    decBuf[8427] = 256'ha7039c03920377036f037603b403ee0331044d043404d3035a03c80266025402;
    decBuf[8428] = 256'h64029002b902c502ba029c028002570232020102d601ba01aa01b801f8014a02;
    decBuf[8429] = 256'had020b0347035203480308039d02fb0138018100dbff6fff83ffb8ff2a009100;
    decBuf[8430] = 256'hd400f800030121013d0166018c01bc01e7011a023c024302ee01510138002bff;
    decBuf[8431] = 256'hf1fd1efdabfccefc2dfdf6fd16ff22001601f40184029e0227023901ddff99fe;
    decBuf[8432] = 256'h72fd65fcfcfbddfbfafb7cfc22fde5fd04ff1100bf001e0102014b0045ff51fe;
    decBuf[8433] = 256'h35fd28fc7afb1bfb38fb52fb99fb30fcbafc13fd64fdaefdbbfdaffd8efd20fd;
    decBuf[8434] = 256'h9cfc1efccdfba1fbc9fbedfb0efc04fcb2fb23fb9afa64fa54fabbfa34fba5fb;
    decBuf[8435] = 256'heffbfdfbc0fb9ffb81fb66fb4dfbfafa6bfabbf9e5f855f83bf823f88ff8f2f8;
    decBuf[8436] = 256'h4bf9bdf924fa67fabcfaf3fa11fb08fbdefa6efabbf9e5f81cf831f793f676f6;
    decBuf[8437] = 256'hc4f66bf784f890f93ffa5efa42fabff919f981f8d1f75af7eef68cf656f687f6;
    decBuf[8438] = 256'heef681f732f8a9f8bef85cf898f7acf6cff5b2f5ccf5a2f6def705f912fa7bfa;
    decBuf[8439] = 256'h9afa0afa1ff903f8a9f665f592f4d2f36af389f3dff396f4cbf5f2f64bf833f9;
    decBuf[8440] = 256'h5df937f989f8eaf75bf70cf7c5f6dbf6a0f646f6f5f5c9f5d6f55cf6d9f66bf7;
    decBuf[8441] = 256'h7ff725f773f69df59af431f451f4a7f492f5aff608f8f0f8c3f936fa59fabbf9;
    decBuf[8442] = 256'h7ff858f7b2f599f434f3a9f27ff2a5f20ef3ebf327f5a2f607f84cf9c7fac6fb;
    decBuf[8443] = 256'h51fc27fc1bfb9bf96af7c9f405f369f189f0cdf002f28bf356f506f7fff853fa;
    decBuf[8444] = 256'h88fbc0fb8dfb02fbdbf982f83df716f60af55bf4fcf319f4d0f4a6f56ff6f2f6;
    decBuf[8445] = 256'h39f723f7c1f668f657f6bff687f78af8c4f942fab5fa93fab5f9ecf801f823f7;
    decBuf[8446] = 256'h5af60cf6c5f505f668f6e5f677f7d9f7ebf79af750f70df701f764f7f7f780f8;
    decBuf[8447] = 256'h21f962f94ff93df92cf91ef946f96af949f917f98ef8b6f7edf602f6a3f5c0f5;
    decBuf[8448] = 256'h77f67cf7fcf861faa5fbccfcf3fc8afcecfbb0fa89f92ff8ebf6c4f551f52ef5;
    decBuf[8449] = 256'h8df58ff60ff8daf98afba3fca2fd2dfeaffda2fc22fb57f9a7f71ef6ebf576f6;
    decBuf[8450] = 256'hf2f723fa2efc82fd3bfe03fe6afd25fcfefaf2f943f9a5f8c2f8a8f81ff9b6f9;
    decBuf[8451] = 256'h67fa3cfb06fcbdfc63fdcffd0afed4fd21fd1cfce2fa67f9cef843f8c1f8cef9;
    decBuf[8452] = 256'h4efbb3fc54feddff76000101830076fff6fd2bfc7bfa63f9caf8f8f8cbf924fb;
    decBuf[8453] = 256'hc5fc4efeb3fff80076019d01ee0092fff1fd68fc9dfa68f930f9c9f90efb31fd;
    decBuf[8454] = 256'h3dff9100c5016e023b02b001dd001d006fffd1fe41febefde9fc59fcd6fb1dfc;
    decBuf[8455] = 256'he0fc68fef1ffbc0175021d038402f90127011a0026ff88fe32fee3fdfbfd67fe;
    decBuf[8456] = 256'h18ffedffb7006e01e401500264022e02dd013b01a400f3ffacff96ffaaff0300;
    decBuf[8457] = 256'h54009e0016018801ef0183020c03650376034903d102fe01fb000700eafe2afe;
    decBuf[8458] = 256'h07fe66fe30ffb70040020b04bc05d40607071f06f8040603a20006ff91fd4dfd;
    decBuf[8459] = 256'h81fe0a00d5010a032304bc048d046304f003cd03ad03ca03b003980301035002;
    decBuf[8460] = 256'h7b01b1009700af0072012802fe028e03dc032404390426041404c2033e037902;
    decBuf[8461] = 256'hc2014b013601bf01a8024304cc05cb0656072c076c06ec042103ec016300caff;
    decBuf[8462] = 256'h9cff6f007b01fb026004a505cb063f071c073e060205870322023a0110018301;
    decBuf[8463] = 256'h770255035704c0041f0502051c05d504bf0484044f043f0430047304af04fc04;
    decBuf[8464] = 256'h2e054a0531050b05c0046604f90391034f034203a5033904c204d4046204a203;
    decBuf[8465] = 256'heb02d4026b039104610696073e080b082307a805a904c1039703bd03e0033f04;
    decBuf[8466] = 256'h22040804c1038003940335044e05a706ec07be083109c908eb07af0634056903;
    decBuf[8467] = 256'h3d01c8ff74fe36fe4eff4b022506c4091e0c670d3c0c780a9407db041703c402;
    decBuf[8468] = 256'he4012802ea01b2014b02330302052e073909050a430a2b09fa06ee0412035902;
    decBuf[8469] = 256'h91029003d504a705ce056505880485031c037b03f104bc06e808c8090c0ad708;
    decBuf[8470] = 256'h4e07b704f30258017700bb00f0017903aa05b50791094b0a830aea09a5082a07;
    decBuf[8471] = 256'hf904ee029a0165009d009c013d03c604c50550067b0654063106cf0699078408;
    decBuf[8472] = 256'h2209cc087807d705de030202480110010f02f7021e04de04d20570060007b707;
    decBuf[8473] = 256'h5d08c908b508f1076906e00415035c0294022d031504e7040e05a5040704ea03;
    decBuf[8474] = 256'h39043e05be06bd07a4087a086e073406640430031702e4011202390346048005;
    decBuf[8475] = 256'h520679061006b1052205d304bb04d104bd04cf042105e005cb06a907ff074807;
    decBuf[8476] = 256'he405b303a801ccff8eff36000102b203ab05ff06b807f007bd07d5060306a904;
    decBuf[8477] = 256'h65039202d201f5019302cf034a05490631070707fb057b0416032e0258026503;
    decBuf[8478] = 256'he404e30512063f05990380028101b0012e02ee02570337031a03000377033a04;
    decBuf[8479] = 256'h2505c305e0059105eb0454041904e303d303a7032e037b02050299018501bb01;
    decBuf[8480] = 256'h4d02fd02a403e503f803c303b203df0321048f04d8049504e0038c0247012000;
    decBuf[8481] = 256'h61ff83ffe2ffac00ff01a10329058e06d307a9079c0691045b0137ff46fda0fd;
    decBuf[8482] = 256'h3cffb1008d02c203fa03c7033c0366038d03b0039003c70273012e005cff35ff;
    decBuf[8483] = 256'h6f00ea01b503ea04220523048202f900faffccfff6ff69008c006c0016003000;
    decBuf[8484] = 256'ha700eb013003ab04de0453042c0386016d00d4ff0300d50048016b01cd00caff;
    decBuf[8485] = 256'hd6fe38fe55fe74ff1a01a3026e042705600561041c03a101d6ff26fe7dfde4fc;
    decBuf[8486] = 256'h6ffd42fe4fff43005f01d2013b021b02ff01e501fc0112024d021702a501e600;
    decBuf[8487] = 256'hfbff1dffc7feadfe24ffbbff6c00e20023011001da006800c6ff2ffff4fe06ff;
    decBuf[8488] = 256'h57ff1700cd007401e001f3015301650009ff21fe4efd28fd91fdadfe07004b01;
    decBuf[8489] = 256'hca013d021a02bb0165011601cf006300daff15ff2afe4cfdbdfc6efc86fcc7fc;
    decBuf[8490] = 256'h78fd4dfeddfe94ffdbff1c005700d40087012d026e0233024b01efff4dfec5fc;
    decBuf[8491] = 256'hc6fb97fbc1fb34fce3fc42fdd1fd88fe2fffc6ff7700ed000301c800270039ff;
    decBuf[8492] = 256'h1dfe10fd62fc03fc59fcdcfc82fd45fec7fedffe9efe3cfe9bfd2ffdf4fc2afd;
    decBuf[8493] = 256'h9bfd5bfe46ffa5ffc2ff3fff6afea0fde9fc73fc88fc9cfcaefc7dfcdbfb18fb;
    decBuf[8494] = 256'h96faadfa9bfb36fda0ffdf0155039903e002e70083fe43fca2f9def78cf741f7;
    decBuf[8495] = 256'h85f73ef8c7f9f8fb03fe57ff8c00c4002b00e6fe14fea1fdc4fd62feb8fe35fe;
    decBuf[8496] = 256'hd1fca0fa95f841f77ff797f862fa12fc0cfed8fe91ffc9ff96ff0bff38fe78fd;
    decBuf[8497] = 256'h84fce6fb56fb08fbf0fadbfac7fab5faa5fad1fa14fb81fb23fcbbfc44fd7afd;
    decBuf[8498] = 256'h69fde5fc44fcd8fbc4fb1dfc11fd05fe64fe47fe91fd2cfc61fa2df984f851f8;
    decBuf[8499] = 256'hdcf8aff9bcfa3bfca0fd42ffeaffb7ff72fe4ffcaef9e9f797f7e2f746fa86fc;
    decBuf[8500] = 256'h91fe5dffa4feabfc47faabf8cbf797f8c3fa64fd28ff7affc5ff71fe3cfdb3fb;
    decBuf[8501] = 256'hb4facdf94ef9dbf844f921fa24fb18fcb6fc60fc75fb58fa98f9bbf998fa0efc;
    decBuf[8502] = 256'h73fd5bfe85fec5fd8bfc10fbabf9c3f899f80cf9bbf998fa61fbe4fb8afcf6fc;
    decBuf[8503] = 256'h80fdd9fdc9fd62fd99fc5dfb36fa76f9c8f8a8f8fef8b5f95bfa49fb27fc29fd;
    decBuf[8504] = 256'hd8fd37fee0fdc1fc1bfb92f92df8fff7d1f82bfa6ffb96fcbdfc54fcb6fb26fb;
    decBuf[8505] = 256'hd8faeffa5cfb6ffb3afba7facff9cdf864f8c3f88cf914fb0dfde9fea2ffdbff;
    decBuf[8506] = 256'h42ffa0fd37fbf7f881f72df674f5acf545f68af759f985fb90fd6cff2500ce00;
    decBuf[8507] = 256'hcfff8afebbfc8ffa19f9c5f788f7c0f759f841f913fad3fa3cfb9bfbf1fb73fc;
    decBuf[8508] = 256'heafc56fd6afdc9fcdbfbbffa65f97df8fff7d9f787f864f914fbc4fcbdfe1100;
    decBuf[8509] = 256'h4f0036ff6bfdc4fa95f772f547f457f5f2f693f9c1fcc0ffea00fa0103018dff;
    decBuf[8510] = 256'h39fe0efc98faccf913f9daf8a7f879f8f7f86bf95ffa7bfb88fc08fe07ffeeff;
    decBuf[8511] = 256'h1900f2ffb8fe3dfd0cfb01f9adf7f4f62cf791f832fabbfb20fdabfd2afe9dfe;
    decBuf[8512] = 256'h05ffa3ff33004d00d7ff92fef1fc68fb03fa1bf945f9b8f9f2fa19fcd9fccdfd;
    decBuf[8513] = 256'h2cfe82fe68fef1fd85fdfcfca2fc72fc80fcdefc4bfdd0fd4dfe7efe8dfe64fe;
    decBuf[8514] = 256'h71fe7cfeaefec9feb0fe4ffea1fdfbfcbafcf5fcb9fda4fe42ff5fffddfed7fd;
    decBuf[8515] = 256'h29fdcafc5afd45fe62ff21008a002b009bff19ffa2fe8cfe79fe67fef5fd53fd;
    decBuf[8516] = 256'he7fcacfc29fdfcfd39ff5f00d300f50097000700b8ffa1ff0d0048007d006d00;
    decBuf[8517] = 256'h4100fefff2ff29008300bf007200dcffc3fe03fe9bfdfafdfcfe7c007b016302;
    decBuf[8518] = 256'h3902c601d2003300ddff2c00d2006901f3010402d401140129000cff00fe0bfd;
    decBuf[8519] = 256'hecfc7cfd03ff6d01ad034d065d07af07cf066b042b028affc6fd2bfce0fb9cfb;
    decBuf[8520] = 256'h55fcfdfcfcfdfbff5f0243053407f908a708c607620523031701c3ff86ff4dff;
    decBuf[8521] = 256'h80ff52ff28ff4effb7ffd4002d027203ed048605b4053605c304140437033402;
    decBuf[8522] = 256'hfa00d3ff13fff1feceff4401a9024a046305960567054004e702a201270028ff;
    decBuf[8523] = 256'h9dfe1cff2800a801730323053c063b07c607f0077d078906ee0465039a016500;
    decBuf[8524] = 256'h4cff19ff48ff1a00740115039e0403064807c607a007f1061406d804b103f102;
    decBuf[8525] = 256'h4202e4018d013f0127016801ca018f024603ec03830434050a060c0701089f08;
    decBuf[8526] = 256'h4808290783051a037e019e005a0013012c0291037904a3041605f30413053005;
    decBuf[8527] = 256'he104c9045d044a045c04ee04c605c806bd075b0804084e07e9058404e302ca01;
    decBuf[8528] = 256'h3101030181018e020e04730514072d08c60851092709b3080508e8062906ef04;
    decBuf[8529] = 256'h1c045c03f4025502c60143015b01c701ed02bd046d06f607f50880095609e308;
    decBuf[8530] = 256'h3408960793065a05de03df0254027e02d8037905020701082f08050845079706;
    decBuf[8531] = 256'hf90569051b05d404be04aa040405d7051307e607a608c908eb07af0634053504;
    decBuf[8532] = 256'haa03d40347043b05d905f605dc0595057f050806f1068f07e50762072e06b304;
    decBuf[8533] = 256'hb4032803fb03540599061707f1068806ab051b053505ac056f06bd06d5066906;
    decBuf[8534] = 256'h2e061c064d069706d906b50610060b051704b80348049b053d073609020ac409;
    decBuf[8535] = 256'h3b087006c004a7030e0399036c042c0520067f06d50623076b072a07c806df05;
    decBuf[8536] = 256'hc3040304540335038b030e048404c50427055d058e05ba05c705bb05b005ba05;
    decBuf[8537] = 256'h0c069b06fe063307c106e405c804bb03520372033b048f05d306fa076d08bf07;
    decBuf[8538] = 256'he2066c0507047c03520378039b03bb039e03b8032f044805a10643087b084808;
    decBuf[8539] = 256'ha6063d04a202c10105023a03e3037c044d04cf03a803cb0369046c0560068006;
    decBuf[8540] = 256'h2a0673059d049a03ec028d027002bf023503f8037b04f1043205460558056805;
    decBuf[8541] = 256'h3c05c304d003dc02bf014c01b401d1022a046f05ed05c7055e05c0046a041c04;
    decBuf[8542] = 256'hd40394033103b40243021602ee01fa010502fb0104020d025002b5022d039f03;
    decBuf[8543] = 256'hcb03d8039c03230370029a019700a3ff44ff28ffaaffdf0006025f03ea031504;
    decBuf[8544] = 256'hee0386032703d002b6029f0232025b0158001eff4bfe25fed3fe2f002d028103;
    decBuf[8545] = 256'hb6047e04e503a00279016d004a006a008600d5008d00cbff14ff3efeaefd94fd;
    decBuf[8546] = 256'h0bfecefeedffad005b017b015e011001990058001d00a0ffedfee8fdf4fc56fc;
    decBuf[8547] = 256'hc6fbe0fb28fc68fcf2fcdafdf7fe9d0026022503b0038902960032fef2fb7dfa;
    decBuf[8548] = 256'h39faf2fa7bfce0fd6bfe95fed5fd6dfd0efd64fd4ffeeaff7301d8020603e001;
    decBuf[8549] = 256'ha0ffbcfc03fa8af7eef5a4f5f8f6a8f811fbf6fde7ffac015901790025fff9fc;
    decBuf[8550] = 256'h84fbb8fa7afa42fa0ffa84f9b1f8f1f788f766f815fabcfc36ff7601c001f400;
    decBuf[8551] = 256'h44ffdbfc9bfa90f8c4f701f83af839f97dfaa4fbb1fca5fd43fe99fe17fe11fd;
    decBuf[8552] = 256'h92fb2dfae8f815f8eff758f8b7f846f995f93bfad2fa83fb59fce8fc03fd8cfc;
    decBuf[8553] = 256'h9efb42fa5af933f873f751f731f74ef768f750f73af79df785f820fa19fcf5fd;
    decBuf[8554] = 256'h2aff62ff63fe65fc01fac1f7b6f5eaf4acf4e4f4e3f5cbf646f8abf9a9fbfdfc;
    decBuf[8555] = 256'h32fe6afe37fe4ffdd4fb6ffa2bf904f891f76ef7cdf723f871f85af8edf764f7;
    decBuf[8556] = 256'he7f6d7f696f7eaf88bfa14fc13fde5fc12fc1ffa43f893f60af571f4a0f472f5;
    decBuf[8557] = 256'hccf610f88bf98afab9fa8ffa82f98ef8b1f721f707f71ef7b6f766f83cf905fa;
    decBuf[8558] = 256'hf1fa4ffba6fb57fbe1fa1efa33f955f88cf7d5f62ff698f55df5b6f5aaf6b5f8;
    decBuf[8559] = 256'hc0fa9cfcd1fd09fe0afd69fb70f91cf8e7f6aff6e2f610f73af761f7f8f699f6;
    decBuf[8560] = 256'h43f691f608f721f87bf9bffa92fbb8fb50fb33fadaf895f717f7f0f659f736f8;
    decBuf[8561] = 256'hfff882f9c9f9b4f92af989f8f2f790f77ef731f836f9b6fa1bfc03fd2dfdbafc;
    decBuf[8562] = 256'hc5fbe8fa1ffa68f921f90bf9d0f877f805f89ef75bf767f7e0f7d4f853fab8fb;
    decBuf[8563] = 256'h5afd72fea5febefd42fc11fa06f82af67af4d2f305f449f519f744f950fba4fc;
    decBuf[8564] = 256'hd8fd10fe77fd33fc0cfbb3f9cbf84cf873f8dbf8b9f982fa39fbb0fbf0fb04fc;
    decBuf[8565] = 256'hf2fbc1fbd0fbdefb02fc23fc19fcfefbb3fb45fbc1fa43faf2f91efab2fab1fb;
    decBuf[8566] = 256'hebfc11fed1fef4fe95fe93fd13fc14fbcff9fdf8d6f8b3f812f9a2f98dfa6bfb;
    decBuf[8567] = 256'h6dfc1cfdbafd10fe2afe42fe2cfecafd71fd9efc9bfba7fac9f93af954f929fa;
    decBuf[8568] = 256'h9ffb04fda6febefff1ffc3ff99ffd9feb6fe57fe3afe20fe7afdb7fc00fc5afb;
    decBuf[8569] = 256'h45fb1cfc92fd5dff0d012602f3016801edff88fee6fc3efca5fb77fbf5fb68fc;
    decBuf[8570] = 256'hd1fc6ffdfffdb6fe8bff1b009e00e500cf006d0085ff68fe0ffdcafbf8fa1efb;
    decBuf[8571] = 256'hccfb67fd61ff3d01ed0295036203d7025c01f7ff0fff91fe6afed3fe71ffc7ff;
    decBuf[8572] = 256'hadff66ff25ff39fffdff1d0176025e03dc0303045403b602b301bf00210058ff;
    decBuf[8573] = 256'hd5febefea8fe0aff63fff6ffa6004d01b9014202bf02f002c4024b029901c300;
    decBuf[8574] = 256'h33007cff35fff4fe2fffacffa000da0155035404820458044b0357027a01ea00;
    decBuf[8575] = 256'h3901af014702d0020603f502e702bf02cb02ec020a034a039403da033e049c04;
    decBuf[8576] = 256'hf1041205e0047b04e80338039102500216024b027c02e3022603630358033a03;
    decBuf[8577] = 256'h310339035e039c03f703340481049f04ba04c204ca04b50496044104bc03f702;
    decBuf[8578] = 256'h0c026e01180166013c02eb039c0524072308af08300870077c069f0549052e05;
    decBuf[8579] = 256'h17050105ed049404430434045c04e20482051a06a306b5066406df053e05d204;
    decBuf[8580] = 256'he604630536063907a1074307b306c805ea0494047a04c104d704ea04b5048404;
    decBuf[8581] = 256'h9304bb044005e105790602077f07d0075508d20844098e0930097a08f2068904;
    decBuf[8582] = 256'hee020d02c901fe02f7045b079b09110b550b170b6f0ad6094b092009fa089108;
    decBuf[8583] = 256'h75071b067a04f1025802e3020a044a06e507f009bc0a7f0a6609010860064705;
    decBuf[8584] = 256'h1405e60464052406d2063107c107db0722086308770865081408360759065605;
    decBuf[8585] = 256'ha80449046604e804ee0527074e08a809900a620b220c450ce60be30aa909da07;
    decBuf[8586] = 256'hae053904e502a702df0278031905a2066d081d0a360b350c630c390c2d0b6709;
    decBuf[8587] = 256'h3c0730055403200277011002f8027304d8051d07ef0763088508e4083b095509;
    decBuf[8588] = 256'h3d09a608a6076d0646053904d003b10307048a043005f305de06bb0784080709;
    decBuf[8589] = 256'h1f09090980089707ba06b705c304e6038f037503ec03af049a057706cd061c07;
    decBuf[8590] = 256'h3407f306df06a9067906f4052f05100403035502f6014c02030338045f051f06;
    decBuf[8591] = 256'h8706a706170660058b04c1030a039402530266029c022e03b8035904f0047905;
    decBuf[8592] = 256'haf05bf057505e20432048b034b03100322035203610354032f030e032c039103;
    decBuf[8593] = 256'h09045a042e04b60303032d029d014f019601d7013902b602e702f602e902c402;
    decBuf[8594] = 256'h8d023302c6015f010101f50000010a010101d800b2009e00b00005018a01e301;
    decBuf[8595] = 256'h1402e8015501a400feff67ff2cff61ffd3ffb000cd01da02ce032d049d03b202;
    decBuf[8596] = 256'h56011100eafe2afec2fde1fd38febafe61ff23000e012b02eb02530334036b02;
    decBuf[8597] = 256'h4b01f2ffadfe86fdc6fca4fcc3fc8cfd78fe94ffa10009012901d300e8ffcbfe;
    decBuf[8598] = 256'hbefd10fdb1fccefc51fdf7fdb9fe70ffb8ffcdffbaff84ff33ffe9fea6fe51fe;
    decBuf[8599] = 256'h1afec0fd6bfd08fdc5fcb9fcdafc70fd33fe1efffbffc50047013001c300ecff;
    decBuf[8600] = 256'haffe34fdcffbe7fa15fa3bfae9fac7fbcafc78fd16fe6cfe86fe9efe89fe75fe;
    decBuf[8601] = 256'h1cfecafd28fd91fc07fcaefbbefbeafb2dfc39fc18fcfafb16fc71fc26fd12fe;
    decBuf[8602] = 256'heffe45fff7fef2fdb8fc3dfb3efa6cfaeafa44fc88fd03ff9cffcbfff8fe9ffd;
    decBuf[8603] = 256'h5afc88fb14fbf2fa11fba1fbbbfb02fcedfb28fc5dfccffc54fdadfdfefdf0fd;
    decBuf[8604] = 256'hadfd58fdc9fc3ffc9ffb07fb7efa01fa8ff963f970f9adf93cfa14fb16fc50fd;
    decBuf[8605] = 256'h23fe96feb9fe99fe09fe87fdb1fce8fbfdfa1ffa90f941f959f91cfa3bfb48fc;
    decBuf[8606] = 256'h81fd54fe7afe58feb9fd2afd73fccdfb8cfb78fbaefbbefbcdfba5fb80fb75fb;
    decBuf[8607] = 256'ha7fb30fc2ffd23fe82fe2cfe75fd11fcacfac4f946f96cf91afaf8fafafbeffc;
    decBuf[8608] = 256'h8dfd56fed9fef0fedbfe2afef5fc7afb15fa2df9aff822f9d0f9edfafafbeefc;
    decBuf[8609] = 256'h8cfd1cfe6afeb1fe9cfe88fe52fec0fde8fce6fbacfad9f966f989f966fa2ffb;
    decBuf[8610] = 256'h4ffc0ffd77fd97fd7afdc9fde0fd21fe0efeb4fd01fdfcfb08fb6afa4dfa04fb;
    decBuf[8611] = 256'hdafbddfc8bfdeafdcdfd4afda4fc0dfcabfb75fb85fbb2fbf4fb62fcabfc09fd;
    decBuf[8612] = 256'h46fd7dfd9bfda4fd6afd17fdcafc84fc57fc70fca4fce2fc0bfde6fca8fc4dfc;
    decBuf[8613] = 256'h10fc31fcb3fc78fd2ffed5fe41ff06ff66fea3fdecfc75fc34fc21fc7afccbfc;
    decBuf[8614] = 256'hf8fceafcc6fc79fc33fcf3fbdafb00fc3efca9fc2efdcffd66fec8fefefecdfe;
    decBuf[8615] = 256'h48fe84fd98fcbbfbf2faa3fa8cfaf8faa8fbaefc5cfd39fe90fe76fefffd93fd;
    decBuf[8616] = 256'h31fd1ffd2ffd96fdbefdb2fd65fde3fc8afc7afcc3fc3cfdcefd09fef7fdc6fd;
    decBuf[8617] = 256'h5ffde7fcb6fca7fceafc57fddcfd35fe66fe57fefafd8cfd08fdd2fcc2fcd1fc;
    decBuf[8618] = 256'hf9fc35fd6cfd8afda6fdcffdd6fdc2fd8afd46fd06fdddfc02fd33fd84fdd1fd;
    decBuf[8619] = 256'heffd0afe33fe68fea6fecffed7fe99fe1dfe7cfdb9fc37fcf0fbdafb3cfcddfc;
    decBuf[8620] = 256'hcbfda8fe38ffbbff0200ecff8affe9fe27fe3bfd9dfc0efcbffb06fc47fcd1fc;
    decBuf[8621] = 256'h95fd18febefe2aff65ff9bff8bff41ffaefeaffdbafc1cfcc6fb14fcbbfc7dfd;
    decBuf[8622] = 256'h34fedafe72ffd4ff0a003a002c00ceff30ff6efe83fde4fc55fc3bfc82fceefc;
    decBuf[8623] = 256'h9ffd74fe3eff29008800de00c4004d00e1ff57ffb7fe4afec1fd8bfd5bfd69fd;
    decBuf[8624] = 256'hc7fd34fe9bfedefe03ff3aff6cffe2ff7500fe001001bf00ffffdffe20fe71fd;
    decBuf[8625] = 256'h52fda8fdf6fd6dfed9fe3bff71ffc2ff0c0019000d00aaff32ffc0fe59fe4bfe;
    decBuf[8626] = 256'ha0fe03ff96ff20005500660057001400d7ffb6ff84ff69ff40fffcfebcfe83fe;
    decBuf[8627] = 256'h7bfeb9fe35ffd6ff98001b0192017c0168010f01be009100690045002400deff;
    decBuf[8628] = 256'h8cff3fffe5fec0fee1fe27ff9eff5100f700ba013c02b302c9028e02c901de00;
    decBuf[8629] = 256'hc1ff02ff53fe34fec3feaeff8c008f01f70156023902eb01a4013801ae003100;
    decBuf[8630] = 256'hbfff58ff4bff87ff2c00610188029503fd031d048d03a20285012c00e7fe69fe;
    decBuf[8631] = 256'h43fe65fe43ff0c002b0138022c03ca0321043b04f3033103460229011c006eff;
    decBuf[8632] = 256'h0fff2cffafff84004e013902d702f4020e03c60286022302ca0179016a015d01;
    decBuf[8633] = 256'h8101b80112027f02e60229031d03d00276020902dd01cf010c02430261026a02;
    decBuf[8634] = 256'h41020c02ea01f0012e0299021e03bf0300043b0405047303c2021c0285012301;
    decBuf[8635] = 256'h110121016b01e3015502bc023403a6030d04360411049803e5026f020302ef01;
    decBuf[8636] = 256'h4802ba0221037f03bc039b035503de024c029b0154013e017901f601c9029303;
    decBuf[8637] = 256'h15045d0472041004b70365031c03d902b402a9029f02bb02f50229033e034403;
    decBuf[8638] = 256'h1103c6028002400238026c02d3025803d5036704c904ff040f05e3046b04b803;
    decBuf[8639] = 256'he202190262014a016001e901ae026503dc0348045b046d045d044e0441041c04;
    decBuf[8640] = 256'hcf0375030803a1022902f801e901f7014b02c4025703e0035d04cf04de04b604;
    decBuf[8641] = 256'h6104d2034803a7023b0228021602470273029b02bf02e0022603af0387045005;
    decBuf[8642] = 256'h07061f0688056104e602810199001b004100f0000c02cc027a0319046f04bd04;
    decBuf[8643] = 256'hd504eb04b00433048003da026d02330268029902c502d30296025f0255028302;
    decBuf[8644] = 256'hee027303f003410450040d04a0033803f602e902f402120352036b0382038803;
    decBuf[8645] = 256'h76037b036c035e033803eb0288021002be01b0010d0293023303cb030604f403;
    decBuf[8646] = 256'hc3037903510345033a031c03ca0251029e012701bb00a800010193011d02e102;
    decBuf[8647] = 256'h98033e04ab04be04ac045b04b90321039802f7018b0150011b010a0137015f01;
    decBuf[8648] = 256'hb40101025b02af0212037003c503fc030604d8037e03e0021d029b01f400b400;
    decBuf[8649] = 256'hc7002101b3016302da021b032f03d5026402fc01b9019501a001be01fe013802;
    decBuf[8650] = 256'h8a02c102f302fc02d302810208027501c5004e0038004c00ed00af0166023c03;
    decBuf[8651] = 256'h9203ac0336039e02150298012601dc009900450024004200a6005401fa019102;
    decBuf[8652] = 256'hcc02970204025401ae0041002e006300d5003c019a01be01df01d501ba01a101;
    decBuf[8653] = 256'h8b015b012201df008d004000e6ffa9ff9effa8ff0d00a0005001f7018e021703;
    decBuf[8654] = 256'h0503b4021202f9009fffb8fee5fdbffde1fdbffe88ffa7006701160275029102;
    decBuf[8655] = 256'h77023002c4013a017600bfff19ff81fe1ffeeafd1afe82fe4aff4d004101df01;
    decBuf[8656] = 256'h35025002d90116015f008afffafeabfe64fe7afe8dfec3fed3fe00ff5dffcaff;
    decBuf[8657] = 256'h4f00cc001d012c01e900330048ff6bfea2fdebfcd3fc14fd9dfd62fe4dff6a00;
    decBuf[8658] = 256'h2a019201f101d4011d011800defe63fd64fc7cfba6fb1afc0efd6afeaeffd500;
    decBuf[8659] = 256'h9501b8019801cf00180013ff1ffe02fd42fcdafbf9fb89fc40fd45fe39ffd7ff;
    decBuf[8660] = 256'hf4ffdaff93ff27ff9dfe68fe37fe46fe38fefcfdaffd55fd18fd0dfd3ffdb6fd;
    decBuf[8661] = 256'h48feaafee0fef0fec4fe81fe44fe23fef1fdb1fd88fd53fd31fd1efd2ffd5dfd;
    decBuf[8662] = 256'haffdfcfd56fe92feb3fea9fe7cfe31fec3fd5cfde4fc92fc49fc3bfc60fcadfc;
    decBuf[8663] = 256'h43fddafd63fe99fea9fe60fee7fd75fdf1fc97fc46fc55fc7dfcd2fc1ffd8dfd;
    decBuf[8664] = 256'hb9fde1fdd5fd9efd80fd65fd5cfd64fd79fd8bfd86fd76fd56fd30fd0cfdebfc;
    decBuf[8665] = 256'hd6fce2fcfafc23fd4afd5afd55fd37fd1cfd19fd3bfd77fdb1fde5fdd1fd8cfd;
    decBuf[8666] = 256'h15fda4fc1ffce9fbfafb43fca1fc0efd75fdd3fddffdd4fdb6fd88fd70fd77fd;
    decBuf[8667] = 256'h70fd5efd20fdb4fc30fcb3fb82fb91fb09fc9bfc4cfdc3fd2ffe42fe0dfefcfd;
    decBuf[8668] = 256'hb3fd8bfd66fd5bfd3dfd10fdc5fc6bfce6fb8dfb7cfbc6fb3efcf1fc97fdd8fd;
    decBuf[8669] = 256'hecfdb6fd65fd39fd11fd35fd56fd88fda3fdacfd95fd65fd20fdcefc6bfc28fc;
    decBuf[8670] = 256'hecfbf7fb15fc67fce0fc52fdd6fd30fe60fe6ffe2cfebffd3afdbdfc8dfc9bfc;
    decBuf[8671] = 256'hdefc33fd6afd60fd20fdc5fc58fc2cfc54fc91fc0afd7cfdc5fd23fe2ffe50fe;
    decBuf[8672] = 256'h5afe3ffe15fee1fd7afdf5fc9cfc2afcfefb26fc7bfcdefc3bfd60fd55fd37fd;
    decBuf[8673] = 256'h09fd11fd55fdb9fd32fe83feaffe87fe32feb9fd47fde0fc82fc46fc0ffcf1fb;
    decBuf[8674] = 256'he8fb11fc54fcb9fc4cfdfdfda3fe0fff4aff38ffe7fe44feadfd24fda7fc55fc;
    decBuf[8675] = 256'h47fc39fc45fc7cfcc2fc14fd77fdd5fd12fe49fe7bfebbfe05ff4bff66ff3dff;
    decBuf[8676] = 256'hccfed9fde5fc07fc77fb5dfba5fb11fcc1fc97fd27fea9fe20ff36ff22ffedfe;
    decBuf[8677] = 256'h9bfe34febcfd6afd03fddbfcb7fcd8fc0afd6efdccfd21fe58fe4efe20fed6fd;
    decBuf[8678] = 256'hb8fdaffde8fd3bfe9efee1feedfeb6fe34feb7fd45fdfbfceefc2afd61fdbbfd;
    decBuf[8679] = 256'hf8fd2ffe61fea1fecafefffef8fec0fe5efee6fd74fd48fd55fdc2fd29fe87fe;
    decBuf[8680] = 256'habfea0fe46fef2fdbbfdb1fddefd18fe4cfe61fe4efe10fee7fdeffd2dfe98fe;
    decBuf[8681] = 256'h1dff9affcaffbcff79ff0cffc2fe7ffe5bfe24fef2fdb2fd57fd33fd3efd98fd;
    decBuf[8682] = 256'h35fef8feafff55009600aa005000beff35ffdbfe69fe20feddfda0fd69fd73fd;
    decBuf[8683] = 256'ha1fd1dfebdfe80ff03004a008b0050001a00c9ff7fff22ffe5fe82fe3ffe1bfe;
    decBuf[8684] = 256'hfafd04fe31fe7cfeeafe6effecff3d0069005c003700eaff90ff3bff04ffd2fe;
    decBuf[8685] = 256'hc9fed2fe06ff6dffd4ff3200870092007400100097ff25ffdcfeb4fea7fedefe;
    decBuf[8686] = 256'h38ffa6ff2a00a700d8000401f700ba006d002700e8ffaeff88ff74ff61ff72ff;
    decBuf[8687] = 256'ha0fff1ff5400b200ee0025012f012601fd00ab0048000500b0ff8fff85ffb2ff;
    decBuf[8688] = 256'h0d006200c5000801450150015a013e011501ef00cd00a10090008b009000a500;
    decBuf[8689] = 256'hc800f20019013301410145013101190109010c0119013801560171017c016c01;
    decBuf[8690] = 256'h4c011e01f200ca00d000e7001e016101a101cb01e101da01bb01aa019b019f01;
    decBuf[8691] = 256'ha401a701a401a101a401b101d401f801fd01df01a5014a0126011b014d019f01;
    decBuf[8692] = 256'h18028a02f10219033e0333031503c2025f02e70175012c011e014301a6010302;
    decBuf[8693] = 256'h7002d80235037203930375032303aa0217028e01350124015101ae011b028302;
    decBuf[8694] = 256'he0024d039703bf03e403ef03d1039103150398020602a4014a015a01a4013702;
    decBuf[8695] = 256'he8028e03cf030a04d403a40377034f035b03500332031703dd02b802b102d002;
    decBuf[8696] = 256'h0303330339031203d902a5029e02e3024703bf0331045d041b04ad032903ac02;
    decBuf[8697] = 256'h9b02c8024003b20319042604ea037103ff02b5028d028102a202c002db020503;
    decBuf[8698] = 256'h4803bf03510402057805e405d105540580047e0344027101fe00db003a010302;
    decBuf[8699] = 256'hee020b04cb047905d805bb056d05f60434047d0306039a025f024d025d028a02;
    decBuf[8700] = 256'hcd0221038403fd034e0498048a0466041904ab0361033903450366039803d803;
    decBuf[8701] = 256'h010418041104e50391032403bd029402a102d8025a03d703480457044a04f503;
    decBuf[8702] = 256'h92034f035b03920300044a0457041b04a2030f03860250028102e8026103b203;
    decBuf[8703] = 256'hde03d103940373037d039903d203e903d403b503820360035a0354033b030803;
    decBuf[8704] = 256'hbc0262023e025f02b90226038d03d003dc03a503730345032d03340357036903;
    decBuf[8705] = 256'h58032003bf024602f501e601f4014802c10233035f0388037b035a0364038003;
    decBuf[8706] = 256'h9903af039a035603df024d02eb016e015d016c01ca011f028202df0204032503;
    decBuf[8707] = 256'h1b03ff02e602df02ca02c402b30285024d02fa01ad0153012f01240156019601;
    decBuf[8708] = 256'hf10145026602700267025f0267027b029a02a00286024a02f0019b0164015a01;
    decBuf[8709] = 256'h63016b0164015d014a0144016801a401de0122023d0256025d0264026a025902;
    decBuf[8710] = 256'h2102cf015601e4007d001f00fbfff0ff0e004d00b9005b01f20154028a027a02;
    decBuf[8711] = 256'h3002b8014601c10068001700eaffddff01004e00a800fd003401520149013001;
    decBuf[8712] = 256'h0b01f600ca00a3007f0068006c008700ae00c800c300ae0093007a0077008500;
    decBuf[8713] = 256'h9d00a00092006a002100dbff9bff83ff8affc8ff12006c00a900e000d600a800;
    decBuf[8714] = 256'h5e000400c7ff90ff72ff57ff5fff67ff7bff9bffabffa6ff98ff83ff7fff91ff;
    decBuf[8715] = 256'hc0ff0b003d0059002f00ecff88ff2affedfee2feecfe2cff66ff9affbdffd0ff;
    decBuf[8716] = 256'hcaffbbff91ff6aff31ff0cffe9fed7fedcfeecfe15ff3dff56ff77ff8cff88ff;
    decBuf[8717] = 256'h7dff5bff31fffffec1fe87fe35fefefdccfdc3fdecfd4dfec6fe37ff9fffc7ff;
    decBuf[8718] = 256'hbbff84ff2affbdfe55feddfd8cfd5ffd52fd5efd95fdeffd44fea7feeafe0eff;
    decBuf[8719] = 256'h19ff0ffff4fecbfe96fe74fe61fe3afe16fee3fdb3fd94fd8efd93fdaafdc8fd;
    decBuf[8720] = 256'hf3fd1afe48fe80fea6febafe9bfe52fef8fd8bfd41fd19fd0dfd18fd36fd64fd;
    decBuf[8721] = 256'h9dfdc3fdd7fddefdc2fd89fd37fd00fdcefcc5fceefc22fd60fd9afdbffdd4fd;
    decBuf[8722] = 256'he7fdecfdf2fddafdb4fd67fdeefc7dfcf8fb9efbaffbdbfb6efc1ffdc5fd5cfe;
    decBuf[8723] = 256'hbefed0fea0fe56feddfd6cfd04fda7fc3afcd2fb90fb53fb48fb7afbdefb71fc;
    decBuf[8724] = 256'hfbfc9cfdddfdf0fdbbfd69fd02fdbffc6afc1dfcebfbbefba5fb9dfbb2fbeafb;
    decBuf[8725] = 256'h2efc5bfc64fc4dfc1dfcf1fbecfb24fc77fcc4fc0afd25fdfcfcc7fc7cfc4afc;
    decBuf[8726] = 256'h2efc15fc0efc15fc28fc38fc3efc26fceffbbbfb8bfb91fbcffb29fc97fce0fc;
    decBuf[8727] = 256'hd3fcaffc78fc46fc18fc10fc17fc10fcf1fbbefb73fb19fbc4fa77fa45fa60fa;
    decBuf[8728] = 256'hccfa6efb30fce7fc2ffd44fd09fdb0fc3efcd7fb94fb57fb36fb04fbc5fa8bfa;
    decBuf[8729] = 256'h65fa7afab2fa23fbd5fbabfc3bfd89fd72fd31fdcffc51fce0fb78fb50fb44fb;
    decBuf[8730] = 256'h39fb2ffb26fb0dfb06fb1afb46fb9bfb08fc6ffcb2fcbefcb3fc6dfc1bfccefb;
    decBuf[8731] = 256'h88fb6cfb75fb6dfb66fb3bfb13fbdbfac4facbfa03fb56fbb9fbfcfb38fc6ffc;
    decBuf[8732] = 256'ha1fcbdfcb5fc8ffc43fce9fb7cfb15fbedfaf9fa1afb60fbc4fb22fc77fcaefc;
    decBuf[8733] = 256'hb8fcc1fcc9fcc2fcc9fcdbfcd6fcbcfc77fcf5fb9bfb4afb59fb9cfb09fc70fc;
    decBuf[8734] = 256'hb3fcbffc9efc6cfc51fc49fc50fc65fc77fc88fc8dfc80fc6afc47fc27fc12fc;
    decBuf[8735] = 256'h0efc18fc35fc50fc68fc84fc98fca9fcbffcc2fcb5fca9fc9efc9cfcb7fce9fc;
    decBuf[8736] = 256'h27fd61fda4fdd2fdeafdf2fdddfda5fd53fddafc88fc7afc87fcf4fc79fdf6fd;
    decBuf[8737] = 256'h47fe56fe2efef1fdbafdc4fde0fd09fe1ffe18fee0fd8efd2bfdcdfca9fcb4fc;
    decBuf[8738] = 256'hfafc5efdbcfd11fe48fe52fe36fe1dfe16fe1dfe30fe40fe50fe4bfe36fe23fe;
    decBuf[8739] = 256'h0afefafdfdfd05fe11fe28fe57fea3fe11ff78ffd6ff1200f1ffbfff6dff20ff;
    decBuf[8740] = 256'h02fff9fe01ff09ffe7fec7feabfeb0feecfe58ffdcff5a00ab00d700af004200;
    decBuf[8741] = 256'hbdff1cff85fe4afe38fe69feb3fe2bff9dff04007c00ad00d900cc008f005800;
    decBuf[8742] = 256'hfeffa9ff5cff2aff21ff4bffacff3f00a100fb002b011d01f500e800f3002501;
    decBuf[8743] = 256'h65018f01960174013b01f800ca00b200aa00cc00050139015c017b018c01b001;
    decBuf[8744] = 256'hec0136029002b402a9024f02b201ef006c002500100099003a01d1015b02b402;
    decBuf[8745] = 256'ha40295026d0248023d021f02f201b80166012f0125015201bd014202bf021103;
    decBuf[8746] = 256'h5a0382038f039a0368033a03df028a023d021f0216025002c0025303dc037d04;
    decBuf[8747] = 256'hbe04aa04750403047e030103d002df02070344039103c303cc03b3038e035003;
    decBuf[8748] = 256'h37034d037e03cf031c043a0443041a04c7037a0334030703fe02240354039903;
    decBuf[8749] = 256'hd903120438044c04530458045d046b049204c004eb0408050205e204ab047604;
    decBuf[8750] = 256'h38040f04170439048a0403055505bc05e405d805b70599056b0563053d050d05;
    decBuf[8751] = 256'hd50483044c041a04100419043e0461048c04d5042f058405e7050f060306cc05;
    decBuf[8752] = 256'h4a05a904e70364034c036203eb038c042405ad05e305f305e405bc05b005a505;
    decBuf[8753] = 256'h9b05a4058b05660536050a05ee04f30426058d0512066b06bc06e906a6065106;
    decBuf[8754] = 256'hc2053805bb048b047c04bf0414058d05fe054806550649062806ce056105fa04;
    decBuf[8755] = 256'h8204300404042c046904b604fc04290542054a0551057c059805a805ac059705;
    decBuf[8756] = 256'h65052705dd04970457044f047404cd045305ac05fd050c06e405a70586056805;
    decBuf[8757] = 256'h84059d05c205d705dd05cc05a80575052a05e40492045b043d0446046f04c104;
    decBuf[8758] = 256'h0e0568058d05980566051405c7046d0448041104df03b203780352034c035e03;
    decBuf[8759] = 256'ha70315049a041705890598055505e8046304c20356031b0309035b03c2033a04;
    decBuf[8760] = 256'hac04f6041e052a050905d704a90470041d04d0039e0383039b03c103f1031d04;
    decBuf[8761] = 256'h2e041404f403d603d203eb03f403da03a603350382020c02f6010a0287021903;
    decBuf[8762] = 256'ha203fc03eb03a2030f0385020802d701c9010b0248027f029d02820269025202;
    decBuf[8763] = 256'h7502ad020003370341030103a60251020402fa012802510285029a02a0029b02;
    decBuf[8764] = 256'h8b027d0271025d023e022002fd01dd01bf01a401a001b001d001ed01f101d901;
    decBuf[8765] = 256'haa015101fc00db00d100da00e200f900f200d200ab008700670063007e00ab00;
    decBuf[8766] = 256'hd700e800ce009200480016000d0036006a009b00ad00a8008e0077006a006e00;
    decBuf[8767] = 256'h80009500aa00a20088006800420028002d0042005d005a003700fbffc1ff8dff;
    decBuf[8768] = 256'h86ff99ffaaffa5ff84ff55ff2aff0efffefefafe06ff0aff07fff1fec6fe8dfe;
    decBuf[8769] = 256'h4afe2ffe26fe4cfe7cfeb4fecbfec4fe98fe7cfe58fe4afe46fe3afe37fe2dfe;
    decBuf[8770] = 256'h2bfe42fe65fe85fea3fea7fe9cfe80fe65fe53fe4afe47fe4afe47fe30fe07fe;
    decBuf[8771] = 256'he0fdb2fd93fd8dfd9cfdbdfddafdeefdeafdd4fda9fd65fd12fdc5fc6bfc47fc;
    decBuf[8772] = 256'h3cfc6efcc0fc0dfd3ffd5bfd31fdeefcaefc64fc32fc16fcfefbf6fbeffbe9fb;
    decBuf[8773] = 256'hfafb32fc85fce8fc2bfd37fd2cfdd2fc7dfc1afcf2fbcdfbd8fbe2fbebfbf4fb;
    decBuf[8774] = 256'h0afc11fc3dfc6ffcadfcc6fccefc9dfc4cfce9fb8cfb67fb5cfb66fb82fb9afb;
    decBuf[8775] = 256'ha2fb8dfb7afb5efb4ffb54fb60fb74fb7efb6ffb49fb11fbcdfaa0fa87fa70fa;
    decBuf[8776] = 256'h85faa4fac0fae4fa0efb1ffb2efb2afbfbfac3fa8efa79fa73fa84fa9efab5fa;
    decBuf[8777] = 256'hcafad6fae0faf0faedfaf0faf7faecfaeafae8fad6fac6fab7faa9faa4faacfa;
    decBuf[8778] = 256'haafaacfaa5fa97fa99faacfaa9fa9efa7efa42fa18fa02fa09fa28fa44fa49fa;
    decBuf[8779] = 256'h29fa03fad4f9b5f9bbf9caf9d8f9e5f9e9f9e5f9e8f9ebf9fef918fa37fa4cfa;
    decBuf[8780] = 256'h58fa39fa01facdf99df996f9bef90bfa58fa9efab9fab1fa9afa86fa7ffa85fa;
    decBuf[8781] = 256'h80fa69fa54fa19fae0f9c9f9c2f9e2f91ffa6afab0facbfac3fa8efa50fa17fa;
    decBuf[8782] = 256'h00faf9f900fa05fa00fae9f9cbf9c0f9b5f9bef9e4f908fa31fa59fa68fa51fa;
    decBuf[8783] = 256'h2bfaf2f9dcf9e3f9f5f91dfa41fa4ffa53fa5efa62fa78fa97faa4fab8fac9fa;
    decBuf[8784] = 256'hccfabefab6faa1fa92fa8afa8dfaa8facbfad9fae6faf1faf5fa11fb34fb4bfb;
    decBuf[8785] = 256'h4ffb2cfbe7faa1fa73fa6bfa91facffa08fb2efb42fb30fb14fb0efb01fbfcfa;
    decBuf[8786] = 256'h00fbfdfa00fb03fbfbfa02fb0dfb17fb2dfb49fb55fb6efb77fb6efb71fb7dfb;
    decBuf[8787] = 256'h87fb9dfbacfba4fb98fb8dfb8ffbaafbe4fb3ffc7bfc86fc7cfc61fc38fc12fc;
    decBuf[8788] = 256'hfdfb04fc15fc38fc59fc6efc89fc8dfc8afc92fc9ffca6fcadfcabfc91fc75fc;
    decBuf[8789] = 256'h64fc54fc5dfc7afc95fcb4fccafcd5fce0fce3fcd5fccdfccffcd5fceffc0ffd;
    decBuf[8790] = 256'h2dfd40fd44fd40fd43fd4bfd5cfd7cfd9cfda9fdb4fdaafd9afd8cfd94fdb3fd;
    decBuf[8791] = 256'hf2fd32fe6cfe83fe6efe29fefcfde3fd08fe46fe90fec2feccfea2fe6efe59fe;
    decBuf[8792] = 256'h53fe6ffe9dfec9fef0fef5fee8fecafeaffe96fe93feadfed3fe02ff21ff3dff;
    decBuf[8793] = 256'h42ff47ff4bff4fff4bff3cff22ff10ff13ff3fff83ffd5ff0c002a0034001b00;
    decBuf[8794] = 256'hf5ffd3ffc0ffc6ffd5ffffff2600400060007e00a100c100d600ea00e600d700;
    decBuf[8795] = 256'hbd00ab00a800b700d300f6000401110115011f012f0143015b016a0173017001;
    decBuf[8796] = 256'h77017e0184019401960188017801720170018301a501c501ec01050213022002;
    decBuf[8797] = 256'h2b0236024c02660270026d02530226020602f60119025f02cd02340377036b03;
    decBuf[8798] = 256'h4a032c03fe02f6020c032f034203470338032103250338035f03ac03e3031504;
    decBuf[8799] = 256'h1e040504c2038203580351038103ad03df030204080402040804150422043604;
    decBuf[8800] = 256'h390423040f04fd03f6030d042f0459048c04bc04ce04df04e404d704d204ce04;
    decBuf[8801] = 256'hc404b404a60494049604ad04dc041a05540579059c05a20591058c057e054f05;
    decBuf[8802] = 256'h2405fc04d804dd040c055005a305f00522062b061206dd05ad0582055a055505;
    decBuf[8803] = 256'h630578059305b305c805e305f505040613061006040602060006050617061e06;
    decBuf[8804] = 256'h0b06f905d505a705a105a605d5050d0650067e069706ad06a606a0068f066b06;
    decBuf[8805] = 256'h5d0640061506f905ea05ee05140643067b06af06c406be06a20688067a068706;
    decBuf[8806] = 256'ha206b306b006850640060106d705d0050e066806bd060a071407e7069c065606;
    decBuf[8807] = 256'h17060e06250647065a0654061c06f605e205e8051b066606ac06da06d206ac06;
    decBuf[8808] = 256'h7c0637060a06f105f8050d062c063d06420650064c0648065306620671067e06;
    decBuf[8809] = 256'h7b06600645061e06f005dd05cc05bd05c205d705e20502060f061a061e061406;
    decBuf[8810] = 256'h0006ee05d405ad0594057305560542053f0548056d059105b205cf05d305b405;
    decBuf[8811] = 256'h8e05550521050c05f9040a0524054405510555054a0534052605190508050605;
    decBuf[8812] = 256'hfc04ec04e604dc04cc04ca04c004b704c004ca04ce04d704d104c204a2048204;
    decBuf[8813] = 256'h640449042a04140409040c041604300441043e0441043904320427041104ec03;
    decBuf[8814] = 256'hbe03850351033c034303530377039803ad03c003bd03a7038703610333031403;
    decBuf[8815] = 256'h0303f302e602c802bc02c702e30206032f034b0346032f030003bc028e025402;
    decBuf[8816] = 256'h3e0229022f02400245025302580263026e0271027402670243021f02ec01bc01;
    decBuf[8817] = 256'h9d018101670150014301470160018201ac01bc01c201a1017b014d011501ef00;
    decBuf[8818] = 256'hcd00ad009d0097009c00a900c400e300010115011101f500bb0081003e001000;
    decBuf[8819] = 256'h08000f002400430049004e0049003c0039004300460038001600daff8fff5dff;
    decBuf[8820] = 256'h30ff27ff4dff7dffb5ffccffd3ffb3ff76ff3cff16fff4feeefee8feedfee9fe;
    decBuf[8821] = 256'hdcfec1fea8fea5feaefec0feccfecefec4feadfe97fe83fe61fe38fe10fee2fd;
    decBuf[8822] = 256'hcffdd5fdf9fd2cfe5cfe6ffe69fe4ffe26fefefde5fdcefdb8fda5fd93fd8afd;
    decBuf[8823] = 256'h7cfd7efd8afda2fdbefdd9fddcfdcdfda7fd79fd41fd1bfdf9fcdafcd4fccffc;
    decBuf[8824] = 256'hd4fcd8fce4fce7fcf0fceefcf0fcf7fcedfccffca8fc70fc3cfc19fc06fc0cfc;
    decBuf[8825] = 256'h26fc46fc64fc8efcabfcbafcbffca1fc6efc3efc13fcf6fbf1fbedfbf1fbf5fb;
    decBuf[8826] = 256'hf1fbfbfb1afc38fc5bfc7bfc77fc5cfc2efceafb98fb61fb43fb39fb63fb97fb;
    decBuf[8827] = 256'hbafbd9fbbdfba3fb95fb88fb85fb8ffb8cfb7efb6bfb4cfb37fb24fb19fb0afb;
    decBuf[8828] = 256'h07fb09fb1afb3afb63fb8bfba4fb97fb79fb5efb37fb1efb10fb03fbf7fafbfa;
    decBuf[8829] = 256'hf8fafbfa08fb0ffb22fb3ffb5afb72fb76fb5cfb27fbf3fab5fa9cfa95fa9bfa;
    decBuf[8830] = 256'hbbfad7fae6faf4fa09fb15fb34fb52fb56fb4cfb2ffbf5faabfa79fa5efa66fa;
    decBuf[8831] = 256'ha9fae9fa23fb58fb5efb58fb47fb38fb21fb14fbf9fad9fab3fa85fa66fa6bfa;
    decBuf[8832] = 256'h71fa91fac8fafdfa2dfb4cfb5dfb58fb4afb24fb00fbcdfa9dfa8afa84fa9efa;
    decBuf[8833] = 256'hd1fa0ffb38fb5efb72fb85fb8bfb90fb82fb6dfb59fb33fb0ffb01fbf4fa00fb;
    decBuf[8834] = 256'h26fb54fb80fb9cfb97fb80fb6bfb57fb54fb5dfb55fb4dfb3cfb1cfbf3fae2fa;
    decBuf[8835] = 256'he7fa07fb47fb87fbb0fbd6fbddfbb1fb95fb67fb54fb4efb53fb61fb6efb81fb;
    decBuf[8836] = 256'ha1fbd8fb0dfc2ffc5bfc6cfc71fc63fc4efc2bfc01fcc3fb9afb92fb99fbc5fb;
    decBuf[8837] = 256'h0efc40fc6efc97fc9ffc98fc85fc52fc22fcf6fbdafbd5fbd1fbccfbd0fbe2fb;
    decBuf[8838] = 256'hfefb38fc82fcb4fce2fcfbfce4fcc2fca2fc86fc77fc72fc6efc72fc8afca7fc;
    decBuf[8839] = 256'hd1fc04fd34fd6cfd92fda6fda0fd79fd36fdf6fcbcfca6fc9ffcbefcdafcfefc;
    decBuf[8840] = 256'h31fd61fd8dfdb4fdbafdb5fd97fd65fd35fd15fd05fd0afd2afd3ffd5afd6cfd;
    decBuf[8841] = 256'h7cfd95fdc3fdfbfd3ffe6cfe75fe6dfe3dfe05fec1fda6fd8dfda4fdc6fdfefd;
    decBuf[8842] = 256'h24fe46fe65fe81fe9bfeb2fec7fec4fea4fe75fe31fe03fedafde1fde8fd07fe;
    decBuf[8843] = 256'h3afe5cfe95fec9feebfe0bff27ff22ff1dfffffed5feadfe89fe85fea3fed5fe;
    decBuf[8844] = 256'h13ff5dff8fffbdffd5ffddffe4ffd1ffb5ff87ff5bff28ff06ff00ff11ff2aff;
    decBuf[8845] = 256'h5dff8dffb9ffd5ffeffffdff0900feffe5ffb6ff79ff3fff28ff21ff4dff8bff;
    decBuf[8846] = 256'he6ff3b007200a400bf00c700b10081005500390029003700550070009000a500;
    decBuf[8847] = 256'hb800d800f600200148015701520146012301f000b200890063005c006f00a200;
    decBuf[8848] = 256'he00009012e0135012f0129012401160112010e01fd00ed00e400f20015015801;
    decBuf[8849] = 256'haa01f7013d0246022d020802d801b801b301c201d901ef01f201fd0106021502;
    decBuf[8850] = 256'h3c026f029102b0029f0271022d02da01a30185018f01b801dd010d0239026c02;
    decBuf[8851] = 256'h8e02a102b202ad02960280026d02540245023602340249027402b902f9023303;
    decBuf[8852] = 256'h58036d0373036d035e033e031703f402ca02ae029e02ac02d30201032c034903;
    decBuf[8853] = 256'h6c0371036d03590348032c030903e902c202b302c102df02190352038703a903;
    decBuf[8854] = 256'hbc03c203c703c203be03b2039a037e03630351034e0362038403ae03ec031504;
    decBuf[8855] = 256'h3a044f04490421040804de03ac0389035d0341033c034a035f038203a303c003;
    decBuf[8856] = 256'he303040421042d042204f403b6038c036703600373038f03b303e60324046e04;
    decBuf[8857] = 256'ha004a904a1046c043c041d040c0407040204ed03da03e40300042b045d047204;
    decBuf[8858] = 256'h78045c043804fc03d303ad03990393038d039c03aa03b703ca03e30305042604;
    decBuf[8859] = 256'h4c04510443042504f303c303a4039e03a303c303ea031804500476049804b704;
    decBuf[8860] = 256'hb2049804780449041104dc03ac038d0387039603ae03d403f8030f0435044404;
    decBuf[8861] = 256'h520446042304f003b203680336031a031203290359039103d40314043e046304;
    decBuf[8862] = 256'h6a04640448040f04cc037a0343031103070341038503c503ee03040419042c04;
    decBuf[8863] = 256'h3d042d040d04cd034403e202ac029c02ab02d302f7022e037403a203dc03f203;
    decBuf[8864] = 256'heb03cc038e033403f702aa028c0271028902af0208035d03aa03f003f903e003;
    decBuf[8865] = 256'hbb038b035f032103d702910251022802200243028702c702120344033a033203;
    decBuf[8866] = 256'hfe02ce029502610231021102f501e601eb010002230256029302cd0202030903;
    decBuf[8867] = 256'he902c2029402750258023f021e02f801d401d001ed0128027202a402ad029402;
    decBuf[8868] = 256'h6f024c022102f901cb01860146011d011601380157017f019801a601b301b701;
    decBuf[8869] = 256'hb3019d0184015d0139011001f300e400e900fe00210154018401b001cc01db01;
    decBuf[8870] = 256'hd601b0016e012e01f400ce00c800c100c700c200bd00ca00ed00160127011801;
    decBuf[8871] = 256'hdc0092004c001e000500fefff7fffdff030027004700650078007c0078007000;
    decBuf[8872] = 256'h630044001500e9ffcdffddff06002e0047004300360022002d00430057004500;
    decBuf[8873] = 256'h2100d4ff71ff49ff3dff48ff52ff49ff40ff48ff5dff7cff8dff92ff84ff66ff;
    decBuf[8874] = 256'h3cff09ffd9fea1fe8afe83fe96fec9fe14ff5aff88ffb1ffb9ffb2ff92ff6bff;
    decBuf[8875] = 256'h47ff27fff8feccfea5fe77fe58fe5dfe8bfec4fef8fe0dff06ffeafec6fea6fe;
    decBuf[8876] = 256'h88fe56fe0afec4fd72fd51fd6ffd9dfdd7fd0bfe2dfe4dfe5efe6dfe5ffe4afe;
    decBuf[8877] = 256'h27fe07fefafde6fddcfdc6fdc3fde0fd1afe75fe99fea4fe86fe6bfe52fe5afe;
    decBuf[8878] = 256'h61fe41feedfd98fd4bfd2dfd48fd72fd97fd83fd63fd47fd4cfd6dfd82fd76fd;
    decBuf[8879] = 256'h42fdfefcbefcb6fccdfcd4fce6fce1fce6fc06fd35fd7afda7fdb0fda8fda1fd;
    decBuf[8880] = 256'h9bfd8afd8ffd8bfd7efd63fd43fd2efd22fd3bfd6afd9afda0fd84fd4cfd08fd;
    decBuf[8881] = 256'hdafcf3fc0afd11fde5fc9cfc56fc28fc20fc45fc75fc88fc83fc73fc78fc8dfc;
    decBuf[8882] = 256'ha8fcb3fca9fca1fca3fcb9fcd8fce5fce9fce5fce9fc08fd37fd4afd39fd15fd;
    decBuf[8883] = 256'hf5fce8fc0bfd22fd1efdfbfcd1fcb5fcbafcbffcc3fc98fc5afc21fc19fc2efc;
    decBuf[8884] = 256'h41fc3bfc0dfce1fbc5fbd4fb10fc4afc70fc69fc63fc68fc8cfcacfccafcc6fc;
    decBuf[8885] = 256'ha7fc78fc65fc76fcaffcf2fc32fd4bfd34fd2dfd1bfd20fd3afd48fd2afdf0fc;
    decBuf[8886] = 256'h85fc3bfcf8fb04fc25fc43fc3afc21fcfcfb03fc2efc61fc76fc56fc0dfcc7fb;
    decBuf[8887] = 256'hacfbc5fbdbfbf0fbf6fbe5fbfffb44fcb2fc19fd41fd4efd2dfd23fd2cfd44fd;
    decBuf[8888] = 256'h3dfd0dfdc8fc9afc92fcb8fcf6fc1ffd26fd1ffd19fd1ffd24fd16fde7fc96fc;
    decBuf[8889] = 256'h33fcf0fbb4fba9fb9ffb95fb9efbc3fb0ffc55fc95fcbefcb6fca2fc9cfc8bfc;
    decBuf[8890] = 256'h90fc82fc75fc5afc50fc5ffc8afcdcfc3ffd9cfdf1fd12fef4fdd9fdc0fda9fd;
    decBuf[8891] = 256'ha3fd83fd3afde0fc8bfc80fc9efcdefc18fd1ffdeffcabfc8ffca8fcdcfcf1fc;
    decBuf[8892] = 256'hb9fc48fcf7fbcbfbf3fb48fcabfcb8fcc4fcb9fcd7fc3cfd99fdd6fdcbfd85fd;
    decBuf[8893] = 256'h57fd4ffd75fdc0fddefdd5fdbcfda6fdc8fd0dfe4dfe66fe31fee5fd8bfd67fd;
    decBuf[8894] = 256'h5cfd66fd5dfd44fd1ffdeffce8fcf9fc13fd21fd25fd29fd25fd28fd26fd28fd;
    decBuf[8895] = 256'h26fd28fd3afd54fd7bfda9fdc8fdeffd13fe3dfe6ffea0feb2feb8fea9fe91fe;
    decBuf[8896] = 256'h85fe81fe84fe8efe9cfe9ffe93fe80fe68fe58fe50fe43fe32fe12fedffdaffd;
    decBuf[8897] = 256'h9cfd8cfd91fd9ffd9afd96fda8fdd7fd22fe54fe70fe68fe33fe1efe25fe63fe;
    decBuf[8898] = 256'h9cfec2feadfe9afea0feedfe7cffdeff37000700bdff95ff89ffc0ffdeffb0ff;
    decBuf[8899] = 256'h55ffd0fe9afe8afef1fe34ff40ff1fffd9fed0fef9fe3dff6bff41ffd1fe3ffe;
    decBuf[8900] = 256'h04fe16fe67fecefedbfecffec4fee2fe34ffadff1f004b005900340029003300;
    decBuf[8901] = 256'h4f00680060003e00120001001b005700a100bf00c8009f006a0064006a007b00;
    decBuf[8902] = 256'h61001c00aeff64ff57ff7bffc8fffaff0300c9ff95ff9cffe0ff33006a006000;
    decBuf[8903] = 256'h2000e6fffcff4800b600e200d500b100bc00ee005201b001d4019d0143010601;
    decBuf[8904] = 256'h27018101a6019b014101d400c50008017501bf0196012901c2007f00a400f100;
    decBuf[8905] = 256'h23010701bd0063005700a400fe00530174015601280130016501b001f6010002;
    decBuf[8906] = 256'hd601a201a901d40129026502860254020202e101ff0151029e02a8025602f301;
    decBuf[8907] = 256'hb001bd010a02500259020e02b40178018301c9011b022602e0017c0153019001;
    decBuf[8908] = 256'hf30151025d022602f401eb014502b302fc020a03b50268027202c40227034f03;
    decBuf[8909] = 256'h4303f602b002b90203035d0369033203c4027b028802dd0214031e03cc026902;
    decBuf[8910] = 256'h41024d02b002f302e7029a0240021b023c02aa0211030403c70290027202d702;
    decBuf[8911] = 256'h4f03c103d00372031d03e60218037d03da03e6038303260301034e03bc032404;
    decBuf[8912] = 256'h1604c1035e0336035b03a803c60398031c039f028f02d90236038b0380032603;
    decBuf[8913] = 256'hd102c60220038d03d703ca0375031203040329038c03e903f603bf038d038303;
    decBuf[8914] = 256'had03ff0336042c04ec03b3039c03b103dc03ed03d403a10371036a039203ca03;
    decBuf[8915] = 256'hd203bd0378033803410366039603a9038d0355033e036003a503f7030204e403;
    decBuf[8916] = 256'ha4037b038303c103fa030204ed03b5038f039603cf03030418040504d203be03;
    decBuf[8917] = 256'hb703c803e203d4039d0359033e0336035b037e03840373035903420357037a03;
    decBuf[8918] = 256'h91039e0383034f033803310350038303b303c603b503a6039803ad03d003f003;
    decBuf[8919] = 256'hfd03da039e0364033f034603580375037a036303340321033d0376039b039403;
    decBuf[8920] = 256'h5c03fa029d0291029c02ce02d702be028a0275028802dc024903750383035e03;
    decBuf[8921] = 256'h110307031103290331030e03d602b102aa02c90212033003390331030c030503;
    decBuf[8922] = 256'h17031d03f902bd0262020d02ec010a02380251023a02fc01d301cc010a026402;
    decBuf[8923] = 256'h89027e023802e601c501cf012102580262023402fa01e40106023e0264026b02;
    decBuf[8924] = 256'h3f0223023202530270024e020802ae01a201c30109022402da014401d8009d00;
    decBuf[8925] = 256'hf7006801b2018a01ec00800045009f0031016c015a01c80066005400c5004a01;
    decBuf[8926] = 256'ha40173010c01ae00d2003501c8010302aa011801b600a400f5005c016a011501;
    decBuf[8927] = 256'h860024003500a70049015f01d60011005aff42ffafff11004600d5ff15ff92fe;
    decBuf[8928] = 256'haafe41ff19006f005500afff43ff57ffd4ff66007a00440091ff4aff34ffbeff;
    decBuf[8929] = 256'h5f009f006500e7ffb7ffe3ff5b00cd00a1000e005dff16ff2bff66ff9cff4bff;
    decBuf[8930] = 256'hc6fe49fe39fe82fefbfe2bffe2fe69fef8fd06fe7ffef0fefffebcfe1ffeb3fd;
    decBuf[8931] = 256'hc6fd43fed6fe10fffffeadfe64fe8cfef9fe60ff88ff64ff01ffd9fee5fe1cff;
    decBuf[8932] = 256'h62ff59fffefe79fe43fe33fe7cfebffe9bfe22fe90fd2efd3ffdb1fd18fe0bfe;
    decBuf[8933] = 256'hb6fd11fdcafce0fc42fdbffdf0fdc3fd30fdf5fc07fd79fd1bfe5cfe48feeffd;
    decBuf[8934] = 256'hbefdcdfd2bfe98fea7fe7efe11fec8fdbafdf7fd2efe4cfe1efee4fdbffdb8fd;
    decBuf[8935] = 256'hbefdadfd7ffd47fd13fdf0fcddfccdfca9fc7ffc58fc48fc5ffc7dfca0fccafc;
    decBuf[8936] = 256'hf1fc0bfd19fd0cfdf8fcf5fc0bfd30fd5efd7efd6dfd53fd45fd5afd95fdeffd;
    decBuf[8937] = 256'h14fe09feebfdbdfda4fdacfda5fd86fd53fdfafcbdfc9cfc7efc63fc4afc33fc;
    decBuf[8938] = 256'h3afc66fc82fc92fc84fc5dfc44fc48fc5efc69fc5ffc43fc2ffc33fc62fca0fc;
    decBuf[8939] = 256'hc9fceefc03fd22fd55fd85fdb1fdcdfddcfdd8fdbafd9ffd78fd54fd2bfd1afd;
    decBuf[8940] = 256'h00fde0fcc2fc9ffc9bfca7fcbbfcc5fcaffc84fc3ffc36fc60fc85fc7efc39fc;
    decBuf[8941] = 256'hd5fb92fb86fbe9fb61fcb3fca4fc97fc8afcd7fc59fdd7fde7fd9dfd25fdf4fc;
    decBuf[8942] = 256'h3efd9bfdf0fdcffd61fdfafcedfc5afdfcfd68fe2dfe8cfdf5fc93fcc8fc3afd;
    decBuf[8943] = 256'h66fd09fd6bfca9fb5afbd1fb68fcf2fc04fdb2fc4bfc3efc93fc22fd84fd72fd;
    decBuf[8944] = 256'he0fc56fc44fcd7fcaefd3efe24feadfd16fd2afdeefdd9fe77ff21ff36fe59fd;
    decBuf[8945] = 256'h02fd85fd5bfeb1fe2efe59fd8ffc75fc4bfd4efe71fe12fe0ffd1bfc3bfccafc;
    decBuf[8946] = 256'h81fdc8fd5cfd84fcf5fb77fc7dfd71fe90fe01fe4afd02fd6ffd6efe1cff3cff;
    decBuf[8947] = 256'hacfec1fda1fdf7fd17ffd7fffaff1cff53fe05fe4cfe0eff91ff4aff5cfe7ffd;
    decBuf[8948] = 256'heffc3dfd13fedcfec2fe1cfe84fd4afdc7fd9afef0fea2feccfdc9fca6fc45fd;
    decBuf[8949] = 256'h47fef6fed6fe46fec4fd0bfef9fe1500d5006d008fffc6fee0fe86ff1e003100;
    decBuf[8950] = 256'h6dff82fe23feb3fe9eff7b009800adffcffe79fefcfea2ffe3ff59ff4dfe8dfd;
    decBuf[8951] = 256'h6bfd09fe0bff74ff15ff4cfe32fe79fe67ff44006100aaff04ffc3fe25ffeaff;
    decBuf[8952] = 256'h6c008400edff63ff75ff2800fe0054013a019400fcffe9ff4200b400c3006500;
    decBuf[8953] = 256'hc7ff5bff48ffc5ff36004500e8ff4affdefef1fe6fffe0ff0d00afff2affd0fe;
    decBuf[8954] = 256'h01ffa3ff3b0075004000efffe0ff58000b01820197010e0191008100e8007b01;
    decBuf[8955] = 256'h0402cf013c018c004500b1003a0193014201a000ddffc3ff3a00d1000c01b300;
    decBuf[8956] = 256'he0ff50ff36ffdcff7300d500a000edff76ff8cff64002d01b001390176002800;
    decBuf[8957] = 256'h40002e014a02bd0255027701ae00c8009e01a1020903aa026e019c00c2007001;
    decBuf[8958] = 256'h4e026a02b401ae00baffdaffa3005a01a1010a01320069ffb7ff8d0056017001;
    decBuf[8959] = 256'hf9000c00adff3c005c011c023f02a001d700bd00630151022f0312035b028501;
    decBuf[8960] = 256'h6801eb019102fd02c302fe017b016401d00159026b02f9013901b700cf003b01;
    decBuf[8961] = 256'h76014001ae002400efff6000e5003f012e01c7008400a9004e01f40135022102;
    decBuf[8962] = 256'ha40173019f011802aa02be028802370228026b02d8023f034d03e0023d02fc01;
    decBuf[8963] = 256'he901420273022902b1011f01e40019016b0179016c01ff00b500a800fd004a01;
    decBuf[8964] = 256'h68012801bc0090009e002301a001f101e301ba01c7012a02bd02460358030703;
    decBuf[8965] = 256'h9f027702b4020103470319039e02200210025a029d02c1025e02cb0169015701;
    decBuf[8966] = 256'ha801d501ac01f7004000f8ff3900ea0061014b01e9006c007c003c012702c502;
    decBuf[8967] = 256'ha802bd011f010201ed010a037d035a037d02b401ce01d302c7036504d603b602;
    decBuf[8968] = 256'hf601d30172023b0355037f0209010a0039006001200242026501290056ffc9ff;
    decBuf[8969] = 256'h0301d601fc014e01f2ff67ff39009301d70202034202080189004901c902c803;
    decBuf[8970] = 256'hf6032403ca019c011a0227031b04fb03f902bf014001b401a8024603b6029701;
    decBuf[8971] = 256'h8a002100c00089010b0295017c006fff92ff300033019b013c013a008bffabff;
    decBuf[8972] = 256'hae00e801660240024b01ad000401230230039803390337028801e701b0029b03;
    decBuf[8973] = 256'hbb03f202070229014601c9019e028202cb019600c3ffeaff520030014d01ca00;
    decBuf[8974] = 256'hc5ff16ff75ff3e00f5003d01d00020007aff8fff67006a01d201b3015d01da00;
    decBuf[8975] = 256'h2101b9019002e702cd025602be018401dd016f02aa027402e2013201bb00d000;
    decBuf[8976] = 256'h5a01b3018201fe00390082ff6affabff0d001f00aeff29ffcffe00ff85ff4a00;
    decBuf[8977] = 256'hcc00b400740039002700990000015d016a0133010101f7004201b001f9012202;
    decBuf[8978] = 256'hfd01c601bc01c501de01c8016e01e9006c00faffceffdbffe7ffdcff96ff69ff;
    decBuf[8979] = 256'h50ff66ff89ff9bff8bff5cff18fffcfe05ff39ff69ff95ffa6ffbffffcff5600;
    decBuf[8980] = 256'hc3002b0153015f0154015e01790182017a014a01f900ac007a008300ac00d200;
    decBuf[8981] = 256'hbd006c001f00d9ffbdffc6ffbeff72fff0fe73fe43fe51feaffeecfee1fe87fe;
    decBuf[8982] = 256'h4afe55fed7fe9cff1e003600caff68ff56ffc8ff87000a01f2008600fdff3200;
    decBuf[8983] = 256'hc5009c01f301a401cf000500ebff6200ce00e200410028ff68fe45fee3fe73ff;
    decBuf[8984] = 256'h8dffe7fef9fd5bfdb1fd9cfe3aff1dff9bfec5fd6ffd26fe2bffd9ffbaff2aff;
    decBuf[8985] = 256'hdcfef3fee1ffbf004e01cc00f6ff66ffb5ffba0068018801bf00d3ff75ffcbff;
    decBuf[8986] = 256'h8200f8008c008dff53fe29fe9cfe4bffaaffe0fe8dfda5fccffcdcfdd0fe2fff;
    decBuf[8987] = 256'h9ffe7ffd0cfd75fd92fe9eff070029ff27febefd5cfe0b004001e901ea00a5ff;
    decBuf[8988] = 256'h27ff9aff19011802ea01c3001dff75fea8fe4900f100be001dff94fd61fdecfd;
    decBuf[8989] = 256'h13ff2000b7ff5bfe17fd98fc0bfdfffd9efe47fe90fdeafc00fdfffdf3fe91ff;
    decBuf[8990] = 256'h74ff26ffaffef0fea1ff4700880074001b000b0037007a009e00930061003400;
    decBuf[8991] = 256'h2b0042003b00f6ff80ff0effc4fe9cfe90fe59fefffdc2fda1fdd3fdeffdf7fd;
    decBuf[8992] = 256'hc2fd77fd59fd86fdf2fd76feacfebcfe90fe83fed7fe66ff17005e004900e7ff;
    decBuf[8993] = 256'hb1ffc1ff2800a100f200e300a0003300eafff7ff1b0052003400beff2bffc9fe;
    decBuf[8994] = 256'h94fe83fe92fe85fe30feb7fd86fd77fdd5fd12fe33fe15fee7fdbefdd4fd2efe;
    decBuf[8995] = 256'h83fed0fedafee3fe1cff8dff1f00810093006200360044009800270162012d01;
    decBuf[8996] = 256'h7a00d4ff93ffceff4b005b00f4ff2bff9bfe81fef8fe64ff78ffb3fe94fdd4fc;
    decBuf[8997] = 256'hf7fc95fd98febbfe1cfe53fd05fd7cfdc0fe05002f006fff7bfe1cfe1fff9e00;
    decBuf[8998] = 256'h9d01cc01a5004bffc0fee7ff8d01a6027302d10049ff16fffdff2401e4013601;
    decBuf[8999] = 256'h5bff7ffd42fd5afebfff4a00ccff26fe0dfddafcc2fd3dff70ffe5febefdfefc;
    decBuf[9000] = 256'h67fd84feddff0b008dffcdfe65fe42ff7e005101c401160138001b006a004001;
    decBuf[9001] = 256'hcf01b501df005000010019008500e700b2001f0096ff19ffe8fed9feccfec0fe;
    decBuf[9002] = 256'h89fe57fe29fe00fef9fd0dfe52feb6fef9fe05ffe4fedafe08ff73ff15005600;
    decBuf[9003] = 256'h4300e9ff98ffc4ff72004801d801be011701ab009800f10063017101f9002600;
    decBuf[9004] = 256'h96ffb0fff7ff6400290088ffc5fe43fe8afef6fe58ff22ffb1fe0efecefd08fe;
    decBuf[9005] = 256'h86fef7fe06ffdefed2fef3fe75fff2ff6400900068005c0067009900c6000001;
    decBuf[9006] = 256'h08010e01150126012b011401f600d300b3008c005e001900c7ff64ff21fffdfe;
    decBuf[9007] = 256'hf2fee8fedffec6feb0fea9fea3fea8fec2fef5fe25ff38ff1bffe3febefee0fe;
    decBuf[9008] = 256'h3effecff6200a30090007e006d00b7003001810190013201c5007b008800f600;
    decBuf[9009] = 256'h5d013501af00ebff9cff85fff1ff53001d008bffdafe34fe4afe85fe02fff1fe;
    decBuf[9010] = 256'ha8fe4afe0dfe70fe1eff95ffd6ff9bff1effedfe37ffe5ff8b00f700e400ae00;
    decBuf[9011] = 256'h7d00a90007017401a00178012301c0009800a400af00a50066000b00b6ff7fff;
    decBuf[9012] = 256'h61ff6aff83ffa8ffa1ff76ff21ff9cfe66fe56fea0fefdfe3aff19ffbffe82fe;
    decBuf[9013] = 256'ha3fe39fffcff7f0096002a00a1ffb3ff45001d01ad019301bd002d001300b900;
    decBuf[9014] = 256'h7c01fe01b701f5000900eaff4000f7000f01770051ff7efe0bfebafe58ffaeff;
    decBuf[9015] = 256'h60ffb9fe22fe0efeaffe72ffc0ffa8ff11ffaffec1fe74ff1a00b1009e002000;
    decBuf[9016] = 256'hcfffdeff56000901af01c50163010901b8008c00b400d800e3009d004b00feff;
    decBuf[9017] = 256'he0ffe9ff23003a001700baff41fff0fefffe42ff96ff8bff31ffacfe53fe63fe;
    decBuf[9018] = 256'he8fe65ffb6ff8aff47ff23ff70ff0600c800e2009b002f00f4ff4d002101ea01;
    decBuf[9019] = 256'h04028d01cb007c0094000001620150019e00c8ff38ff87fffdff69005600d9ff;
    decBuf[9020] = 256'h26ffaffec5fe27ffa4ffb4ff6bffd7fe75feabfe1dffa1fffbffcaff80ff73ff;
    decBuf[9021] = 256'hc8ff5700e0003a01e80064000a003b00a2001b016c012201c40070009100eb00;
    decBuf[9022] = 256'h3f014a01dc003a00ceffbafff0ff410050000d0088ff0bffdafe06ff64ff88ff;
    decBuf[9023] = 256'h67ff21ffe1fec9fe0cff83ffd4ffe3ffbbff96ffa1ff0f00b10049015c012701;
    decBuf[9024] = 256'h95005a006c00bd0024014c01f700940051008e00070158012c017e00a8ff52ff;
    decBuf[9025] = 256'ha1ff17008300490084ff99fe79fecffebbff59003c00b9ff13ffd2fe5cff2000;
    decBuf[9026] = 256'h6f00270065ffe2fefafebcffa80046012901a6005f007500fe007b018b010701;
    decBuf[9027] = 256'h6600faff0d008a00fc00ed00ab0056003500530093009b005700ceff45ff0fff;
    decBuf[9028] = 256'hfffe0eff1bfff7feecfe0aff4affa5fff9ff30004e0058007000780063002b00;
    decBuf[9029] = 256'he7ffccfff5ff5700cf0020011201cf00aa009f00e5003801590113018a000000;
    decBuf[9030] = 256'ha7ffb7ff1e0047002200bfff62ff3dffa0ff330095008400f1ff19ff8afea4fe;
    decBuf[9031] = 256'h1bffddfff7ffe0ff73ff39ff6eff2100c7000801cd002c00c0ffd4ff51000401;
    decBuf[9032] = 256'h4b010a01810027003800da009c01eb01a401b600d8ff82ff9cff13005400f2ff;
    decBuf[9033] = 256'h2dff76fe5efef6fef5ffa3008400f4ff3dfff6fe0bffbcff33004800e6ff45ff;
    decBuf[9034] = 256'h05ff67ff2b00e200590118018f00120022006c00c900d5009e003000e7fff4ff;
    decBuf[9035] = 256'h6100ab00ee00e200c1008f0085007d005800f1ff89ff11ff01ff0fff38ff44ff;
    decBuf[9036] = 256'h65ff6fff9cffe7ff190034000b00c7ff75ff54ff72ffa0ffb8ffcfffe4ff0f00;
    decBuf[9037] = 256'h6400e9001f014f015e015101450150013201bb00080062ff21ff5cffb5ff2700;
    decBuf[9038] = 256'h53002b00efffceff00002d003600f2ff69ffe0feaafedbfe42ffa0ffc4ffb9ff;
    decBuf[9039] = 256'h9bffb7fff0ff5200950089005200f8ffbbffc6ffe4ffffff29003f006f00b400;
    decBuf[9040] = 256'h180176019a016301f500710017000700f8ffebffc6ff63ff06fffafe5dfff0ff;
    decBuf[9041] = 256'h79008b00190095ff17ff07ff51ff94ffa0ff3dffdffea3fedafe70ff5e00fc00;
    decBuf[9042] = 256'h1801ca00b2009d00d8000d01fd00d1005800e7ffbaffe2ff37009a00c200cf00;
    decBuf[9043] = 256'hc400920052001800d4ffa7ff8eff96ff81ff55ff2eff14ff35ff74ffc6fffdff;
    decBuf[9044] = 256'hdfffb2ff89ff90ffc0ffdfffb8ff6bfff2fee2fe67ff2b00e20029011401b200;
    decBuf[9045] = 256'h7c00ee007301cc017b019d0081ff0eff76ff5400e300c90023000affe4fe4cff;
    decBuf[9046] = 256'h6900750153013600ddfef5fd1ffe2bff2000000037ff4cfeedfdb6fe0a00f100;
    decBuf[9047] = 256'h1c01a800b4ff55ffe5ff0501c4015c017e007cff59fff7ffc0004301fc003900;
    decBuf[9048] = 256'hb6ff9fff61004c016c011601f6ff36ff14ffb2ff41009000eafffcfe5efe41fe;
    decBuf[9049] = 256'hf8fecdff5d000f0069ffd1fe96fe13ffe7ff760091001a0082ff6fffc8ff7b00;
    decBuf[9050] = 256'h21013701d500580027007100040166015401a100cbff75ff8fff3600cd00e100;
    decBuf[9051] = 256'h40007dff2fff76ff0d006f003a0067ff9dfe4ffe96fe59ff1000f8ff8cffdbfe;
    decBuf[9052] = 256'hc3fe5bff3300fc004a01d400e6ff87ff6aff21009800d9009e002100cffffcff;
    decBuf[9053] = 256'h8f003f018701460195001e00ddff18004e007f003500d7ff6aff5bff9efff3ff;
    decBuf[9054] = 256'h1400e2ff90ff2dff05ff11ff48ff52ff37ff0dff06ff36ff94ff4200b800ce00;
    decBuf[9055] = 256'hba0085007500a100c900d500b4005a00edffc1ffe9ff5600bd001b010f01d800;
    decBuf[9056] = 256'h7e0072007d009b006d00f1ff50ffb9fea5fefffe50ff9aff8cff50ff45ff8bff;
    decBuf[9057] = 256'h140076008800160091ff38ff48ffafff0d001900f8ffdaff0800830024016501;
    decBuf[9058] = 256'h2a01ad003b000f0052008f00b0007e003e0014002b006900b300bd008f003500;
    decBuf[9059] = 256'he0ffa9ff77ff37ff0effd9feb7febdfef0fe3bff95ff02006a00ad00b9008200;
    decBuf[9060] = 256'h2800ebffcaffe8fff1ffe9ffc3ffafffdbff2f00cd00390174013e010d01e100;
    decBuf[9061] = 256'hee00ca0093002500a0ff23ff13ff5dffbaff0f001a00fcffe1ffc8ffdeff0100;
    decBuf[9062] = 256'hfbffdeff92ff45ff13ff09ff43ffa5ff02003f004a00680071008a00af00b600;
    decBuf[9063] = 256'h8a003600e1ffc0ffdeff4300bb00ec00dd009a0076009700f100460125018f00;
    decBuf[9064] = 256'ha1ff03ffe6fe00ff77ffb8ffa4ff4bff1aff64ff1100b800f9009600f6ff5eff;
    decBuf[9065] = 256'h23ff59ffcbff140007009aff50ff5efffbffbe0075018c012001be0089009900;
    decBuf[9066] = 256'he300f000b30024009bff65ffb7ff3b00950084001d00a5ff74ffa0fffeff3b00;
    decBuf[9067] = 256'h1a00acff44ff1cff71ffd4ff32002600efffa9ff9fffd9ff2c0063006d002d00;
    decBuf[9068] = 256'hd2ffaeffcfff3d00a400e700db00ba009c009300ab00d100ca0092003000d3ff;
    decBuf[9069] = 256'h96ffa1ffbfffdaffd2ffbcffa7ffbaffe1ff190030000e00d5ffa1ff9affb9ff;
    decBuf[9070] = 256'hcaffc5ffaeff90ff94ffc8ff1b00680072006900400047006900a200d600cf00;
    decBuf[9071] = 256'ha40066003c0026003b005a006b005b002800ebffa0ff82ff9effd7ff0c002100;
    decBuf[9072] = 256'h0100cfffacffb3ffe5ff23003c000700a0ff56ff64ffa0ff030046003a000300;
    decBuf[9073] = 256'hbdffb4ff0f009400ee00dd00b100530017002200680095009e005a001a00e1ff;
    decBuf[9074] = 256'hf7ff270046003600f3ff8fff66ff73ffc0ff1a0026000500abff56ff61ffbbff;
    decBuf[9075] = 256'h280072006400f7ff72ff3dff6efff2ff6f00a0005600f9ffbcff09009f003701;
    decBuf[9076] = 256'h710118016500efffaeff100069009a003300a0ff16ff04ff76ff180084007100;
    decBuf[9077] = 256'h1700a6ff79ffa2fff6ff2d002300d1ff6eff46ff6bffb8fffeff19000000dbff;
    decBuf[9078] = 256'he2ff0d0056008800a4008b0066005f006500810090008c007f00640044001e00;
    decBuf[9079] = 256'h0500e4ffcfffc3ffc0ffb6ffaeffa1ffb1ffd1ff04001900edffafff75ff5fff;
    decBuf[9080] = 256'h8fffc7ffdeffbbff77ff37ff60ffd0ff6300c500d70085003c0049008600d300;
    decBuf[9081] = 256'hf100b1003500b8ffa8ff0f006d00a90072001800c3ffceff000040003800d6ff;
    decBuf[9082] = 256'h5eff2dff3cff9affd6ffe1ffafff6fff67ffabff0f0037001300b0ff52ff46ff;
    decBuf[9083] = 256'h7dffebff350042003600150047009900fc0024011801cb00850058003f002800;
    decBuf[9084] = 256'h1400e8ffb5ffa1ffa7ffc3fff1ff04000a00faffe3ffc5ffa2ff79ff51ff38ff;
    decBuf[9085] = 256'h2aff2eff42ff61ff7fffa2ffb9ffdfff0d0045008900a4008c00570027001400;
    decBuf[9086] = 256'h3c007e00ac00b4008000420029004e008c00b60090002900a4ff6fff7fffc9ff;
    decBuf[9087] = 256'h0b00ffffb2ff58ff34ff6bffc5ff1a000f00b5ff2ffffafeeafe33ff91ffb5ff;
    decBuf[9088] = 256'h94ff76ff7fffcaff4c00c900fa000801c500890068008600b300bc0078002600;
    decBuf[9089] = 256'hd9ffcffffdff5700940073004100efffceffecff1a001100ceff69ff0cffcffe;
    decBuf[9090] = 256'hf0fe36ff64ff6cff47ff40ff52ff9cffe2ff0f001700100009001c0038004700;
    decBuf[9091] = 256'h39002d0031005e009600bc00a7006f003a0041008600c600ce008b000200a0ff;
    decBuf[9092] = 256'h8effbfff08003000f4ff91ff33ff27ff74ffcefff2ffbbff4dffe6febefefbfe;
    decBuf[9093] = 256'h5effa1ffc5ffbaffb0ffb9fff3ff45009200d800e100c9008500330012001c00;
    decBuf[9094] = 256'h5c0096008e004300e9ffdcff2900ab000501f5007000abff29ff70ffdcff1700;
    decBuf[9095] = 256'he1ff2eff88fe47fed1fe95ff4c0034009dff14ff02ff74ff3300b6006f00d7ff;
    decBuf[9096] = 256'h27ff0fffa6ff7e000e01280182001600dbff3400c600290117018400d4ff8dff;
    decBuf[9097] = 256'hcdff3000650075004900ecffafffa4ffc2ffddffc5ff81ff2ffff8feeefe1cff;
    decBuf[9098] = 256'h55ff7bff82ff88ffa4ffdcff20006000580032000200efff0b002f0046003a00;
    decBuf[9099] = 256'h0f0009002d007300e1000d01e5009000430011002c0034002d00fdffb8ff78ff;
    decBuf[9100] = 256'h70ff95ffb8ffd7ffd1ffb8ff97ff8bff8fff8bff82ff6eff6bff7cff9bffbcff;
    decBuf[9101] = 256'he2fffcff130042006d007e0079006b004d003a00300020002300300045006500;
    decBuf[9102] = 256'h7a0086007b006c005800550053003b000c00b3ff76ff3fff49ff77ff90ffa6ff;
    decBuf[9103] = 256'h9fff99ff9fffc3ffecfffdff0200ebffd6ffcaffc7ffcaffd2ffe5ff08004100;
    decBuf[9104] = 256'h66007b0075005900530074009a009f0076003800fefff6ff1900510068005300;
    decBuf[9105] = 256'h1b00e6ffd2fff1fff6ffe7ffb4ff76ff5eff74ff96ffb6ffbbffacffbafff1ff;
    decBuf[9106] = 256'h350062005a002500e8ffbeffd5ff050031002000f2ffdffffbff4800ab00d300;
    decBuf[9107] = 256'hc70090005e0055006e00750053000e00bcff85ff8fffbcffd5ffecffe5ffd2ff;
    decBuf[9108] = 256'he3ff1100300036000800c3ff95ff8dffa4ffd4ffe7ffd6ffbcffc1ffefff4100;
    decBuf[9109] = 256'h8e00ac00a300790045003e00440055005a00430025000a00070023004d006a00;
    decBuf[9110] = 256'h6f00580031000d00f6fff2ffdfffc6ffa4ff83ff88ffa3ffd0fffcff0d001200;
    decBuf[9111] = 256'h0d00230046005d0050001e00e0ffb6ffcdff0b0045004c0037000c001d005500;
    decBuf[9112] = 256'ha700de00e8009600490003000c0036003d001b00d6ff96ff9effd3ff2c005100;
    decBuf[9113] = 256'h46001400d4ffccfff1ff21002700f5ffa9ff77ff93ffddff37005b003a001c00;
    decBuf[9114] = 256'h13003c008000ad00b600810036000400faff340069007d006b0043001f002400;
    decBuf[9115] = 256'h39005c0061004b001100d8ffb2ffabffbeffe5fff5fff9ffe4ffe0ffebff1a00;
    decBuf[9116] = 256'h4a005c004c0028000700f2fff6ff00000400fbfff8ff090029006e008c009500;
    decBuf[9117] = 256'h7d0075008a009c00a2007e003900f3ffd7fff0ff2500470034000200d2ffcbff;
    decBuf[9118] = 256'h0900530071004400e9ffacffa1ffd3ff13001c00f6ffaaffa0ffceff29007e00;
    decBuf[9119] = 256'h9f006d001b00faff2c007e00b500ab0059000c00eeff09006400a000ab007900;
    decBuf[9120] = 256'h2700f0fffaff3a0063006b002d00e3ff9dff94ffbdff0f0030003a001f00e5ff;
    decBuf[9121] = 256'hcfffe3ff0f0036003c001b00e4ffbeffb8ffe3ff2c005e0068004f0038003100;
    decBuf[9122] = 256'h51008300a600ac00790049002a00300049006000540029000200f2ff09003800;
    decBuf[9123] = 256'h57003b000d00d5ffbeffd3ff0b0022001b00e3ffbdffb6ffd5ff080038003e00;
    decBuf[9124] = 256'h2200fefff1fffdff28005b0061004f00330023003100570085008c007b005700;
    decBuf[9125] = 256'h370021002500370040002c001400fefff6ff030018002c002a001e0013000900;
    decBuf[9126] = 256'h0100f8ffebffdbffd1ffcfffd7ffe9fff5fff7fff9ff02001700310049004d00;
    decBuf[9127] = 256'h4a0042003b003d0047004900440039002d0032003c0049004a00400033002500;
    decBuf[9128] = 256'h2300240020001200fbffdfffdbffedfffcff0500fdffe3ffd2ffceffe8ff0100;
    decBuf[9129] = 256'h17001400f7ffd4ffbdffd2fffdff2f0044004a002300fffffaff18004b006d00;
    decBuf[9130] = 256'h67003f00fdffe1ffeaff0f004d00660040001e00f2ffecff1000430058003900;
    decBuf[9131] = 256'h0600d6ffb7ffc7ffebfff9ffecffcaffb2ffaeffc9fff7ff16001c000c00f5ff;
    decBuf[9132] = 256'he8fff4ffffff0e0011000e000700010007001700260034004000410034001d00;
    decBuf[9133] = 256'h0700040012001d001b000500e0ffd1ffd5fffbff34004a002800f0ffcaffc3ff;
    decBuf[9134] = 256'he3ff0a001900f0ffa7ff75ff6bffa5ff07004a003d000600d4ffcbffe4ff1900;
    decBuf[9135] = 256'h3b0035000200b6ff98ffa2ffcbffffff2f00360030002100130028003b004600;
    decBuf[9136] = 256'h43002300ecffa8ff8dff85ffaaffdafffaffffffe6ffcfffcafff5ff28002e00;
    decBuf[9137] = 256'h1c00deff94ff76ff91ffcbffe1ffdaffbbff9fffaeffeaff24004a004300feff;
    decBuf[9138] = 256'hbeffa5ffcbfffbff1a00feffc6ffa0ffa7ffdfff320069004b000b00c1ffa3ff;
    decBuf[9139] = 256'hbefff8ff0e00faffb5ff75ff6dff92ffdeff10001900f0ffcaffb6ffbcffd8ff;
    decBuf[9140] = 256'he8ffd0ffaaff86ff82ff97ffbaffdaffdeffe2ffe6fffcff1b0031001d00f7ff;
    decBuf[9141] = 256'hc9ffa9ffbaffd4ffe2ffddffc2ffaaffb3ffdeff17003c002700fcffbeffa5ff;
    decBuf[9142] = 256'hbcffd0ffe3ffc7ff8eff69ff70ffa8ffddffffffecffc5ffabffb0ffd6ffe5ff;
    decBuf[9143] = 256'hd8ffa0ff7bff66ff92ffdbff0d000400dbffb5ffbcfff4ff29004b002c00d8ff;
    decBuf[9144] = 256'h83ff78ff96ffe8ff1f001500d5ff9bff85ffb5ff06003d003300f3ff88ff5cff;
    decBuf[9145] = 256'h4eff8bffc2ffe0ffc5ff7aff48ff64ffaeff08002c000b00b1ff75ff6affb0ff;
    decBuf[9146] = 256'hf0ff0800e3ff97ff65ff81ffcbff250049001200b8ff94ff9fffe5ff25003d00;
    decBuf[9147] = 256'hfaffa8ff71ff7bffbbfff4ff0b00f6ffb2ff84ff7cff92ffb5ffd4ffceffb5ff;
    decBuf[9148] = 256'h94ff7fff7bff94ffa9ffc9ffd6ffd2ffb2ff8cff87ff9effcdfff9fffeffdaff;
    decBuf[9149] = 256'ha8ff93ffa6ffe4ff1d002500f5ffbcff97ffacffd7ff0a000300d7ffa5ff90ff;
    decBuf[9150] = 256'ha3ffd5fff8ffe5ffbeff90ff89ffa5ffc9ffd7ffc2ff97ff7bff80ffb3ffd6ff;
    decBuf[9151] = 256'he8ffc1ff9dff8fff9cffbfffdfffe3ffc8ffb0ffadffbbffd8ffebffefffe5ff;
    decBuf[9152] = 256'hddffe5ffecfff2fff0ffddffcbffc3ffcaffd0ffd2ffc6ffb6ffabffb1ffbdff;
    decBuf[9153] = 256'hccffdaffd5ffbcffa4ff94ff9dffb4ffcaffd9ffccffb6ffa2ff9fffbaffe0ff;
    decBuf[9154] = 256'hfafffeffe9ffbeffa2ffb2ffd2fff8ff0800faffdcffc1ffc4ffe1ff03001100;
    decBuf[9155] = 256'h0500e9ffcaffbdffc9ffdaffe4ffe1ffceffc3ffc0ffcaffdaffe1ffdbffc7ff;
    decBuf[9156] = 256'hbaffb8ffbaffbcffc1ffc3ffc1ffc3ffc9ffd5ffe4ffeefff3ffeeffe4ffe0ff;
    decBuf[9157] = 256'hebfff8fffefff9ffe8ffd9ffd7ffddffefff04000700ffffeeffdfffd1ffd3ff;
    decBuf[9158] = 256'hdfffe6ffeaffe4ffdeffd7ffd3ffd6ffdfffeefff8fffafff2ffdeffccffc5ff;
    decBuf[9159] = 256'hd0ffdeffedfff4ffeeffe1ffddffe7fffcff100018000c00f9ffe6ffdfffe1ff;
    decBuf[9160] = 256'he7fff4fffcfffafffeff02000300000003000c0016001a000d00f5ffd6ffc9ff;
    decBuf[9161] = 256'hcdffecff0a0016000400eeffe6fff3ff1600300035001700f4ffddffeaff0c00;
    decBuf[9162] = 256'h1a0016000300f1fff4ff14003a003f0028000200deffecff12002c0027000100;
    decBuf[9163] = 256'hc9ffc1ffe3ff280056005e002a00ecffd3fff8ff3600600058001a00e0ffcaff;
    decBuf[9164] = 256'hecff25004a0043002400080003002c005400630039001200f8ff060024003f00;
    decBuf[9165] = 256'h35001200f2ffeeff11004300660053002000f0fff7ff13003700570042000f00;
    decBuf[9166] = 256'hdfffe5ff020030004f00550045002e0021002d0045004f005200450034003200;
    decBuf[9167] = 256'h3000320033003b003f0045004d004c004100320028001f002700320036002800;
    decBuf[9168] = 256'h18000e000c0018003000490052004a00420031002f0031003d0049004a004100;
    decBuf[9169] = 256'h33002a00320049005f0067006a005e0058005e00660068005d00490035003200;
    decBuf[9170] = 256'h430056005e004d0031001e0029004b0075007a0061002400fbfff4ff24005c00;
    decBuf[9171] = 256'h730050002400fdff02003e008900a7009d0064002f00280048008500af009800;
    decBuf[9172] = 256'h68003c002b0045008100aa00a300730054004300520072007f0064003e002400;
    decBuf[9173] = 256'h1f003d0060006e0050002d0016002b005e00800086005f003100120022005100;
    decBuf[9174] = 256'h7c008d00690040002f0048008500ae00b50093007400580067007e0093009700;
    decBuf[9175] = 256'h7f0063005f006900790087007a0060005500520061006e006700470026002200;
    decBuf[9176] = 256'h2e004d006b006f005d003b002d003a00650081009a0083005d0043003f005c00;
    decBuf[9177] = 256'h8f00b100ab008f006b00540069008c00b600b000960063004f00490065008900;
    decBuf[9178] = 256'h8d00780055003e004b005e0069005f0045002d00300044005c005f004b003300;
    decBuf[9179] = 256'h2a0044007100900096007200480038005b008e00b1009e007700530057007500;
    decBuf[9180] = 256'ha700bc00a900770054005b00770090008c006e004300320042006b007c006d00;
    decBuf[9181] = 256'h3a0018001e004500690080005a001700fcff040039007700a00089004c002200;
    decBuf[9182] = 256'h2a005a009f00ba00a1006d002f0027004c008a00b300ac007c0043002d004200;
    decBuf[9183] = 256'h6d0089007a00500029000f001400320045003b001f000300000010002f003c00;
    decBuf[9184] = 256'h30000a00fafff6ff14003e004f0035000c00f0ffffff290067007f0069003900;
    decBuf[9185] = 256'h0d0007002b005e0080007a00480017000500160039005a005e003b000800f4ff;
    decBuf[9186] = 256'hfaff160030002b000d00e3ffd2ffe1fff8ff16001a000100ecffe3fff5ff1400;
    decBuf[9187] = 256'h21001d00feffe8ffe4ff0400220035002b000e00f3fff0ff0c002f003d003000;
    decBuf[9188] = 256'h1500f5ffe9ffecff05001b0018000600f5ffe6ffe8fff4ff0600170019000b00;
    decBuf[9189] = 256'hf8ffebffedfff8ff0e00270032002900140007000a00210037004b004e003d00;
    decBuf[9190] = 256'h2a002200290038004e0057004f003e002f0025001d001e002c0031002c001f00;
    decBuf[9191] = 256'h12000000f9ff08001a002600240012000100fbff0100180027002a001d001100;
    decBuf[9192] = 256'h0f0025003f0050005400450033003f0056006c006f005c003e0031003c005500;
    decBuf[9193] = 256'h7100750055002f0016001a0038005300570034000100dfffd9ffeaff03001100;
    decBuf[9194] = 256'h0400e1ffcaffbeffc9ffe2fff1fffaffedffd7ffc9ffc6ffd2ffeafff9ff0200;
    decBuf[9195] = 256'hfffffdfff7fff1fffdff0f001f0026002800220017000d000e0017001f002a00;
    decBuf[9196] = 256'h2e0027001e0017000e000c0019002100220019000b00fbfff9fffbfffdfffeff;
    decBuf[9197] = 256'hfaffeeffe5ffe1ffe0ffd9ffcfffc3ffbeffbcffbeffbaffabff95ff7cff71ff;
    decBuf[9198] = 256'h81ff95ff97ff87ff67ff50ff43ff56ff6fff7fff70ff59ff43ff40ff52ff76ff;
    decBuf[9199] = 256'h8fff94ff87ff7cff7fff95ffafffc7ffcbffcdffd5ffe1fff4ff07000e001400;
    decBuf[9200] = 256'h1e002a003600430045003d00380034003d004700430038002a001b0010001200;
    decBuf[9201] = 256'h14000c000100efffdaffcbffbeffbcffbeffb8ffb3ffabffa0ff97ff90ff8bff;
    decBuf[9202] = 256'h8aff92ff99ff9cff95ff84ff73ff75ff7bff8eff9cff9eff8fff75ff6bff6eff;
    decBuf[9203] = 256'h76ff7eff7cff6dff4fff31ff1eff21ff2bff2eff1bff01ffe2feccfec1fec4fe;
    decBuf[9204] = 256'hc1feb3fea6fe8bfe7afe77fe7afe77fe75fe73fe71fe79fe81fe8cfe93fe8dfe;
    decBuf[9205] = 256'h87fe92fea5febdfed3fedcfed4fed6fed8feeafe09ff1eff32ff2eff1fff16ff;
    decBuf[9206] = 256'h19ff29ff3cff49ff47ff41ff33ff26ff28ff33ff34ff33ff2bff1cff04fffbfe;
    decBuf[9207] = 256'hf2fef0fee9fee7feddfed0fec5fec0febafeb6feb5feb2feadfeaefeaafe9efe;
    decBuf[9208] = 256'h96fe8ffe90fe9efeb8fec4fec0feb7feaefeb6fed5fefbfe15ff23ff16ff12ff;
    decBuf[9209] = 256'h1dff3fff72ff94ffa7ffadffbcffcafff0ff1e004a0050005f00640079009c00;
    decBuf[9210] = 256'hb300c800c400c100ca00de00f100fd00f600e000cc00c400cb00d200c800ad00;
    decBuf[9211] = 256'h8b006a0055004900460036001c00f6ffd2ffbbffaeffa2ff91ff81ff6dff56ff;
    decBuf[9212] = 256'h40ff37ff34ff32ff30ff32ff34ff2fff2aff23ff22ff26ff35ff43ff49ff4bff;
    decBuf[9213] = 256'h46ff3fff48ff56ff66ff6cff66ff5aff4bff39ff32ff34ff32ff26ff1bff04ff;
    decBuf[9214] = 256'he2fed4fec7feb4fea9fe94fe6efe55fe2bfe1afe0bfeeafdcdfdb1fd8bfd71fd;
    decBuf[9215] = 256'h63fd4efd33fd1bfdf2fcd6fcc6fcb9fca3fc88fc62fc3efc1dfc11fc15fc18fc;
    decBuf[9216] = 256'h02fcddfbaffb8ffb8afb99fbb0fbacfb99fb72fb59fb54fb69fb8cfba3fba7fb;
    decBuf[9217] = 256'ha4fba0fbb0fbd5fb0dfc33fc63fc76fc87fcb5fce1fc1efd69fd9bfdb6fdf0fd;
    decBuf[9218] = 256'h15fe61fea7fef9fe1aff4cff7affa3ffe6ff2600600086009a00ad00c900f700;
    decBuf[9219] = 256'h2f0155016a0163015e016d018401a201b501b901a30189017f0188019601a301;
    decBuf[9220] = 256'h98017c0169015e015b0169016c016001550147013f01470157015e0164016901;
    decBuf[9221] = 256'h71018801a401b701d701ec01ff012602540273029a02be02df0205033d036303;
    decBuf[9222] = 256'ha103da03000430045c048304bc04f00412053e055a056a0581059f05ba05d905;
    decBuf[9223] = 256'hee05f205ef05ec05f405fc050306f405e605cc05b105a705aa05960583056e05;
    decBuf[9224] = 256'h540549054d054f055d055f0554055e0575059705ca05fa051a06360664069c06;
    decBuf[9225] = 256'hef0652079507e90720086608b9081c097909ce091b0a610a8f0ac80a0c0b4c0b;
    decBuf[9226] = 256'h860bab0bc00bc60bcc0bd10bdf0bd20bb70b890b510b0d0bce0a940a500afe09;
    decBuf[9227] = 256'h9b095809eb08a1084408ef078c074907dc0692064f06fa05ad057b052905f204;
    decBuf[9228] = 256'hc00493047a047204500431041504f103da03d503ca03b80390035d032d030103;
    decBuf[9229] = 256'hcf029e0266020502a7015201d9008800030086fff4fe43fe9dfd06fd55fcaffb;
    decBuf[9230] = 256'hecfa35fa5ff9d0f819f873f7b0f6f9f553f5bbf432f491f325f39cf21ff2cdf1;
    decBuf[9231] = 256'h66f123f1fff0def0acf090f078f070f085f0a4f0c0f0e4f0f2f007f13af16af1;
    decBuf[9232] = 256'h95f1d3f1ecf103f233f239f255f279f27ef279f275f241f21bf215f2e9f1b6f1;
    decBuf[9233] = 256'h86f128f1cbf08ef041f0fbefbbef50efe9eea6ee39eeefedaced6fed22edf0ec;
    decBuf[9234] = 256'h9eec67ec49ec40ec38ec3fec2bec31ec4dec71eca4ecf0ec36ed63edadedf3ed;
    decBuf[9235] = 256'h46eebfee30ef98eff5ef4af0adf025f197f1fef177f2c8f212f36ff3c4f311f4;
    decBuf[9236] = 256'h7ff4acf4eef42bf54cf57ef5bef5e7f50df63df643f649f681f698f6acf6d8f6;
    decBuf[9237] = 256'hdef6cef6eff6fbf60ff73cf736f725f72af713f706f721f709f7e7f6cff690f6;
    decBuf[9238] = 256'h50f627f6d4f587f52df5a8f407f49bf3eaf244f2acf1d5f00bf020ef43ee40ed;
    decBuf[9239] = 256'h4cec6feb6cea78e95be89be7a7e6cae500e54ae4a3e30ce3aae274e264e255e2;
    decBuf[9240] = 256'h7de2eae252e300e405e53fe666e70ce995eac6ecd1ee35f119f4d2f64bf92ffc;
    decBuf[9241] = 256'haffff902f8053e0a170db710f214cb176a1ba61f7e221e266929422dd92f2333;
    decBuf[9242] = 256'h4735ff37793ab83cc43e1840c841e142e043c7444645b945964576455a45d744;
    decBuf[9243] = 256'h31446e434f428f415540da3edb3d3a3cb13ab239103887368835e733ce32cf31;
    decBuf[9244] = 256'h8b30642fa42ef62d182dc22c3f2cc92bb32b9f2b8e2bbe2beb2bf82b652caf2c;
    decBuf[9245] = 256'hf22c772df42d452eca2e242f752fbf2f01300e302f301130d12f862f042f642e;
    decBuf[9246] = 256'ha12d822c752b3b2ac028f52645254c237021c81e4f1c0f1a6e17f5141112580f;
    decBuf[9247] = 256'h2a0c2b09ac05610262ffaafc7bf97df6c4f34bf167eeaeebeae9aae79fe54be4;
    decBuf[9248] = 256'h9ae282e183e0f8df79df06df29df49dfd8dfc4e0a1e117e37ce41de616e8f2e9;
    decBuf[9249] = 256'h99ec13ef53f1f3f36df6adf84dfbc7fd07001202760411061c08f809a90bc10c;
    decBuf[9250] = 256'hc00da80e7b0fee0f1110f10f9b0f180f430e400d060c8b0a260984078b05af03;
    decBuf[9251] = 256'h840178ff14fd79fb6ef90af76ff563f387f1d7ef4eeee9eca5eb29ea2ae943e8;
    decBuf[9252] = 256'h70e7b0e602e6a3e54de532e51be505e540e552e5a3e5ede530e66ce6a3e6c1e6;
    decBuf[9253] = 256'hcae6f4e6dde6c9e6a9e660e606e6b1e54ee5f1e484e4ffe382e3efe266e2e9e1;
    decBuf[9254] = 256'h77e1d5e03ee0b4df37dfc5de5edee6dd94dd68dd40dd4cdd83ddc9dd2edec1de;
    decBuf[9255] = 256'h71df18e0dae0c5e163e266e315e4f2e4bbe5a6e644e747e8f6e894e996ea45eb;
    decBuf[9256] = 256'h22ecebeca2ed49ee36ef95ef25f0a8f0eff005f167f131f141f150f10df1d1f0;
    decBuf[9257] = 256'hdcf06ef024f016f079ef0defabeec2ede5ec55ec01eb60e947e87ce651e445e2;
    decBuf[9258] = 256'he1dfa2dd01dbd2d7d4d41bd2edce13cb74c729c450c0b0bc66b98cb5edb1b1ad;
    decBuf[9259] = 256'hd9aa39a7eea3f0a0379e739c339abd9879983c987498d999d79b3b9e1fa166a5;
    decBuf[9260] = 256'h62a913af61b495ba15c225c966d12ad93ee2c9eac5f42afeb506b110c51ce524;
    decBuf[9261] = 256'h3b2fa0389b43fd4a63547d5a41624c67b76de271ac751e79ff7a907b157c9c7b;
    decBuf[9262] = 256'h2f7b3d79c4763b73006f046b52650460d159fb53a54b1946093fc9363d312d2a;
    decBuf[9263] = 256'hc223ec1d9e18cb136a0f6d0bd7087d0634050a046404b7040105dd060909aa0b;
    decBuf[9264] = 256'hd80ed7111d161a1ac21e24234428162d783198360a3a6b3e6842fe445847a148;
    decBuf[9265] = 256'hcb4971497a480447a0441741dc3cbc37ea32072c9c251b1e07157c0cb804a0f9;
    decBuf[9266] = 256'h4aefe4e55add5ed3f8c96ec1aab99ab259aa95a2859bf0961a91cc8b5a883985;
    decBuf[9267] = 256'h8483f6818d80fa802582e983ce864d8a898ea8937b985e9fc9a5f4ae7fb743bf;
    decBuf[9268] = 256'h57c852d3a8dd0ee709f25ffcc405c010161b7b24062dca34de3df843bc4bc750;
    decBuf[9269] = 256'h32575d5bab601d643e67176aa56b1d6c8b6c276c636ac768916593624c5e505a;
    decBuf[9270] = 256'ha7550550b74ae4454240783c45361a32502e7d291c254322a31e491c4b195917;
    decBuf[9271] = 256'h9515fa131913d512981240133f148415a717481ac21c4a2095239326da2ab32d;
    decBuf[9272] = 256'h5231ac33ab369c38613a573b383c7c3c3e3c253bc0391f38b535d132522f162b;
    decBuf[9273] = 256'h1a277222cf1c81174e11ce09be0253fcd2f4c2ed82e5beddaed643d06dcaa3c6;
    decBuf[9274] = 256'hd0c16fbd96ba08b99fb70db870b880b9c0bb60be8fc168c511cab3cf01d595dc;
    decBuf[9275] = 256'ha5e3e6ebaaf3befc4905450faa18a523072b6d34f73cbb44cb4b61503656005a;
    decBuf[9276] = 256'h725d94604962cd624663fd61d3600e5f2a5caa586f544f4f7d4a9a432f3dae35;
    decBuf[9277] = 256'h9a2c8026841c1f13940ad002c0fb55f5d5edcae85ee233de69da58d878d6c2d4;
    decBuf[9278] = 256'h3ed4c5d333d45dd522d762d96ddbe1de2ce205e6aeea50f09ef5d1fba701f506;
    decBuf[9279] = 256'h280dfe124c181e1d40203c24d2263c28a928462836279b2590231c20d11c1c18;
    decBuf[9280] = 256'hbb139b0e68089202c0fb7ff3bbebabe46bdc6fd209c97fc0bbb8a6af1ca7589f;
    decBuf[9281] = 256'h4898b293dd8d8f881d853c83878102818a80d281c4833d86c689118dc5916897;
    decBuf[9282] = 256'hb69ce9a269aa79b1bab97ec192ca1dd319dd7ee609ef05f96a02840848105315;
    decBuf[9283] = 256'hbe1be91f2f22a1254126d3264f26d625b323c121481fbf1b84178713d60d8808;
    decBuf[9284] = 256'h55027ffc29f465ec55e514dd50d53ccc22c65ebe4fb7b9b2e3ac19a9a7a586a2;
    decBuf[9285] = 256'hd1a0439fcb9e5d9efa9d549e4b9f969feaa0a3a1bca221a465a5e1a6aca85caa;
    decBuf[9286] = 256'h55acb9ae54b0cab1a6b35fb497b4cab4e2b3bcb27cb098addfaab1a7d7a338a0;
    decBuf[9287] = 256'hfc9b00986a951f92fb8fd18e0c8dba8c058dd18d068f6f91af93e596bf9a5e9e;
    decBuf[9288] = 256'h8aa3bea93eb14eb88ec08aca9fd6fee148efcbfb2a077414f62016296c33d13c;
    decBuf[9289] = 256'h5c45204d2b5296586c5eba638c682f6ef9716b758c78657bf27c5b7ec97e2c7f;
    decBuf[9290] = 256'h1d7e817c767a0277c772cb6e1969cb63985dc2577452414c6b461d414a3ce937;
    decBuf[9291] = 256'hec334d30022d042a4b27872547233c21e81fb31e9a1d011d8d1d0b1e181fdd20;
    decBuf[9292] = 256'h0923a925d828d62b8f2e723209356337613a533c623d593ea43e603ea73d8e3c;
    decBuf[9293] = 256'hc33a9738f635c832c92f4a2c0f2812246a1fc8197a14e50cd6056affeaf7d6ee;
    decBuf[9294] = 256'h4be687de73d5e8cc24c515bea9b7d4b186ac52a627a25d9e4c9c2b997697e895;
    decBuf[9295] = 256'h709502956695c0955c976799539cd29f0ea451aa27b0f9b664bd8fc61acfded6;
    decBuf[9296] = 256'hf2df7de879f22ff9b9017d098d10ce185a1e6a25d52baa317c38123de842b246;
    decBuf[9297] = 256'h844ba64ea2522f548956f7565a57005765555953f5506d4d224a4846a9426e3e;
    decBuf[9298] = 256'h713ad2368733ae2f0e2cc428c5254622fb1e211b821737143911b90d5f0b6108;
    decBuf[9299] = 256'h6f06ab04b40369032503df038704ec053107ac08770a270c400da50ee90f1011;
    decBuf[9300] = 256'hd0117e12dd126d13f0136614d314351547159815a71599157515d0149b132012;
    decBuf[9301] = 256'hef0fe40df80a3f085c04bc0072fd98f9f9f59ff3a0f0e8ed6eeb2ee9b9e765e6;
    decBuf[9302] = 256'h30e5a7e3a8e207e15ee05fdf31dfb3de8cdeafde4ddfc3e08ee235e5afe793ea;
    decBuf[9303] = 256'h12ee5df112f673fa70fe0f025a053309d30c1d101c13d4154e18321b241d5220;
    decBuf[9304] = 256'h76222e25a82743294e2ba22c522efb2e942f092f362edd2c3b2b42296627bf24;
    decBuf[9305] = 256'h90216d1fb41c3b1a57179e142512e50f440dcb0a8b08ea0571038c00d4fda5fa;
    decBuf[9306] = 256'h82f8c9f550f310f16feeabecb4ebd4ea08eacae992e95fe9eae968ea8feaf7ea;
    decBuf[9307] = 256'h17eb34eb4eeb36eb4ceb5feb4eeb5eeb8aebcdeb52eccfec21ed88edcbedefed;
    decBuf[9308] = 256'h26eef4ed6bed93ec91eb11ea12e971e778e59ce3ebe1f2df9edeeedc65db00da;
    decBuf[9309] = 256'hbbd895d788d694d5b6d4edd302d325d25bd1a5d02ed018d005d05ed0f0d0c8d1;
    decBuf[9310] = 256'h3ed309d5b9d622d962db03de7ce061e319e693e877eb68ede2ef22f2c2f487f6;
    decBuf[9311] = 256'hc7f8d2fa26fc52fec7ff9300c801e10214039f03750302035302370191ff08fe;
    decBuf[9312] = 256'hd7fb36f971f78df4d5f15bef77ecbee945e705e564e2ebdfabdd0adb46d906d7;
    decBuf[9313] = 256'hfbd4a7d37bd170cf1ccee7cc5ecb5fca1bc948c888c7dac63cc6acc5c1c4e3c3;
    decBuf[9314] = 256'h54c369c28bc188c04fbfd3bd6ebccdba44b979b7c9b540b40fb299b0bdae89ad;
    decBuf[9315] = 256'h00ac01abbca9e9a8c3a85aa8b9a883a939aa9eab69ad10b03eb318b7b7bae4bf;
    decBuf[9316] = 256'hb6c458ca2ad196d716df26e667ee2bf63afd5107b61041190521192aa3329f3c;
    decBuf[9317] = 256'h5643e04ba453b45a4a5f1f656d6a406f61723a75d0773a79827ae67a8b7a9479;
    decBuf[9318] = 256'h897725759c71526e786ad0656e612b5b55550750344b92454440723bcf350532;
    decBuf[9319] = 256'h332dd128f8255922ff1fdb1db11ca11b4f1b041b481b021caa1c0f1e6a20aa22;
    decBuf[9320] = 256'h4a25c4274d2b972e963115356038393cd03e2a414d433f454e46454790474c47;
    decBuf[9321] = 256'h17468e445d42bc3f8e3cb4380c34aa2f8a2a5724d71ccb178b0fc707b70076f8;
    decBuf[9322] = 256'h7aeec4e739df3dd5d8cbbec5c2bb0cb5f2ae2ea723a28d9d6299989526924690;
    decBuf[9323] = 256'h908e0c8e848ef28ee390a8928c95d299f29ec5a3a8aa13b193b8a7c132ca2ed4;
    decBuf[9324] = 256'h93dd8fe8e5f24afcd504d10e3618c120bd2a22343c3a004210497b4f51559f5a;
    decBuf[9325] = 256'h715fd363cf67666ac06c2d6d916d366d3f6c346a4867c9638d5f915be9564651;
    decBuf[9326] = 256'hf84b26478341353c02362c30de2a0c26aa218a1cb81756135a0fb10a90079403;
    decBuf[9327] = 256'hfd00a3fe80fc55fbfbfa04fa4ffa93fa4cfbd5fc3afe7fff4e01fe0287045206;
    decBuf[9328] = 256'h87071009750a5d0b2f0cef0c9d0dfc0d530e380e210ee00d560db60cc80b6c0a;
    decBuf[9329] = 256'hca08d106f5044e02d5fff0fc71f926f628f36ff0f6edb6eb15e951e7b5e540e4;
    decBuf[9330] = 256'h74e3bae282e2e9e1bbe1e5e158e2c1e29ee367e4bbe55ce756e9baebf9ed30f1;
    decBuf[9331] = 256'h2ef4e7f6cafa6afeb401b30432087d0b7b0e3411ad13ed15f817d419851b9d1c;
    decBuf[9332] = 256'h021eea1e1120842032219121e8210222ea21a921d120ce1f951e191db41bb619;
    decBuf[9333] = 256'hda17af15a313c71117108e0e290d880bff090009bb0794063b05f603d002c301;
    decBuf[9334] = 256'h8900b6ffaafe70fd9dfc91fb57fa84f9c4f8d0f732f769f6e6f56ff503f553f4;
    decBuf[9335] = 256'hdcf3eef211f2d4f0aeef07ee7fecb4ea88e87de629e5fde287e1abdf7fdd0adc;
    decBuf[9336] = 256'hb6da05d97cd7b1d501d408d2b4d004cf7bcdb0cb7bcaf2c8f3c70bc739c6c6c5;
    decBuf[9337] = 256'he9c508c698c64fc7b3c818cab9cbb3cd8fcf36d2afd4efd690d909dceede6de2;
    decBuf[9338] = 256'hb8e5b6e836ec80ef7ff2c5f69ef93efd880087033f066e09910b830d470fe210;
    decBuf[9339] = 256'hc311071244120c120d118210070f3c0d8c0b9309b7078b05ea02bcff98fd19fa;
    decBuf[9340] = 256'hcef6d0f389ef8debf6e8bbe4bfe028dededadfd727d5add212d107cfb3cd02cc;
    decBuf[9341] = 256'heacaebc903c984c811c8a9c74ac7f4c671c62ac6bec55bc5bbc423c473c3fcc2;
    decBuf[9342] = 256'h64c2b4c10ec14bc060bf43be37bdb7bbecb93cb843b6dfb343b2ceb0f2aebdad;
    decBuf[9343] = 256'ha4aca5ab77abf5ab68ac5cadf8ae80b017b346b61fbabfbdebc21ec9f4ce42d4;
    decBuf[9344] = 256'hd6dbe6e227ebebf2faf91104c70ac2151820ce26ca31203c8545104ed455e35c;
    decBuf[9345] = 256'h4f632469726ee47146761f79ac7a067d4f7eb27e0d7fba7e457d697bc1789375;
    decBuf[9346] = 256'hb971116daf688f635c5d86573852054c2f46e140ae3ad8348a2fb82a56267d23;
    decBuf[9347] = 256'hde1f841d3b1c4a1aef199d19e819b41a6d1b151ce01d911ffa213a24db26092a;
    decBuf[9348] = 256'he32d8231bd35ba39593da440a24394450d480449e449284a6f49e64781462644;
    decBuf[9349] = 256'h4241c33d87396734952ff3292123b51c3515250ee40520fe11f7faec44e649db;
    decBuf[9350] = 256'he7d382caf7c1fbb745b1baa82ea31e9c89975e93948f838d618ad0894b89c489;
    decBuf[9351] = 256'h0c8bfe8c778f5b92db95169a59a02fa601ad6cb397bc22c5e6ccffd755e2baeb;
    decBuf[9352] = 256'h45f441fea607a212041a6923f42b80318f38fb3ed0441e4af14e53534f57e559;
    decBuf[9353] = 256'h3f5c635ec65e215fce5e595d7d5bd558f2545251264c5447b141633c30360532;
    decBuf[9354] = 256'h332b9d26c8207a1ba7164512490eaa0a6e067202d3fe88fb89f8d1f557f318f1;
    decBuf[9355] = 256'ha2efd6ee1dee55eeeeeed6ef51f1b6f2b4f490f640f839fa15fc4afdd3fe3800;
    decBuf[9356] = 256'h7d014f020f037803160433044d0464042404c1038c03fa0297021a022701edff;
    decBuf[9357] = 256'h72fea7fc7bfadaf761f57cf2c4ef4aed0bebffe8abe7f2e64ae617e645e66fe6;
    decBuf[9358] = 256'h2fe7dde77ce80be98ee964eaa0eb1bede6ee12f11df381f565f8e5fb2fff0903;
    decBuf[9359] = 256'ha806f309cd0d6c11a7158018201c7a1e78216a23e3257e275f282b29e4291c2a;
    decBuf[9360] = 256'hb52a402b132c392c5c2c7c2c252ca32bcd2a572926271b252f22761f481c241a;
    decBuf[9361] = 256'ha5164b1428126f0fab0d0f0c9a0abe08890700069b0456032f02d60035ff1cfe;
    decBuf[9362] = 256'hb7fccffba8fae8f93af95df806f8ecf704f845f8a7f800f972f9f7f92dfa3dfa;
    decBuf[9363] = 256'hf3f945f96ff833f7b8f553f4b2f229f1c4ef22ee0aeda5ebbdea42e943e8fee6;
    decBuf[9364] = 256'h2fe57fe3f6e1c5dfb9dd55db16d975d6b0d471d2fbd0a7cf72cecacd97cd68cd;
    decBuf[9365] = 256'h93cd06ceb4ced1cf91d0cad1f1d2fed37ed5e3d684d87ddae1dc21dfc2e13be4;
    decBuf[9366] = 256'h1fe79feae9edc3f162f5adf8acfb2bff760299048b060409fb09710b3d0cf60c;
    decBuf[9367] = 256'h9e0dd10da30dcd0da70d3e0da00cd70b4f0a56087a06d203a400a5fd5ff963f5;
    decBuf[9368] = 256'hc3f188ed8ce9ece5a1e2c8de28dbded7dfd427d2adcfc9ccd8ca5ec8c3c64dc5;
    decBuf[9369] = 256'h71c33cc224c125c03dbf13bfa0be7dbe1bbfabbf96c0f2c136c306c5b6c6cec7;
    decBuf[9370] = 256'h33c91bca45ca6cca49caabc91bc998c822c88ac7dac633c69cc5c4c4c1c388c2;
    decBuf[9371] = 256'h0cc141bf91bd98bb44ba94b87bb77cb64eb6cfb5f6b5a4b642b745b80aba36bc;
    decBuf[9372] = 256'h6cbf46c3eec750cc93d269d83bdf7ce708ed18f458fc1c042c0b6d13311b4524;
    decBuf[9373] = 256'hd02ccc363140bc4880508f57d05f5c65676afd6e2873f2760379e47a997c277e;
    decBuf[9374] = 256'h9f7e0d7fe27d1e7cde7912767372466d7468d262845db158ce51384d63471542;
    decBuf[9375] = 256'he13b0c36be308a2a60261221a01d3e196516d8146f1326128a12e41292127213;
    decBuf[9376] = 256'h3e14f71480164b18fb19d51c8e1fbc229626352a802d5931f0333a375e39883a;
    decBuf[9377] = 256'h4d3c9f3c543c103cdc3a5339ee379335af322f2ff42ad42501215f1b8d14220e;
    decBuf[9378] = 256'h4c08f6ff32f822f1e2e81ee109d87fcfbbc7abc06ab8a6b09bab30a55a9f909b;
    decBuf[9379] = 256'h1e98bd9307927a90118f7e8f1b8f2a90c59166949597499caba0eea66fae7eb5;
    decBuf[9380] = 256'hbfbd83c59cd0fed763e15fecb5f61a00a508a112061c9124552c6935833b4743;
    decBuf[9381] = 256'h564aec4ec254105a825da3607c63096572660566a1659264ae61f55e125b6956;
    decBuf[9382] = 256'hc750794b4545703f223aee33192ecb289722c21c7417a112ff0c35096204c0fe;
    decBuf[9383] = 256'hf6fa23f602f329f093ed39ebf1e954eafae9f0ea66ecbaedefee58f1f3f2fff4;
    decBuf[9384] = 256'h63f7a2f9aefb12fef600e7026105a107ac09100cab0d210f75102e114712e012;
    decBuf[9385] = 256'hc813461406156f154f15bf14a013fa1101109d0d5d0bbc084306a7043203de01;
    decBuf[9386] = 256'h24017c0049001b009cff76ff82fe65fd0cfcc7faf4f9cef9abf949fa4cfb86fc;
    decBuf[9387] = 256'h01feccfff8010304df058f078809640b900d9b0fff113f144a162618521a5d1c;
    decBuf[9388] = 256'hb11de61eff1f98208021fb22fa239b25b426b3279b28c229352a582ab929b728;
    decBuf[9389] = 256'h37276c25bc2333226820b81e2f1dca1b851ab319f318b9173e16d91437133e11;
    decBuf[9390] = 256'h620f360d2b0b4f09230718053c038c01030038fe88fc6ffb70fa88f9b6f8f6f7;
    decBuf[9391] = 256'h02f724f65bf53cf4e2f29ef17aef6fed93eb67e95ce708e658e4cfe2d0e1e8e0;
    decBuf[9392] = 256'h15e055df1bdef5dc9bdb57dadbd876d732d6b7d4b8d373d2a0d1e1d078d058d0;
    decBuf[9393] = 256'h02d050d0c7d08ad1a9d24fd4d8d5a3d7cfd9dadb3eded9df4fe12be3dbe4f4e5;
    decBuf[9394] = 256'hbfe7ebe9f6eb5aee3ef1f7f325f724fadcfca1fee1005602aa03df048705ba05;
    decBuf[9395] = 256'h46061b0642061f06c0053005790474033a021301baff19fe00fd9bfbfaf971f8;
    decBuf[9396] = 256'ha6f67af4d9f1abeeaceb2de8e2e409e172de18dc1ad9efd72bd634d5bed3f2d2;
    decBuf[9397] = 256'hbed135d0d0ce2ecda5cb40cafcc829c869c701c720c73dc78bc702c843c8ccc8;
    decBuf[9398] = 256'hb5c992ca95cb15cd14ce58cfd3d038d220d39fd378d310d371d235d10ed002cf;
    decBuf[9399] = 256'h0ece6fcd19cdcbcc84cc43cc6bcb68caa3c877c6d6c3a8c0a9bdf1ba77b837b6;
    decBuf[9400] = 256'hc2b46eb339b271b23eb26cb293b353b4d3b504b8a5bad3bdadc155c6f7cbc9d2;
    decBuf[9401] = 256'h35d90adfdce547ecc8f3d8fa1803dc0af113ec1e4229a732a33d05456a4ef556;
    decBuf[9402] = 256'h815c90632668516c976e09722a75df767679d07b187d437e527f007f207ebc7b;
    decBuf[9403] = 256'h7c79b0750871a66c63668d603f5b0c55364fe849b543df3d0d37a230772c2927;
    decBuf[9404] = 256'h5622f51d1c1b7c171316f013c512b6116411ee0f3210f40fbc0fbb10a3117213;
    decBuf[9405] = 256'h191693181c1c57205324f3273d2b172fad31073450357a368a37383757368b35;
    decBuf[9406] = 256'h5734ce3203315b2ee22b59281e2445219d1cfa16ac11790ba305d1fe91f6cdee;
    decBuf[9407] = 256'hbde77cdfb8d7a4ce8ac8c6c0bbbb4fb57aaf2caabaa699a3c0a0299ec09c9d9a;
    decBuf[9408] = 256'h399a949ae69ac69ba29d539f9ca2e7a59caa3eb010b77bbdfbc410ce9ad65ede;
    decBuf[9409] = 256'h73e7fdeff9f9af003a09fe100e184e20da25ea2c55332b39793eac44d748254e;
    decBuf[9410] = 256'h9751b8546e5604597d590f59ac58e756a7540752234e844a57458540233c0337;
    decBuf[9411] = 256'h31328e2cc428f223901f701afe169d127d0d0b0aa9058a0018fdb6f8baf423f2;
    decBuf[9412] = 256'hc9ef81ee56edfcec4eed2eeefaeeabf0a4f208f547f753f9b7fbf6fd97005c02;
    decBuf[9413] = 256'h9b043c07b609f50b010e65104913011630192e1cae1f08222b241d26e127d828;
    decBuf[9414] = 256'h2329df2826280d270e26c9244e23e921a5207e1f711ec31da61c4d1b4f197317;
    decBuf[9415] = 256'h4715a612e210fd0d450b160818055f0231ff0dfd1cfb57f9bcf746f602f649f5;
    decBuf[9416] = 256'h11f5aaf5d8f502f6c2f671f790f7e7f7ccf7b5f74cf824f99afa65fc90fe3101;
    decBuf[9417] = 256'hab038f060e0a590d58101013d51414178a18de19131b2b1cc41c501d221e491e;
    decBuf[9418] = 256'h6b1e4c1ef61d3f1dc81caf1b551a1119411716150a13a6101e0dd309fa055101;
    decBuf[9419] = 256'haffb61f68ef12ced30e991e546e248dfc8db6ed970d6b7d389d08acdd2caa3c7;
    decBuf[9420] = 256'ha5c425c1cbbe83bd58bcfebbacbbf6bb3abc78bc20bd85becabf99c14ac343c5;
    decBuf[9421] = 256'ha7c7e7c9f2cb56ce96d0a1d27dd42dd626d802dab2db1cde00e1b9e3e7e6e6e9;
    decBuf[9422] = 256'h9eec18efb3f029f26df2aaf2e2f215f3e7f211f338f3a0f3fff355f4a4f4bbf4;
    decBuf[9423] = 256'h4ff49ff3f8f2b4f1ccf0a5ef4cee64ed3dec7deb89eaace9a9e86fe748e6a2e4;
    decBuf[9424] = 256'h19e31ae232e160e086e063e001e191e1abe194e153e1a2e0ccdf3ddf86deb0dd;
    decBuf[9425] = 256'h5addd7dcbfdc00dd8add72de8fdf02e06ae0c9e039e0b7df11df23de85ddf5dc;
    decBuf[9426] = 256'h72dc5adc45dcbbdb62db31dbe8dadada17dbf6daecda07dbcddac6da12db1cdb;
    decBuf[9427] = 256'h49db51dbf0da78da26daa2d948d917d9ced8c0d8e5d8dad8e4d8c8d84dd888d7;
    decBuf[9428] = 256'h9dd641d559d4ded279d134d00dcf67cd4fcc84cad3c84bc780c5cfc346c247c1;
    decBuf[9429] = 256'hbcc092c0b9c021c13ec24ac3cac495c645c85ec98fcb9acd86d0cdd4c9d87ade;
    decBuf[9430] = 256'h4ce5b8eb38f348fa89024d0a5c11c817481f5826c32c4334583d7143354b4a54;
    decBuf[9431] = 256'h645a28623367c96bf36fbd732f771079c57a4a7bb37c207d847d747cd97ace78;
    decBuf[9432] = 256'h5a751f71226d71672362ef5b1a56cc50984ac344753fa23a0035b22fdf2a7e26;
    decBuf[9433] = 256'h5e218b1c29182d148e10340e100cad0b520ba50b5a0b260cdf0cf80dc30f7311;
    decBuf[9434] = 256'h6c13d01510181b1a071df91e27224b243c26b628f52ad62b2a2d672dbf2c8c2c;
    decBuf[9435] = 256'h472bcc2901285a252b22521ea91948152810550bb305650032fab1f2a6ed65e5;
    decBuf[9436] = 256'hd9dfcad85ed289ccb7c521c14bbbfdb52bb1c9accda82da5d3a2b0a0be9e649e;
    decBuf[9437] = 256'hb69e969ffaa13aa470a725ac46af66b499ba6fc0bdc5f0cbc6d198d8d9e09de8;
    decBuf[9438] = 256'hacefc3f979000309c710dc196622f227022f6d35ee3cf9418f46b94a834ef551;
    decBuf[9439] = 256'h1755cc565057b9582759fc57ed56f655eb538751a34eea4b074867442c400c3b;
    decBuf[9440] = 256'h3936d831942bbf25f521c11b97174912760d14093b069c0261feabfc15fabbf7;
    decBuf[9441] = 256'h72f648f538f48bf440f484f43df556f655f7f6f8effa43fcebfe640148048f08;
    decBuf[9442] = 256'h8b0c341195159219281c731f962188234c25e7265d28b129612bea2cb52eea2f;
    decBuf[9443] = 256'h73317232fd3227331b325530ae2d342b50289825d3239321f31ec41bc6180d16;
    decBuf[9444] = 256'h9413af10300dd60afd0666040c02e9fff7fd33fc97fa22f9cef71df695f430f3;
    decBuf[9445] = 256'h8ef105f0d2ef01f0d3f079f273f44ff67af886faeafc85fefbffc700fb011403;
    decBuf[9446] = 256'hdf048f06f908380b440da80fe711f313cf157f172718c018ef181919f218cf18;
    decBuf[9447] = 256'h7118a71725171f165a14aa12d00f510c0609080688022e0055fcbef974f675f3;
    decBuf[9448] = 256'hf6ef9cedc2e923e6e7e1ebdd4cda10d614d274ce1bccf7c9cdc8bdc76bc78bc6;
    decBuf[9449] = 256'h47c68dc555c588c5b7c535c65bc60ac7a8c7abc82acaf5cba5cd9fcf03d242d4;
    decBuf[9450] = 256'h4ed63ad9f2db6cde50e108e482e666e958eb1cedb7ee2df0f9f02ef246f345f4;
    decBuf[9451] = 256'h2df5a8f6a7f749f9d2fad1fbb9fc8bfdb2fd8ffdaefd92fdacfdc3fd57fd1cfd;
    decBuf[9452] = 256'h0bfd99fc6dfc5ffcf2fb6dfbccfa0afa53f90cf9f6f831f9aef920fa87faaffa;
    decBuf[9453] = 256'h42fa65f948f8eff6aaf5d8f4cbf3d7f278f222f208f21ff260f274f262f2f0f1;
    decBuf[9454] = 256'h13f1b7ef16ee8dec28ebe3e911e9eae882e823e893e7a8e64ce564e43de331e2;
    decBuf[9455] = 256'hc8e12ae19ae080e098e02fe107e297e2e5e22ce395e2bde1f4e0d4df15dff2de;
    decBuf[9456] = 256'h51df1ae0a2e12be3f6e4a6e64ee74de8d8e8aee888e8d9e7bde663e51fe4f8e2;
    decBuf[9457] = 256'h85e2d6e138e1a9e0f2dfecdef8dd9cdc58dbddd978d87ad626d575d3ecd187d0;
    decBuf[9458] = 256'he6cecdcdcecc8acb0bcbe5ca7cca9cca2ccbaecb13cdaacf23d250d670db43e0;
    decBuf[9459] = 256'ha5e4e8eabdf00bf63ffc14026207960d6b13b9184e205d279e2f9a3950404c4b;
    decBuf[9460] = 256'hae52135c2d62b967c96e8971b475fa770b7aab7a607cee7d667ed47e377fdd7e;
    decBuf[9461] = 256'h417d367b4a78cb748f70706b3c65675f195a8452794d3845ac3fa13a3634b62c;
    decBuf[9462] = 256'haa273f21691b9f17cd126b0e920bfc08a20659052f041f03cd02ed01a9016b01;
    decBuf[9463] = 256'ha3013c0224039f04d0067109a00c7910191463173d1bca1c241f6d20d0207620;
    decBuf[9464] = 256'h2320431fef1d3f1c461a6a18b916c014d4111c0fed0b3907d70294fcbef670f1;
    decBuf[9465] = 256'h3deb67e595de2ad8aad09ecb33c5b3bda7b812b43cae72aa00a7dfa306a182a0;
    decBuf[9466] = 256'h09a077a0a1a1b1a24ca457a633a8dbaa09aee3b18bb62dbcffc26bc9ebd0ffd9;
    decBuf[9467] = 256'h8ae286ecebf576fe7208d711f117b51fc526302d0633d8396d3e43449149644e;
    decBuf[9468] = 256'hc552c2565859a35ceb5ddd5f825f305fba5d565b7258f354b750974bc5462341;
    decBuf[9469] = 256'hd53ba1357631282c5627b321e91d1719b514b910100caf078f02bcfd5af95ef5;
    decBuf[9470] = 256'hb6f0d5ee20ed92eb0bec78eca3ed67ef02f1a3f31df601f9b9fb33fe1701d003;
    decBuf[9471] = 256'hfe06fd09b50c2f0f1312cb144517291a1b1c941e2f203b2217244b256426fd26;
    decBuf[9472] = 256'h2b27ad26a025db23af21791e9f1a0017c512a50d330ad105d50135feebfaecf7;
    decBuf[9473] = 256'h34f5baf27bf06fee0beccce92be7b1e472e266e08ade56ddaddc7adc05ddd8dd;
    decBuf[9474] = 256'h31df2fe10be3b3e52ce8b5eb0feee8f17ff4c9f7c8fa47fe9201910449070e09;
    decBuf[9475] = 256'h4d0bc30c170e4c0f641063114b12ca123d13a5138613301379127311ae0f820d;
    decBuf[9476] = 256'he20ab307da033a00effc16f97ff635f35befc5ec7ae97ce6fce2b2dfb3dc34d9;
    decBuf[9477] = 256'hdad6dbd3ead125d02ecf4ece0acecccd75cea8ce33cfb1cfbed0b2d10ed353d4;
    decBuf[9478] = 256'hced599d749d942dba6dd8ae07ce2f5e435e740e91cebcdec55eebaeffff026f2;
    decBuf[9479] = 256'h33f39bf339f490f475f45ef41df493f316f364f2bdf126f19df01ff0ceef67ef;
    decBuf[9480] = 256'h09ef6ceed4edd5ec27ec49ebbaea6bea54ea69eacbea90eb7bec98eda4eedeef;
    decBuf[9481] = 256'hb1f071f11ff2bdf2c0f36ef48bf598f646f763f86ff963fa01fbcbfbe5fb2cfc;
    decBuf[9482] = 256'h42fc55fc67fcb8fcaafc9cfc90fc17fc85fb86fa06f9a1f7a3f5c7f317f28ef0;
    decBuf[9483] = 256'hc3ee13edfaeb95ea50e92ae81de7e3e5bce463e31ee2f7e0ebdf3cdf9ede0ede;
    decBuf[9484] = 256'h8cdd45dd04ddc9dcdbdc0bdd55ddcedd60de10dfe6dfe9e097e1b4e2c1e3b5e4;
    decBuf[9485] = 256'h92e595e643e7e1e771e8bfe866e9d2e934eab1ea80ea37ead9e923e9a0e859e8;
    decBuf[9486] = 256'hc2e738e7bbe6c8e5d3e475e4abe329e3b2e299e18ce00ddf42dd91db98d9bcd7;
    decBuf[9487] = 256'h90d51bd43fd20ad1f1cff2ce67ce95cd21cdb9cc1bcc8bcba0ca44c95cc889c7;
    decBuf[9488] = 256'hcac6a7c6c6c61dc708c824c97eca1fcc88ce24d0c4d23ed522d869dc65e016e6;
    decBuf[9489] = 256'h64eb98f16df73ffeab04800ace0f02162d1a7b1fae25842b5632963a5a426a49;
    decBuf[9490] = 256'hab516f597a5ee56465672f6b416d216fd7706472dc7225748874e3749174b073;
    decBuf[9491] = 256'hd471a96f086dd96900666062345dc2592054d24e004a5d448b3d20374a31782a;
    decBuf[9492] = 256'h0d24e21f941a221742156912db10720f2a0ec60db70c1c0b3b0ae70837078f06;
    decBuf[9493] = 256'hf60524069f076a09960bcc0ea6124516811a591df920432467269127a128f328;
    decBuf[9494] = 256'h3e29ea27b526bc24e0223920bf1ddb1a2318a915c512450ffb0b2108790317ff;
    decBuf[9495] = 256'hd4f8fef2b0ed7de7a7e1d5da3fd66ad01ccbaac748c36fc0d9bd7fbb36ba0cb9;
    decBuf[9496] = 256'hb1b804b979baddbc1dbfbec1ecc4ebc731cc2ed0d6d438d97bdf51e523ec8ef2;
    decBuf[9497] = 256'h0efa1e015f09231133187320ff250b2b7631a1356b393d3e9f427845204a424d;
    decBuf[9498] = 256'h1a50b152fc5544576f587e592c59b657da5533534f4fb04b74475542823d2039;
    decBuf[9499] = 256'h01342e2fcc2ad0262722061f0a1b73181a16f6133e11c40ee00b2709ae066e04;
    decBuf[9500] = 256'hcd0109006efe8dfdd1fd8bfea3ffd4017504ee06770ac20d9b1132147c17c518;
    decBuf[9501] = 256'hb61a7b1c161ef61e4a207f21982231235f23de236a230223242222215c1f311d;
    decBuf[9502] = 256'h251b3918811552122f10760dfd0a190899044e0175fdd5f99af59ef107efbdeb;
    decBuf[9503] = 256'hbee8cde653e45ce3e7e11be161e029e0f6dfc8df46e0b9e0f3e16ee305e67fe8;
    decBuf[9504] = 256'h08ec52ef51f2d0f52af84efa3ffc04fe4300b9011d045d066808cc0a0c0dad0f;
    decBuf[9505] = 256'h71110c138214c61404155c145d137512fa102f0f7e0d150bd508340606030700;
    decBuf[9506] = 256'h88fc3df964f5cdf273f075ed83ebbfe924e8aee6d2e4a6e29be0bfde0fdd86db;
    decBuf[9507] = 256'h21da96d96cd992d940da9cdb3edd37df13e1c3e24ce4b1e599e6c0e7cce84cea;
    decBuf[9508] = 256'hb1ebafed8bef3bf134f310f5c1f649f8aef9f3fa1afcdafc42fda1fd85fd6afd;
    decBuf[9509] = 256'hf4fc5cfcacfb35fb72fabbf915f927f84af7baf638f6f0f5aff54df5d0f41df4;
    decBuf[9510] = 256'h48f345f251f173f0aaeff3ee7dee10ee24ee36eea8ee85efa2f0fbf19cf325f5;
    decBuf[9511] = 256'h8af6cff7a1f815f9c3f961fa2afb15fcf3fcbcfda7fe06ff23ff71ff59ff19ff;
    decBuf[9512] = 256'h53ff1effedfea3fedbfdd8fc9efb23fa58f82cf68bf312f12eee75ebfce8bce6;
    decBuf[9513] = 256'h46e56ae3b1e228e129e088deffdc9adbf8d9e0d8e1d756d72cd705d76ed7cdd7;
    decBuf[9514] = 256'h5cd848d925da61db88dc95dd14df79e0bee139e39ee4e3e50ae716e80ae9e8e9;
    decBuf[9515] = 256'h24eb4bec57ed91ee64efd7ef85f0e4f0c8f0e2f06bf0a8eff1eeecedf8ecdbeb;
    decBuf[9516] = 256'hcfea95e9c2e869e724e6fde4a4e3bce23ee2cbe1a8e149e1b9e0cedf72de74dc;
    decBuf[9517] = 256'h98dae8d8efd69bd566d44dd31ad3ecd216d389d338d415d5ded52dd6a3d6b9d6;
    decBuf[9518] = 256'ha5d6b7d608d735d7fdd73ad9b5da80dcabde21e085e2c5e4d0e6bce93ced86f0;
    decBuf[9519] = 256'h3bf59df9e0ffb505030bd60f7815c61a991fba22b6265f2bc12fe034143be940;
    decBuf[9520] = 256'h3f49cb4edb55465c1c62e6655869396bee6c726ddc6e496fe66e406fee6e0e6e;
    decBuf[9521] = 256'hba6c096ba068bc653c62015ee1580e54ad4f69499443463e12383d326b2b0025;
    decBuf[9522] = 256'h2a1f5818ed11c20d7408020521036c01d5fe5dfef0fdc5fc6bfc18fccefb8afb;
    decBuf[9523] = 256'hc7fb70fcd5fd76ffdf01c40443088e0b670ffe1148154718381afd1b981d0e1f;
    decBuf[9524] = 256'hda1f93205b20c21fda1e0b1ddf1a3e1810151112920e470b6e07ce0393ff97fb;
    decBuf[9525] = 256'he5f597f064ea8ee4bcdd51d77bd12dcc5bc7f9c220c08abd30bbe7b9bdb8adb7;
    decBuf[9526] = 256'h5bb77bb6bfb6fcb6a5b7a4b8a2ba06bd8fc0cac4c6c878cec6d3f9d97ae185e6;
    decBuf[9527] = 256'hf0ec70f480fbeb016c097c10e716671e7223de29092e5733c836a938823b0f3d;
    decBuf[9528] = 256'h693fb2406a432f456f47e448384af24a494a7e4852468742e73eac3ab0360732;
    decBuf[9529] = 256'he62eea2a5328f925fb220921901eab1bf3187916f1129710730e820c720b7c0a;
    decBuf[9530] = 256'h310aed092b0af209250a540ad20a450b7f0ca60de60f2512311495163018a619;
    decBuf[9531] = 256'hfa1ab31beb1b1e1cf01bc61bec1b0f1c6e1cfd1c181d2f1dc31c9d1b221af117;
    decBuf[9532] = 256'h50152112480ea80a6d069403f5ffaafc87facef7a0f4a1f1e9eebaebbce803e6;
    decBuf[9533] = 256'h3fe4ffe189e0bddffbdfc3dff6df24e04ee075e052e0b4df5ddf78df1ee062e1;
    decBuf[9534] = 256'h1ae460e85decfcef47f345f6fef8c2fab9fb99fc65fda3fddbfd74fefffed2ff;
    decBuf[9535] = 256'h4500ae000c0129010f019800aaff8efe34fd93fb0afa3ff88ff606f5d5f234f0;
    decBuf[9536] = 256'hbbed7bebdae861e621e416e24ae191e0c9e0fce087e105e2c5e22ee38de3a9e3;
    decBuf[9537] = 256'h5be3e4e2f6e158e102e185e1b9e2dde47ee7acea86ee1cf167f48af6b5f7c4f8;
    decBuf[9538] = 256'h17f961f91df95bf993f9c6f9f5f9c7fad4fb0efd35fea8fe10ff30ff67feb0fd;
    decBuf[9539] = 256'hdafc11fc26fb48fa0cf991f72cf62ef452f2a2f089ef8aeeffed80edc1ec58ec;
    decBuf[9540] = 256'hf9eba3eb89eba0ebb6ebcaebdcebcbebdaebcdeb09ec98ec70ed73eeadefd4f0;
    decBuf[9541] = 256'h2df2cef3e7f44cf6edf706f96bfab0fb2efca1fcc4fca4fc88fc6efcf7fb5ffb;
    decBuf[9542] = 256'h88fa4bf97cf747f64ef4faf2c5f13cf0d7ee36ed3deb61e9bae640e400e260df;
    decBuf[9543] = 256'he6dca6da9bd837d69cd426d35ad21cd2e4d117d2a2d2cdd240d3a8d346d4d6d4;
    decBuf[9544] = 256'hc1d5ded637d835da11dc3dde48e034e3ede566e8a6ea1cecf8eda8efc1f026f2;
    decBuf[9545] = 256'h6af391f49ef5d8f6aaf76af819f9f9f869f8e7f782f61df5d9f35ef25ff11af0;
    decBuf[9546] = 256'hf3eee7edf2ec57ebcee969e86be68fe4dfe256e157e06fdf48ded5ddb2dd93dd;
    decBuf[9547] = 256'h23ded9de80dfecdfffdfcadf99df8adfcddf53e0d0e0a3e16ce257e335e471e5;
    decBuf[9548] = 256'h44e650e744e8e2e839e987e96fe9b0e9ebe944ea18eb54ec7bedd4ee19f040f1;
    decBuf[9549] = 256'h99f297f4fbf6dff926fe2202cb062c0b290fd11333182f1ccf1f0a240628af2c;
    decBuf[9550] = 256'h51329f37723c5443c049954f6756fd5ad3609d64ae668f68446abf69386aca69;
    decBuf[9551] = 256'h67695768bc664665f2634262d95f995d635a8956e1517f4d3c476641943a2934;
    decBuf[9552] = 256'ha82c9d2732215c1b92175f11340d6a09f805d70222018bfe22fdb4fc8afb2ffb;
    decBuf[9553] = 256'hddfa28fb6cfb25fccefc33fe77ff9e0091026d041407f80a970ed312cf166519;
    decBuf[9554] = 256'hb01cd31efe1f0d2160211521d1209c1f131eae1c531a1418dd14df115f0e060c;
    decBuf[9555] = 256'h2c088d04420168fdc9f98ef591f1e9ec87e867e395def2d8a4d333d0d1cbd5c7;
    decBuf[9556] = 256'h47c6edc380c31cc377c312c588c6ecc8d0cb4fcf9ad274d61cdb3dde3ae2e2e6;
    decBuf[9557] = 256'h44eb64f097f66dfc3f03aa092a113a18a51e2626352da133cb37193d8b40ad43;
    decBuf[9558] = 256'h6245f8476149aa4a9b4cf64ced4d374e7b4ec24d1a4d4f4ba8482e46a5426a3e;
    decBuf[9559] = 256'h6e3ac5356331672dbf285d246120c11c7719531762159d1302128c10c00f070f;
    decBuf[9560] = 256'hee0dbb0dd30c550c2f0c510cb00cb30ded0e111147144517c51a001fd9216f24;
    decBuf[9561] = 256'hc926ed28172adc2b2e2c792cad2bf42a4b2a4c2964283d273126b124e6223f20;
    decBuf[9562] = 256'hc51de11a621726132a0f820adf0491ffbffa1cf5ceeffcea9ae69ee207e09ede;
    decBuf[9563] = 256'h7bdc50db41da4ad9ffd833d87ad742d70fd7e0d60bd7cad704d9d4daffdca0df;
    decBuf[9564] = 256'hcfe2cde54de988ed84f11bf456f82ffbc5fd1f0043026d03c8031a0465049903;
    decBuf[9565] = 256'he00237023801500029ff1dfe29fd0cfcb3fa11f918f73cf510f305f1a1ee61ec;
    decBuf[9566] = 256'hc1e992e694e3a2e129dfe9dc73dba7da69da31dafed989da5cdbb5dc57de50e0;
    decBuf[9567] = 256'h2ce2dce365e5cae60fe836e98fea30ecb9ed1eef1cf1f8f2a0f519f859fa64fc;
    decBuf[9568] = 256'hc8fe08011303df039804600461037902a7019a00ecff51fec8fc97fa8bf837f7;
    decBuf[9569] = 256'h03f6eaf451f423f4a4f3e4f236f219f173efeaedb9ebaee94ae7afe5a4e350e2;
    decBuf[9570] = 256'h1be1e3e016e1fee1cde3f9e504e8e0e990eba9ec0eee53ef79f0d3f117f3eaf3;
    decBuf[9571] = 256'haaf458f5f6f54df69bf6e2f6f8f65af790f7e1f748f856f819f8b6f7edf624f6;
    decBuf[9572] = 256'h39f5ddf33cf243f0dfedfaea09e98fe650e444e2e0df45de3adc5eda32d8bcd6;
    decBuf[9573] = 256'h68d534d48bd358d387d305d4c5d4b9d515d759d829da55dc60de3ce0ece194e2;
    decBuf[9574] = 256'h93e37be4a2e548e7b2e996ec4eef7df27bf5fbf846fc44ff3601af03a604f104;
    decBuf[9575] = 256'had046f045603f101ad0086ff79fe85fda8fca5fb25fa5af82ef6b9f4ddf2a8f1;
    decBuf[9576] = 256'h8ff090ef4cee7cecccead3e86fe62fe424e2c0df25de44dd00dd3edd57de22e0;
    decBuf[9577] = 256'hd2e1cbe31fe554e66de706e891e8bbe894e8b7e816e96ce958ea35eb38ece6ec;
    decBuf[9578] = 256'h84ed14ee97eeaeeeefee2aef18ef28ef55ef12efedeeb6ee34eedbedaaed61ed;
    decBuf[9579] = 256'h53ed78ed83edf1edceeea8f094f3dbf7d7fb8801d606a90b0b102b159c18fe1c;
    decBuf[9580] = 256'hfa20a325052a012ea9320b372b3c5e423448064f9c537159bf5e316252650867;
    decBuf[9581] = 256'h95680e69a0683d687866dd64d262e65f2d5db45a2b57e05307505e4bbc456e40;
    decBuf[9582] = 256'h3b3a6534932d28275221801aea156a0e5f09f302c9fe7bf909f6e7f20ff081ee;
    decBuf[9583] = 256'h09eec0ec24ed7eedd1edb1eef5eeaeefc7f0c6f10af3daf405f73cfa3afdba00;
    decBuf[9584] = 256'hf504f108910ceb0ee911db13ea1498144d14091450133712d210d40e700c8c09;
    decBuf[9585] = 256'h0c06d101f8fe50faeef5f2f152ee17ea1be672e110dd14d96cd40ad0eaca18c6;
    decBuf[9586] = 256'hf6c2fabe6dbd03bcbbba1ebbe3bc7ebe89c075c32ec65cc95bccdacf16d436d9;
    decBuf[9587] = 256'ha7dc4ae21ce9b1ed32f542fcad022d0a3d11a8177e1d5024e628bb2e09347b37;
    decBuf[9588] = 256'hdd3bb63e43409d42e54310456a45bd45dc449844df433743d2418d406a3e5e3c;
    decBuf[9589] = 256'h7239f335b731bb2d1329f125f521561e0b1b0d18541590135011da0f0e0f550e;
    decBuf[9590] = 256'hac0d790d4b0d750d820ebc0f371102132e15a3167f18301a481b131dc31e4c20;
    decBuf[9591] = 256'h7d228924ed262c29cd2bdd2c782ec32e072f4d2ea52dda2b2a2ac0278125e022;
    decBuf[9592] = 256'h6620821dca1a9b17c2132210d70cd90959060f03100091fc46f948f68ff361f0;
    decBuf[9593] = 256'h3dee85eb0be9cbe656e58ae44ce484e41de505e62ce785e827eaafeb7aeda6ef;
    decBuf[9594] = 256'hb1f18df3b9f52ff70bf940fac9fb2efd72feedffb801ed020604050533055d05;
    decBuf[9595] = 256'h370514053704fa027f014eff43fd67fb3bf99af621f4e1f140ef12eceee936e7;
    decBuf[9596] = 256'h71e5d6e3cbe177e0c7de3eddd9db37daafd8b0d724d7fad66dd762d87ed9d8da;
    decBuf[9597] = 256'h1cdcecdd9cdf95e1f9e339e644e8a8ea43ec4eeea2ef53f1dcf241f485f5acf6;
    decBuf[9598] = 256'hb9f7f3f819fad9fa88fbe7fbcafb7bfbd5fabcf9aff830f765f539f32ef1caee;
    decBuf[9599] = 256'h8aec7fea2be9f6e7dde644e6b9e5e7e4dae32ce30fe24fe1a1e042e0ecdf06e0;
    decBuf[9600] = 256'heedf2fe0b8e07de19ce2f6e33ae50ae7bae843ea74ec7fee5bf00bf224f3bdf3;
    decBuf[9601] = 256'h48f4c6f4edf410f56ff5fef5e9f6c7f790f847f9bef9a8f946f9edf83af894f7;
    decBuf[9602] = 256'hfcf6fdf5c3f448f37df151ef46ed6aebbae9a1e8a2e774e74ae723e700e7e1e6;
    decBuf[9603] = 256'h8be608e632e569e47ee3e0e250e236e2ade244e31ce4e5e4d0e5aee6b0e7a4e8;
    decBuf[9604] = 256'hc1e91aeb5fec2eee5af0d0f1acf35cf575f674f7fff729f84ff872f813f8f7f7;
    decBuf[9605] = 256'h11f8f9f70ff84af814f8e3f7d4f727f751f64ef514f445f295f02beeebebe0e9;
    decBuf[9606] = 256'h04e8d8e563e497e362e22ae291e162e138e1c5e017e079dfafde61de49de8ade;
    decBuf[9607] = 256'h14dfd8dfc3e0e0e139e37ee4a5e5b1e6ebe7bee8cbe904eb80ece5ede3ef37f1;
    decBuf[9608] = 256'h6bf214f347f3bcf2e9f190f0eeee65ed00ecbceae9e976e90de96fe819e82ee7;
    decBuf[9609] = 256'h11e6b8e4bae2dee02edfa5dd0cdd3add64ddbede02e029e1cfe2c8e4a4e64ce9;
    decBuf[9610] = 256'h7aec2ff190f5d4fb5403640acf104f185f1fa0272c2d3c34d138a73ef543284a;
    decBuf[9611] = 256'hfe4fd0563b5dbc64cb6b377261762b7a3d7cdd7c287b9a7940774274fb6fff6b;
    decBuf[9612] = 256'h5667f562f85e595b2d56f94f244a5243113b4d33392a1f245b1c47132d0d6905;
    decBuf[9613] = 256'h5e00f2f91df4cfee5deb3ce863e5dee466e4aee5a0e719eaa2ededf0a1f5c3f8;
    decBuf[9614] = 256'hbffc55ffa0029e051e09590d5611fe15a01bee2022274d2b9b300c342e37e338;
    decBuf[9615] = 256'h703af839b038be364534bc30802c8428d322851db218cf113a0d64071602e3fb;
    decBuf[9616] = 256'hb8f76af236ec61e68fdf23d94ed37ccc11c6e6c11cbe0bbc2ababcba40bb9abd;
    decBuf[9617] = 256'h98c051c334c7d4ca0fcf0cd3bdd80bde3ee414eae6f051f7d2fee1054d0ccd13;
    decBuf[9618] = 256'hdd1a48211e27f02d5b34313a7f3f514472474b4ad94b424df94bcf4a55487145;
    decBuf[9619] = 256'hb9423f40ff3df43b183a713742344431c42d89298d25e420421b7817a512440e;
    decBuf[9620] = 256'h6b0bd4085c081307b0060a075d073d0809093e0aa70ce70e1d121c159b18e61b;
    decBuf[9621] = 256'he41e9d211624fa26ec28652ba52db02f1432b03325357936ae37e63719388e37;
    decBuf[9622] = 256'hbf359333f2300f2d6f2925264b22a31d411945159c103a0c1b074802a6fc58f7;
    decBuf[9623] = 256'he6f384ef88ebf1e8a7e583e392e1cddfd7de61dd95dcdcdba3db0adb39dbb7db;
    decBuf[9624] = 256'hc4dc89de30e15fe45de7a4eba0ef37f281f580f838fbb2fd4dff5801ac02e103;
    decBuf[9625] = 256'hfa04f905e106b307c0086e098e09ab09f408bf07f005c403b90155ff70fcb8f9;
    decBuf[9626] = 256'h89f666f4e6f08cee69ecb0e9ece751e6dbe487e3cee225e2f2e1c4e1eee161e2;
    decBuf[9627] = 256'h10e3aee377e496e5a3e623e8eee919ec25ee11f102f37cf5bbf75cfa21fc60fe;
    decBuf[9628] = 256'h6c004802f8038105e60671079b078e0654058503d5014c00e7fefffd81fd0efd;
    decBuf[9629] = 256'h5ffc82fb46fa76f84af6aaf37bf07dedc4ea00e9c0e6e0e59ce5d9e512e611e7;
    decBuf[9630] = 256'h55e8d4e893e9b6e9d6e99feabfeb65ed5eefc2f102f477f553f77ff9f5fa59fd;
    decBuf[9631] = 256'hf4feff00db02100499059806dd070309100a040b630bd30ae8094d085406f003;
    decBuf[9632] = 256'h5502df008bff56fecdfc68fb24fa00f8f5f591f351f1b0ee37ec53e961e79de5;
    decBuf[9633] = 256'ha6e4c6e382e344e39be268e281e1aee0eedf85df66dff6df78e04ee151e2ffe2;
    decBuf[9634] = 256'hdce3dfe48ee52ce6bbe672e748e811e931ea3deb31ecd0ec26ed0ced65ec4ceb;
    decBuf[9635] = 256'h8cea98e9fae8a4e88ae8a2e8e2e8cfe8bde8ade845e8b2e702e7cde5a6e44de3;
    decBuf[9636] = 256'h65e292e1b9e167e284e3dde4c5e543e66ae601e663e5d3e485e49ce48ae5a7e6;
    decBuf[9637] = 256'h00e8a2e92beb90ecd4edfeed25eebceddfec4fec01ece9eb55ec06edaced43ee;
    decBuf[9638] = 256'hcdee97ee05ee2dedb7ebb8ead0e9fee88ae8ade88ee871e8eee748e72fe6d6e4;
    decBuf[9639] = 256'h34e3abe146e002dfdbdd81dcf6db78db05dbe2da41db97db1adcefdcb9dda4de;
    decBuf[9640] = 256'h00e0e8e063e22ee4dee5d7e73bea1fedd8ef06f3e0f688fb2b017906ac0c8212;
    decBuf[9641] = 256'h5419bf1f3f274f2ee532ba38083edb423d47394bd84e14533458065d68618866;
    decBuf[9642] = 256'hfa691b6dd06e556feb6dc86b4868fe6424617c5c1a58fa52284ec649a644d43f;
    decBuf[9643] = 256'h313a5f33f42c7425641ef9172312510bbb06e60098fb26f8c4f3ebf055eeecec;
    decBuf[9644] = 256'ha3eb40eb9aeb91ec32efabf134f56ff98ffe010263065f0afe0d49112315b917;
    decBuf[9645] = 256'h041b021ebb20e9230d26c5288a2a252c9b2ddf2d252d9d2b062922257a20181c;
    decBuf[9646] = 256'hd515ff0fb10a7e04a8fed6f795ef09eaf9e264de8ed840d30dcde2c894c322c0;
    decBuf[9647] = 256'h01bd28ba9ab831b7e9b54cb6f2b5e9b65eb8c2ba4bbe86c2cac89fce71d5dddb;
    decBuf[9648] = 256'hb2e184e8efeec5f497fb0202d807aa0e40131519631e36239827942b2a2e8430;
    decBuf[9649] = 256'ha8329934a935a036ea36a636ed35f4339031072ecc29d0252721c51cc9182a15;
    decBuf[9650] = 256'hd012ac10bb0ef60c5b0be5099108e1065805590471034703ba03f40418072309;
    decBuf[9651] = 256'h870b6b0e5d108b13af152e19791c771ff72241264029f82b272f4a3175328433;
    decBuf[9652] = 256'hd733f632a231f22ff92d952bb128f825ca22cb1f851b8917e0127e0e820ada05;
    decBuf[9653] = 256'h780158fc85f724f304ee31e9d0e4f7e157defddbdad9e8d7d9d687d63cd608d7;
    decBuf[9654] = 256'h3dd855d920db4cdd57df43e2fce475e7feea49ee47f1c7f402f9dbfb8300a503;
    decBuf[9655] = 256'ha107370a820da50fd010df113212e7111b116210490fe40d430cba0a55095707;
    decBuf[9656] = 256'hf304b3027dff7efcfff8b4f5dbf144eff9ebfbe809e790e4f5e27fe1b3e07edf;
    decBuf[9657] = 256'h46dfadde7fdea9de1cdf10e06ce10de377e5b6e757ead1ecb5efa6f120f460f6;
    decBuf[9658] = 256'h6bf847fa73fce8fdc4fff900820281030c048b04b1044804aa036e029f00eefe;
    decBuf[9659] = 256'hf5fc91fa51f846f66af43ef29eef24ed89ebe8e824e788e57de329e270e1c8e0;
    decBuf[9660] = 256'h2fe05de087e047e1f5e151e396e4bde563e77be8e0e9dfebbbed6bef44f2fdf4;
    decBuf[9661] = 256'h2bf82afbe2fd11013403260535062c070c08500813084b087e084f0825086507;
    decBuf[9662] = 256'hb7069a05f4036b023a002ffe53fca3faaaf856f72af5b4f3d8f128f02fee53ec;
    decBuf[9663] = 256'hace9e7e7a7e532e456e29ce1f4e05be02de003e029e092e030e1bfe176e21de3;
    decBuf[9664] = 256'h89e3c4e3b2e381e372e380e3ede38fe47de55ae65de70be86ae887e86de855e8;
    decBuf[9665] = 256'h14e8b2e759e7e7e662e6e5e594e50fe5d9e4a9e49ae4a7e4fce433e5a1e508e6;
    decBuf[9666] = 256'h66e6ebe68ce7f8e7d0e89ae9b9eac6eb8bed3bef34f110f33cf547f7abf947fb;
    decBuf[9667] = 256'h52fd2effde00670266034e04cc043f0562050305e7043004b9034d03c3022302;
    decBuf[9668] = 256'hb601df00dcff5cfe91fc65fa5af8f6f512f359f0e0edfcea0ae991e6f5e480e3;
    decBuf[9669] = 256'h2ce272e1abe178e103e22de253e276e2d5e2f2e240e387e3f3e32ee488e43ae5;
    decBuf[9670] = 256'h10e613e74de8c8e92deb72ec41ee76effff064f2a8f323f588f6cdf7a0f8acf9;
    decBuf[9671] = 256'h15fab3fab6fb64fc41fd7efea5fffe00fc02d8047f07ae0a870e3013d218201e;
    decBuf[9672] = 256'hf3225427742ce62f48342137c03a1a3d18409843e346e149284e0051a955ca58;
    decBuf[9673] = 256'ha35b395ea25f1060ac5fe85da85b72589854f04f4e4a0045cc3ea13a5335202f;
    decBuf[9674] = 256'hf52aa725d520731c53178012de0c1409e102b6feecfa7af718f363f1d6ef7ced;
    decBuf[9675] = 256'h0eed72edcced0cf0adf2dbf5b5f95dfebf02df07b10c13113316a519061edf20;
    decBuf[9676] = 256'h7623df2402272d283c29332a132bdf2b992cd12c382cf32a7b289824f820db1a;
    decBuf[9677] = 256'h0615b80f84090402f9fc8df6b8f06aeb97e6f5e0a7db35d8d3d3fbd064ce0acc;
    decBuf[9678] = 256'hc2ca5ecab9caafcb25cd89cf6dd2edd538d911ddbae15ce7aaecddf2b3f885ff;
    decBuf[9679] = 256'hf005700d80141619ec1ebe25532a7e2e4832ba359b37743a013c793ce73c833c;
    decBuf[9680] = 256'h293c8e3a1839b436d0335030062d072a88263d23631fc41b89178c13ed0fa20c;
    decBuf[9681] = 256'ha409eb0627058b03ab02df011d0236039b04f506da09920cc10f9a133a17841a;
    decBuf[9682] = 256'h831d02214d244b27042a322d562f0e3288346c37253a9e3c393e1a3fe63f2c3f;
    decBuf[9683] = 256'h143ee33b42395f35bf31932cc0271e22d01cfd179c137c0ea90948054b01a3fc;
    decBuf[9684] = 256'h82f985f5eff2a4ef81edc8ea04e9c4e6b9e465e3abe273e20ce351e420e6c8e8;
    decBuf[9685] = 256'hf6ebd0ef6ff3aaf7a7fb46ff91028f0548080c0a4c0cc20d9e0f4e11d7123c14;
    decBuf[9686] = 256'hc71445156c154915ea145a143b132e12af10e40e330dab0be0092f0836065a04;
    decBuf[9687] = 256'haa02b1004dfe0dfc02faaef879f7d1f69ef629f750f8a9f94afb44fd20ff4b01;
    decBuf[9688] = 256'hc1029d04d205ea0683076b083e094b0a3f0b5b0c680d5c0efa0e500f9f0f580f;
    decBuf[9689] = 256'heb0e140e110d910bc6099a078f05a302ebffbcfc99fae0f7b2f48ef29df023ee;
    decBuf[9690] = 256'h88ec12ebbee989e871e772e6e7e5bde5e3e506e6a4e66de78de899e919eb7eec;
    decBuf[9691] = 256'h7cee58f084f28ff47bf76cf9e6fb26fe9bff7701ac0255038803b6038c031903;
    decBuf[9692] = 256'h6a02cc01c9001b003eff01fe86fcbbfa90f8eff575f3edef93edb9e923e7c9e4;
    decBuf[9693] = 256'hcae112df4dddb2db3cdae8d8b4d79bd602d677d5a4d47ed45bd4bad44ad500d6;
    decBuf[9694] = 256'hd6d6d9d742d8e0d86fd9bed964da52db2fdcbfdc42dd89dd9fddb2dda0dd70dd;
    decBuf[9695] = 256'h26ddc8dc5bdcb9dbf6da0bda2ed92bd837d759d657d5a8d449d4bad36bd383d3;
    decBuf[9696] = 256'h99d322d4e7d49ed573d676d76ad8c6d967db61ddc5df04e210e4fce6b4e92eec;
    decBuf[9697] = 256'h6dee0ef1d3f212f51ef7faf8aafa33fcfefdaeff370136021e039c0376035303;
    decBuf[9698] = 256'hb50278015200f8fefafc1efb6ef904f7c5f44ff3ebf0abeea0ec3ceafce7f1e5;
    decBuf[9699] = 256'h8de34de1d7dffbddc7dc3edbd9d937d88fd790d662d68cd6ffd668d784d891d9;
    decBuf[9700] = 256'h10db41dd4ddfb1e1f0e3fce550e784e89de936ea1eeb9ceb0fec78ec98ecb4ec;
    decBuf[9701] = 256'h66ec1fecdeeb55ebfbea89eae7e950e99fe89ae7ece64de684e5cde427e464e3;
    decBuf[9702] = 256'haee296e280e20ae316e455e695e861ec09f16bf5aefb2f033e0aaa107f16511d;
    decBuf[9703] = 256'hbd239229e02eb33355391f3df2415346504af84e5a533356d2592c5c755dd85d;
    decBuf[9704] = 256'h145cd45908566051fe4cbb46e540133ad2310e2afe22931c1315030e98071700;
    decBuf[9705] = 256'h08f99cf2c7ec79e7a6e285dfacdc16daadd864d701d75bd7f6d802dbeedd6de1;
    decBuf[9706] = 256'h99e66ceb0ef1e0f74bfecc05db0c4713c71ad21f682493285d2c6e2e4f300432;
    decBuf[9707] = 256'h893201336e330b33fb31bc2f1b2dec2913266120131b7f13700c040684fe74f7;
    decBuf[9708] = 256'h33ef6fe760e0f4d9cad57cd0a9cb88c8afc518c3afc142c1a5c100c240c4e0c6;
    decBuf[9709] = 256'hc4ca63ce8fd3c3d998dfe6e47bec8af3f6f9cbff9d06080d89149419ff1fd525;
    decBuf[9710] = 256'h232bf62f1733cc345a36e13574354934d031902f5a2c8028e124a520a91c0a19;
    decBuf[9711] = 256'hce14d210290cc807a802d5fd74f977f5d8f18dee6aec3febe5ea37eb17ec7bee;
    decBuf[9712] = 256'h5ff1dff41af93afe0d03af08fd0dd0127218441fda23af29fd2ed033f136ed3a;
    decBuf[9713] = 256'h843dde3f01422c43d142da416540893e663b673821342530732a2525f21e7117;
    decBuf[9714] = 256'h6210f609760266fb26f39aed8ae6f4e11edc54d882d361d088cdf1ca88c91bc9;
    decBuf[9715] = 256'hb7c8c7c962cb98ce97d1ddd5d9d982de24e4eee7c1ec63f22df600fb61ff8104;
    decBuf[9716] = 256'hf307550c2e0fcd1218163b182d1a3c1b8e1b441bf019bb18c216e614ba121910;
    decBuf[9717] = 256'ha00dbc0a0308d504fb0065fe0bfc0cf91bf756f516f336f26af12cf1f4f08df1;
    decBuf[9718] = 256'h18f2ebf2f8f377f542f76ef979fb65fe1e014c044b07030a7d0cbd0ec8101c12;
    decBuf[9719] = 256'h5113f9132c14fe132b13d2113010370e5b0cb4093a07fb045a02e0fffcfc44fa;
    decBuf[9720] = 256'hcaf78af5eaf270f030ee25ec49ea1de8a8e654e59ae4f2e325e40de534e627e8;
    decBuf[9721] = 256'h03ea2eeccfee49f188f329f6a3f887fb78fdf2ff3202d2049706d7084c0a180b;
    decBuf[9722] = 256'hd20b990b660b7f0a030938070d056c02f2ffb3fda7fb43f95ff6a7f32df1edee;
    decBuf[9723] = 256'he2ec7eea3ee833e657e422e39ae19be0b3df34df0edf31dfcfdf5fe07ee1d7e2;
    decBuf[9724] = 256'h1ce497e562e712e90ceb60ec10ee99ef64f198f2b1f316f55bf682f78ef83df9;
    decBuf[9725] = 256'h9bf97ff9fcf8f7f7bdf642f577f3c7f1cdeff1ed41ecb8ea53e90fe8e8e628e6;
    decBuf[9726] = 256'h7ae5dbe4bfe4a5e4bce428e5b2e59ae6b7e710e9b2ea3aec9fed9eef7af12af3;
    decBuf[9727] = 256'h23f587f7c7f9d2fbbefeaf00de030106f3076c0a080ce80c2c0d6a0d320d990c;
    decBuf[9728] = 256'h0d0ce70ada092c090f084f071506ee049503f4016b00a0feeffc67fb02fabdf8;
    decBuf[9729] = 256'h96f7d6f628f68af5faf4acf464f44ff462f474f4c5f42df5a5f558f62ef730f8;
    decBuf[9730] = 256'h6af991fa51fbbafb18fcc2fb74fbfdfa66fa04faaaf99af98bf999f9bdf9c8f9;
    decBuf[9731] = 256'h82f9f9f821f8abf646f548f36cf141efcbedefebbaeaa1e9a2e8bbe7e8e6dbe5;
    decBuf[9732] = 256'h2de58fe4ffe3e5e3fde312e4c3e4c8e502e7d1e8fdea08ed6cef51f242f4bcf6;
    decBuf[9733] = 256'ha0f991fb0bfe4b005602ba049e07e50be10f9215e01a75228429f02fc535133b;
    decBuf[9734] = 256'h474171453b49ad4c8e4e4350da5243548b55b656c5576159ab59ef593659ad57;
    decBuf[9735] = 256'h1655e8510e4e6f4a434570400e3cef36bb30902c422770220e1eee181c14790e;
    decBuf[9736] = 256'h2b09b90558017ffee8fb8ff946f8e3f7f2f8e9f95ffb3bfde2ff10030f068e09;
    decBuf[9737] = 256'hca0dc6116e16d01af01fc3242429212db72f1132343426368036d3368836bc35;
    decBuf[9738] = 256'h03357a33af31832fe22c692a3c263f22971df517a712730c9e0650011cfb47f5;
    decBuf[9739] = 256'h7df1aaec89e98ce5f6e28de144e0e1df86dfd9df4ee1a2e253e4bce6a0e920ed;
    decBuf[9740] = 256'h6af044f4ecf84efd6e024007e30cad107f15e119dd1d7420ce22cc25f726bb28;
    decBuf[9741] = 256'h0d29ee29aa29f02848287d265124b121821e841b0418c913f010470c26094d06;
    decBuf[9742] = 256'hae02540056fd64fba0f904f88ff63bf581f4b9f452f597f666f80efb3cfe1602;
    decBuf[9743] = 256'hb505f109100fe3134518641d37229926952a352e70324935d6363039793a153a;
    decBuf[9744] = 256'hbb39c4384e37fa354a34e031a12f002d862afe26b323ff1e9d1aa116ef10a10b;
    decBuf[9745] = 256'hce062c01defb0cf769f19fed2dea0ce757e5c9e360e2f3e156e266e301e50ce7;
    decBuf[9746] = 256'he8e814ebb5ed2ef013f3cbf5faf81dfbd6fd4f008f023005a907e9098a0c4e0e;
    decBuf[9747] = 256'h8e10041258131114b914ec146114e313d61256118b0f600d540b7809c8073f06;
    decBuf[9748] = 256'hda0496036f02af0101016200d3ffb9ffd0ffe6ff4800a100f3007701f5014602;
    decBuf[9749] = 256'hcb020003310340034d03290334032a032103390332031d03f1029d02e7019400;
    decBuf[9750] = 256'hf2fef9fc95fa55f8b5f586f288efcfec56ea16e875e5fce260e1ebdf1fdfeadd;
    decBuf[9751] = 256'h41dda8dc7adca4dc17dd80dd1ede21df15e0f2e0f5e12fe356e4afe5f4e66fe8;
    decBuf[9752] = 256'h3aea6feb87ececedd4eea7ef1af0c8f0e8f03ef158f111f1d0f020f04aef81ee;
    decBuf[9753] = 256'hf9ec70eba5e979e76ee592e366e15bdf07ded2dc49db4ada62d990d869d8bbd7;
    decBuf[9754] = 256'h9bd77fd764d77cd714d876d83ad925da03db06dc85dd84dec9df44e143e288e3;
    decBuf[9755] = 256'h5ae41ae583e521e63ee658e66fe62fe6f4e59ae5e8e412e449e329e2d0e08bdf;
    decBuf[9756] = 256'h64debedc35dbd0d92fd816d7b1d56dd49ad341d259d1dad01bd0b2cfd2cfeecf;
    decBuf[9757] = 256'ha5d0dad155d3bad415d7b0d851dbcadd66df06e2cbe30be616e8f2e9a2eb9bed;
    decBuf[9758] = 256'h77efacf035f29af3dff405f6c5f6e8f608f7b2f62ff689f5c6f4a7f39af2a6f1;
    decBuf[9759] = 256'h89f07def43ee1ced0fec1bebffe93fe990e8b3e723e7a1e6cbe53be5ede4a5e4;
    decBuf[9760] = 256'h90e4cbe400e531e5b6e533e6e6e6ebe7dfe8fce908ebb7eb94ec24ed72ed8aed;
    decBuf[9761] = 256'ha0ed3dede4ec31ec2cebf2e977e812e714e5c0e394e11ee0cade1add02dc03db;
    decBuf[9762] = 256'h1bda9cd929d9c1d862d8d2d784d70dd7ccd66ad658d689d6f0d69ed7a3d8ddd9;
    decBuf[9763] = 256'h04dbaadc33de98df39e1c2e227e46ce5e7e6e6e771e844e950eaffeadcebdfec;
    decBuf[9764] = 256'h19eeebee45f02cf153f2f9f312f5ddf68df816fae1fb0dfeae002703b006fb09;
    decBuf[9765] = 256'hd40d7d12de16fe1bd1207326c12b94303636003ad23ef441cc446347bd49054b;
    decBuf[9766] = 256'h304c3f4d924d474df34bbe4ac54861467d43fd3fb33cd93831348e2e40296e24;
    decBuf[9767] = 256'hcb1ef9178e11b90b6b069801f6fb2cf859f338f083eef5ec8cebf9eb5dec21ee;
    decBuf[9768] = 256'h61f097f396f6dcfad9fe8103e307df0b8810e914091a7b1ddd21b6245528af2a;
    decBuf[9769] = 256'had2dd82e9c30ef3039316d30392fcf2c902a59278023e01fb41ae21580113d0b;
    decBuf[9770] = 256'h1207c401f1fc4ff785f3b2ee50ea78e7e1e497e173df49de84dc32dc7ddc49dd;
    decBuf[9771] = 256'h7ddee7e0cbe34ae786eb82ef2bf48cf8acfd7f02e006dd0a7c0eb81290153019;
    decBuf[9772] = 256'h7a1c9e1e562166225d23a7236323aa222121bc1f611d221b811807162313a40f;
    decBuf[9773] = 256'h4a0d4b0acc0672047301bbfe8cfb69f977f7b3f5bcf471f4b5f46ff587f6ecf7;
    decBuf[9774] = 256'h47fa2bfde4ffc7036707b20a660fc813c417641b902002246328602cff2f4a33;
    decBuf[9775] = 256'h48360139c53abc3b9c3c583c233b9b39d0372835af32cb2f122d992ab427fc24;
    decBuf[9776] = 256'hcd21cf1e4f1b0518061587114b0d730ad30688036501acfe9dfda6fc5bfc9ffc;
    decBuf[9777] = 256'h59fde2fead00d802e40448072c0a1d0c970e7b116d13e6152618311a0d1c421d;
    decBuf[9778] = 256'hcb1e641fef1f1920a61f3d1f601e5d1d691c8c1b891a9519b7187b175416ae14;
    decBuf[9779] = 256'h25135a11aa0f910e920daa0c2c0c060c290c480c9e0ced0c340d4a0d5d0d930d;
    decBuf[9780] = 256'hc40d2b0ed90ede0f18113f124b13fa139814b51432145c1320125110a00e370c;
    decBuf[9781] = 256'hf709ec071006e40344017fff9bfce2f969f785f4ccf153ef6eec7deab8e81de7;
    decBuf[9782] = 256'h3de6f9e537e6dfe678e7bde838ea9deb3eed37ef13f1c3f24cf417f6c8f750f9;
    decBuf[9783] = 256'hb5fa57fc50fe2c00dc016503ca04b2053006a306c606670611065a058504bb03;
    decBuf[9784] = 256'hd002b401a700b3ff96fe3dfdf8fb7dfa18f977f7eef589f4a1f323f3fcf2d9f2;
    decBuf[9785] = 256'h77f3cef385f45af524f60ff7adf73df8bff836f9a2f904fa81fad3fafffa27fb;
    decBuf[9786] = 256'h03fbb6fa34fa93f9a5f8c7f78bf664f50bf423f3a8f143f0feee2fed7feb86e9;
    decBuf[9787] = 256'h22e786e5e6e221e186df10debcdc7edcb6dc4fdd94de0fe0dae18ae384e560e7;
    decBuf[9788] = 256'h10e999ea98eb39edc2ee8df034f3aef592f811fc6bfe6a0122049c063708ad09;
    decBuf[9789] = 256'h790a320b6a0b370b090b360a76093c0816076f0576039a01f3fe2ffdeffa4ef8;
    decBuf[9790] = 256'h8af6eef479f325f2f0f0d7efd8ee4dee7aed07ede4ecc5eca8ecf6ec6ded30ee;
    decBuf[9791] = 256'h4fefa9f04af243f41ff64bf8c1f915fbc5fcddfd76fe5eff31005700c000a000;
    decBuf[9792] = 256'h11005aff84fe48fdcdfb68fac6f85df61df412f226ef34ed70eb30e9bae766e6;
    decBuf[9793] = 256'hade594e4fbe370e39ae374e351e3b0e3cde34fe425e528e6a8e773e923eb8ced;
    decBuf[9794] = 256'h27ef33f187f2bbf364f4fdf4cef4a4f47ef4d0f371f3e1f25ef2e8f17bf1f2f0;
    decBuf[9795] = 256'h99f027f067efb0ee0aee1ced7eec61ec47ecbeec02eea4ef9df189f441f770fa;
    decBuf[9796] = 256'h49fef2025407970d6c133e1aaa207f26d52e6134713bdc410746554bc74ea850;
    decBuf[9797] = 256'h5d52eb5372530553da51cb50e64d2e4b95463442f03b1b36492fde285d214d1a;
    decBuf[9798] = 256'he2130d0e3b07cf00a4fc56f784f222ee26ea8fe745e421e2f7e0e7dfdee054e2;
    decBuf[9799] = 256'h40e5bfe8ebedbef2a1f90c008c079c0e0715dd1a2b20fe24a02a6a2edc31bc33;
    decBuf[9800] = 256'h7235ff3687363e3514349a31b62e372bfb26ff22561eb4186613940e320a1205;
    decBuf[9801] = 256'h3f00defbe1f739f397edcde95be63ae361e0d3de6addfddc27deecdf74e3bfe6;
    decBuf[9802] = 256'h74ebd5eff5f428fb53ffa1047409160fe012521673194c1cda1d431f8b20ef20;
    decBuf[9803] = 256'h94204220f71f2b1f7b1d821b1e1995154a12710ed10a96069a02f1fdd0fad4f6;
    decBuf[9804] = 256'h34f3eaefc6ed0eebfee963e818e8d4e712e89be966eb0dee3cf115f5b5f8f0fc;
    decBuf[9805] = 256'hec008c04c708c30c6310ad138717261b711e7021ef2449276c295e2b6d2cc02c;
    decBuf[9806] = 256'h0a2d3e2c852b8c29b027842579231521d51e351cbb19d716e514b711930fa20d;
    decBuf[9807] = 256'hdd0b420acc08f006c504b9026501310088ff55ff27ffa5ffccffa9ff89ff33ff;
    decBuf[9808] = 256'hb0fe0afe73fdc2fc1cfc84fbfbfa7efa4dfa3efa16faf2f94df948f80ef73ef5;
    decBuf[9809] = 256'h8ef395f1b9ef09ee80ec81eb99eac6e953e976e914ea17eb97ecfced9def26f1;
    decBuf[9810] = 256'hf1f2a1f40af74af955fbb9fdf9ff9a025e04fa050508e109160b9f0c9e0d290e;
    decBuf[9811] = 256'hff0dd80d2a0d8c0c890b950afa08710740059f0271ff72fcf3f8b7f4def136ed;
    decBuf[9812] = 256'h15ea3ce7a5e43ce3cfe26be2c6e218e338e2f4e13be102e1cfe05be12de220e4;
    decBuf[9813] = 256'hfce5a3e81deb5ded68efccf167f3ddf431f666f77ef8e3f928fba3fc08fef0fe;
    decBuf[9814] = 256'hc2ff9cffa8fe4cfd4efb62f8a9f57bf27cefc4ec4aea0be895e641e50ce4d4e3;
    decBuf[9815] = 256'h07e435e460e486e41de47fe329e372e22be2c2e2e9e3b8e55fe8d9ea18edb9ef;
    decBuf[9816] = 256'h7ef119f3f9f3c5f47ef5b7f584f555f52bf56bf403f464f362f2e2f017efebec;
    decBuf[9817] = 256'hb5e9dce53ce201de04da6ed723d400d20ed0ffce64cd83cc3fcc02cc3acc6dcc;
    decBuf[9818] = 256'hf8cc76cde9cd23cf9ed0cfd2dbd4c7d77fdaf9dcdddf95e20fe5f3e7aceadaed;
    decBuf[9819] = 256'hfeefb6f2c6f361f5acf578f6b5f6edf620f7f2f674f6b4f57af4abf2faf091ee;
    decBuf[9820] = 256'hadebf4e87be63be4c5e2f9e1bbe183e150e122e1a4e0e4df35df16df32dfb5df;
    decBuf[9821] = 256'heae065e2cae3c8e5a4e7d0e946eb9aecceed77ee76efbaf08af231f5aaf78ffa;
    decBuf[9822] = 256'h80fc90fd86fe3cfef8fdc3fc3afb3bfaf6f87bf77cf694f5c2f44ff4e6f387f3;
    decBuf[9823] = 256'h31f37af275f13bf0c0ee5bed16ec44eb84ea61ea41ea5eea78eaefea30ebb9eb;
    decBuf[9824] = 256'h7eec00edd6ed66eee8ee5fefcbef55f03df15af266f3a0f4c7f5d4f6c8f766f8;
    decBuf[9825] = 256'hf6f844f92cf917f98df8ecf755f7a4f6fef53cf550f434f38ef105f0d4ed5eec;
    decBuf[9826] = 256'h82ea4de9a5e872e8fde8d0e929ebcaec53ee1ef053f16cf26bf353f422f64ef8;
    decBuf[9827] = 256'heefa1dfef6019f06010bfd0ea5130718271dfa219c27ea2c1d33f338c53f5b44;
    decBuf[9828] = 256'h8548cb4a7c4b1c4c674ad9487f465c446a42f13fb13d103b97380e35d330d72c;
    decBuf[9829] = 256'h25275320e8191214c40e910866042002aefe8dfbb4f81ef6c4f3a0f1afef9fee;
    decBuf[9830] = 256'h4dee98ee74f09ff2d6f5aff94ffd8a01aa061c0a7d0e9d130f17711b6d1f0d23;
    decBuf[9831] = 256'h662565288f299f2a4d2a022a362901287826ad248222e11fb21cb4196d159512;
    decBuf[9832] = 256'hf50eaa0b8709ce060a05ca02bf00e3fe3cfc77fa37f8c2f6f6f5b8f5f0f5eff6;
    decBuf[9833] = 256'h34f8aff9e0fbebfd4f008f029a0476062608af097a0ba60db10f1512b0132615;
    decBuf[9834] = 256'h6a15a815001567142213a711dc0fb00d0f0b96085606b503a602af01cf000300;
    decBuf[9835] = 256'hc5ffacfe13fe88fdb2fdbffe84002c03a505e507c50891094a0a830a820b230d;
    decBuf[9836] = 256'h1c0ff8102413c5153e18221bdb1d0921082432258d25df259425d8251626be26;
    decBuf[9837] = 256'h5727cc26a52566238220901ecc1c1e1d691dbd1ef11f2920901fa91e821dc21c;
    decBuf[9838] = 256'h9f1c7f1cd61cf01c071d741dd61d771e391fbc1f751fdd1eb71de71b371aae18;
    decBuf[9839] = 256'h491705168a14bf120e11850f200edc0cb50b5c0a1709f3065304d90199ff24fe;
    decBuf[9840] = 256'hd0fc92fc5afcf3fc21fd4bfd25fdbcfc1efc8efb40fb87fbccfc26ff0b025106;
    decBuf[9841] = 256'h710be30e0412b9134715ce143c159f156417ff180a1be61ca01d681dcf1ce71b;
    decBuf[9842] = 256'hc01a001a0c19ef1749165014ec11ac0f0b0d920af7085606910452024600f2fe;
    decBuf[9843] = 256'h39fe91fd5efd19fc9efa07f88ef54ef3d8f194f1d2f17af213f39ef374f334f4;
    decBuf[9844] = 256'h6ef592f732faacfc47fe27ff6bff37fe1efdb9fbd1faaaf99ef864f73df6caf5;
    decBuf[9845] = 256'ha7f506f695f64cf794f727f777f672f57df41ff43bf4f2f4c8f591f614f75bf7;
    decBuf[9846] = 256'hc7f751f85df903fb8cfc8bfd73fe9dfe76fe53feb2fe7cff0301fd026105fc06;
    decBuf[9847] = 256'h7208b608fc077306a804f8026f017000e5ff67ffa7feb3fd18fcaef9caf612f4;
    decBuf[9848] = 256'h2ef098ed4dea29e8ffe6a4e69be77be847e901eac9e996e9aee887e714e7f1e6;
    decBuf[9849] = 256'h8fe792e811ea76ebbbec36ee35ef7af0a1f1faf23ff465f525f6d4f672f702f8;
    decBuf[9850] = 256'h21f97afa1cfc34fd67fddcfc61fb30f925f749f599f3f0f223f3aef381f48ef5;
    decBuf[9851] = 256'hc7f69af7a7f80ff9f0f8d3f850f839f879f8a0f96ffb16fe900074036605c005;
    decBuf[9852] = 256'h12065d061906db05a30570054205c4049d0435041504bf03a5032e0340022301;
    decBuf[9853] = 256'h7dff84fda8fb7cf9dcf617f5d7f2f7f12bf169f181f2e6f388f5a0f69ff72bf8;
    decBuf[9854] = 256'h55f82ef80bf82bf80ef828f840f881f80af917fa70fb11fd9afe99ffc8ff9dff;
    decBuf[9855] = 256'h2affabfd46fc48fae4f7a4f599f3bdf10cf013eebfec8aebe2ea49ea1beaf1e9;
    decBuf[9856] = 256'h17ea80eadeea6eebf1eb38ec22ec0fecb5eb44eb17eb25ebaaeb93ecafedbcee;
    decBuf[9857] = 256'hb0ef4ef0def0f8f06ff1dbf13df2def24af30ff36ef22af12cefc8ec88ea7de8;
    decBuf[9858] = 256'ha1e6e7e520e6b9e6b7e81bebffedb7f031f315f695f9d0fdcc017e07500ebb14;
    decBuf[9859] = 256'h911a6321f825ce2b1c314f377a3bc8409b45fd49d54c7550de5171514650824e;
    decBuf[9860] = 256'hf94aae47d5432c3f8a393c34092e33286121f61a75136a0eff07d40386feb3f9;
    decBuf[9861] = 256'h52f555f1bfee74eb2cea01e9a7e89de913ebffed7ff1baf5dafaacff0e042e09;
    decBuf[9862] = 256'h010ea313f118241f4f239d280f2c302f093296330f34c6329c31222f9a2b5e27;
    decBuf[9863] = 256'h6223b91e1719c913f70e5409060434ffd2fab2f540f21fef46ecb0e956e732e5;
    decBuf[9864] = 256'hcfe429e57ce5f1e645e87ae993ea92ebd6eca6ee4df131f5d9f93bfe5b03cc06;
    decBuf[9865] = 256'hee09a30b300db80c260d890de40d360e810e3d0e080d9e0a1607da02bbfde8f8;
    decBuf[9866] = 256'h46f37cef0aece9e833e7a6e54ce303e2d9e0c9df77dfc2df8ee03ee237e49be6;
    decBuf[9867] = 256'h80e938ecb2ee96f115f560f85efbdefe29022705e007590a990ca40e700f2910;
    decBuf[9868] = 256'hd2106b115312791386143415541551148c12dc10530f540e250e500ec30ea00e;
    decBuf[9869] = 256'h410eb10d630dda0df30e991092126e14a3152c17c517ac18d319931afc1adc1a;
    decBuf[9870] = 256'h4c1a9619c0183018ad17d81662153113fb0f210c820837053902470019fd3ff9;
    decBuf[9871] = 256'ha0f573f0a1eb80e8a7e519e4b0e21ee381e327e379e3c4e390e440e639e825eb;
    decBuf[9872] = 256'ha5eeeff1c9f568f9a4fda0013f058a08880b080f621185133e1602189e19131b;
    decBuf[9873] = 256'hdf1b991cd11c9e1c6f1c451c391bb9192217f3131a10710b1007130374ff29fc;
    decBuf[9874] = 256'h2bf972f644f345f0c6ec6cea6de743e633e586e5d0e59ce64de8d6e9a1ebd5ec;
    decBuf[9875] = 256'heeed21eef3edc8eda2ed50ee6defc6f00bf2def2b7f209f22cf19cf082f099f0;
    decBuf[9876] = 256'h06f119f178f034efd9ec99ea63e740e587e278e181e036e002e137e24fe3e8e3;
    decBuf[9877] = 256'hd0e44fe575e523e640e7e6e850eb8fed9befeff023f2ccf2cbf36cf5f5f626f9;
    decBuf[9878] = 256'h31fb85fcbafdf2fd59fdcefc50fc43fb09fa8ef85df6bcf343f15eee6deca8ea;
    decBuf[9879] = 256'hb2e9d1e805e84ce714e77be6f0e51de55de4afe311e3bbe26ce284e21be3cce3;
    decBuf[9880] = 256'hd1e4c5e5a3e6f9e647e75fe7a0e778e8eee9b9ebe4ed5aef26f0e8ef60eefbec;
    decBuf[9881] = 256'h59eb41eaa8e9d6e9ace9d2e9afe950e9fae8e0e8c8e834e9e5e98bea23ebd3eb;
    decBuf[9882] = 256'h1bec5becbeecacec9becc8ec0bedc0ed48ef22f2a1f5ecf810fb01fd11fe63fe;
    decBuf[9883] = 256'haefe6afea7fe6ffe3cfeb1fd36fc6bfac4f74af5c1f168ef69ec78eab3e8bce7;
    decBuf[9884] = 256'h72e7b6e778e7b0e717e78ce662e6d5e683e7a0e8ace915ea74ea91ea77eabeea;
    decBuf[9885] = 256'h80eba0ec93eef7f0dbf393f6c2f9c0fc40008b03ae0567087609c809e8080c07;
    decBuf[9886] = 256'h6504eb0107ff16fd51fb5afae5f881f641f40bf10cee8dea42e71ee52de368e1;
    decBuf[9887] = 256'h72e091dfc5de03df3bdfa0e0e5e10ce318e452e579e61fe818ea7cecbceec7f0;
    decBuf[9888] = 256'h1bf250f3f9f392f4d6f5fdf60af8fef85df979f9c8f93ffa01fb84fb6cfbd5fa;
    decBuf[9889] = 256'haef933f868f6aff596f4fdf372f34bf2f2f051ef38ee05eeedeebcf063f3ddf5;
    decBuf[9890] = 256'hc1f8b3fa2cfd6cffa2025707f90c4712db19e61e5225272b7530a9367e3c4840;
    decBuf[9891] = 256'h7c46fc48c64c764d574fc54e4a4fe04d734dba4a4148144417406f3b0d371133;
    decBuf[9892] = 256'h682e472b4b27a222411e21194e14ed0ff00b510806050802160007ffb4fe95ff;
    decBuf[9893] = 256'he90014034b064909020c300f0a13a916e51ae11e7721d123f525e627f628912a;
    decBuf[9894] = 256'h072c5b2d142e2d2f602fd42e022ea82c4e2a6927ea239f20a11de81aba17bb14;
    decBuf[9895] = 256'h3c11f10d3d091b061f0289ff10ffa3fe06ff16006800de01aa025a045306b708;
    decBuf[9896] = 256'h9b0b8d0d510fa40fee0f3210ec10041269135114cf14f614d314f3140f159215;
    decBuf[9897] = 256'h3816231623151813e20f2e0b0c0810047a011000a3ff78fe69fdcefbedfa21fa;
    decBuf[9898] = 256'he4f98cfa8bfbd0fc4bfe1600c601bf039b054208bc0a450e8f11b3136b163018;
    decBuf[9899] = 256'hcb19411b1d1dcd1e56205521e021b621f620761fab1d801bdf18b015b212c010;
    decBuf[9900] = 256'h470e500dda0b960b590b210bee0abf0a410a670a160b320c250e01102d123814;
    decBuf[9901] = 256'h1416c417bd19991bc51d3b1f0720c020692102228d220b237e23162338228920;
    decBuf[9902] = 256'he21d681b84180415c910cd0c2408c303c6ff1efbfdf700f461f007eebeeccdea;
    decBuf[9903] = 256'h72eac5ea0febdbeb10ed99eecaf0d5f2c1f57af8a8fba7fe260271054a09f30d;
    decBuf[9904] = 256'h55122d15c4172d19761ad91ae91b3b1c861cca1c8c1c731b0e1a101834168414;
    decBuf[9905] = 256'h6b130612c210f20e420dd90a99088e062a04ea0149ff85fd45fbcff903f94af8;
    decBuf[9906] = 256'ha1f76ef740f76af7ddf75df98efb2ffea8004302240368032a038202e9010101;
    decBuf[9907] = 256'hdaff34fe3bfcd7f9f2f601f587f291f1b0f0e4ef2bef12ee13ed72ebe9e91ee8;
    decBuf[9908] = 256'he9e6d1e56ce484e306e3dfe28ee368e554e8d3eb0ff0e8f27ef5e7f630f893f8;
    decBuf[9909] = 256'h58fa97fcceffcc0285059406e6069c0658069e0566059905c8059e05de045e03;
    decBuf[9910] = 256'h2d018cfe13fc8af830f632f379f000ee09ed29ec6decaaec72ecd9eb4eeb7cea;
    decBuf[9911] = 256'h08eae6e905ea95ea4cebf2ebe0ecbdedc0eeb4ef13f069f04ff0d8ef6cefe3ee;
    decBuf[9912] = 256'h66eef4ed52edbaecbbebc7eaabe951e869e797e6d7e528e54be4bbe339e3f1e2;
    decBuf[9913] = 256'h07e369e3e6e358e484e45ce407e4fce356e40ce594e6fde899ea0eec62eda0ed;
    decBuf[9914] = 256'h49ee48ef2ff0fff1aff3a8f5fcf6b5f75ef891f879f9f7f9b7fadafa7bfa3ff9;
    decBuf[9915] = 256'h6ff7bff5a6f4a7f31cf346f320f3b7f219f2ddf0b6ef5dee75ed4bed24ed8ded;
    decBuf[9916] = 256'h2bee2eefdcefbaf0bcf1b1f28ef31ef46cf484f499f486f4dff451f5f3f58bf6;
    decBuf[9917] = 256'hedf6dbf669f6c7f504f582f40bf4caf38ff312f33ff275f18af0adef1def9bee;
    decBuf[9918] = 256'hf4ed5dedd4ec56ec46eccbecd7ed30efd2f0eaf183f255f2d7f117f1aef0d1ef;
    decBuf[9919] = 256'h7bef95efacef19f0a2f01ff1b1f162f2d9f245f380f36ef3dcf204f2c7f04cef;
    decBuf[9920] = 256'h4deec2ed44ed1dedb5ecd7eb9beacce81ce793e52ee446e31fe25fe16be04edf;
    decBuf[9921] = 256'hf5dd0ddde6db26db78da5bd94fd85bd7bcd6d9d6f9d79fd908dc91dfdbe2dae5;
    decBuf[9922] = 256'h59e995ed91f13af69bfa98fe4003a207c20cf512cb18191eeb228d28572c2a31;
    decBuf[9923] = 256'h4b342437c43a1d3d663e5740b240bb3f453e593bda37ae32db2d79295a24871f;
    decBuf[9924] = 256'h251b291781121f0eff082c04cbffabfa39f718f43ff1bbf033f17bf26df4e6f6;
    decBuf[9925] = 256'h26f931fb0dfd39ff44013004b007eb0bc40e6412ae15d217fc18c11a5c1c3c1d;
    decBuf[9926] = 256'h901e40205921f2217d22532293219f20431fa21d891c8a1b461a1f1979177f15;
    decBuf[9927] = 256'ha313fc10830e9e0bad099d08a7075c07a00762079a076707dc065e0637065a06;
    decBuf[9928] = 256'h3807e7088e0b080ea30f1911d5101b10930ec80c930b0a0aa508a706bb030201;
    decBuf[9929] = 256'hd4fdd5fae4f81ff729f6def512f562f368f18cef61ed80ec3cecf6ec7feee4ef;
    decBuf[9930] = 256'h85f19ef29df328f44ff55bf6dbf740f928fafafabafbf4fcc3feef0090030906;
    decBuf[9931] = 256'ha507ef0723076a06c205f505390760086d090409690700051c0263ff54fea6fe;
    decBuf[9932] = 256'h86ff520087019f0238037d04a106d709d50c1c11f5138b16f4173d19671a771b;
    decBuf[9933] = 256'hb71d5720d1226c24b72473243e234521e11e461da51a2b1847158f12600f620c;
    decBuf[9934] = 256'h700af70712055a02c1fd60f963f5c4f179ee31edcdec73ecc5ec10ed54ed0dee;
    decBuf[9935] = 256'hb5ee1af0bcf145f376f581f76dfa25fd0901a804e408bd0b5c0fb611d9139216;
    decBuf[9936] = 256'h0b194b1bc11c8d1d4f1da71cdc1ab0180f1696135611e00f8c0ed30d9b0dce0d;
    decBuf[9937] = 256'hfc0dd20d120d1e0cc20a7e0903086a073b0711073707a007c00716089908e008;
    decBuf[9938] = 256'h21095c0902092f08f3067805ad03fc01730074ff8dfe66fd0cfc0efa32f88bf5;
    decBuf[9939] = 256'hc6f32bf220f044ee18ec77e9fee6bee4dee39ae3cfe458e623e857e98fe95ce9;
    decBuf[9940] = 256'h2ee958e965ea70ec3cf0dbf326f724faddfc56ff96013704fb053b081b095f09;
    decBuf[9941] = 256'h9d09650998096a0994092109b808db079e0623055803a801afffd3fd23fc9afa;
    decBuf[9942] = 256'hcff89af711f646f496f20df142ef92ed09ec0aeb7feaa9ea69eb5dec3aed3dee;
    decBuf[9943] = 256'ha6ee86ee30eee1ed9aeddbed64ee05ef9defd7ef7eefecee14ee4bed94ec1dec;
    decBuf[9944] = 256'h2feb13ea6ce8e4e619e5e4e3ace3dfe3c7e442e641e729e8fbe8bbe924eac2ea;
    decBuf[9945] = 256'h8beb76ec93edecee8ef087f263f413f60cf860f919fac2fa5bfb89fb07fc7bfc;
    decBuf[9946] = 256'h29fd88fddefdf8fde0fda0fd8cfd9efdaefdbdfd44fd51fc46faa5f776f453f2;
    decBuf[9947] = 256'h61f09deea6ed5bed8fec52ec19ec4cec91ed60ef8cf102f356f40ff547f5e0f5;
    decBuf[9948] = 256'hc8f69bf7f4f8dcf95afa34facbf92df9d7f889f841f8d5f74cf787f6d0f52af5;
    decBuf[9949] = 256'hbef483f44ef4fcf378f3b3f230f2baf122f199f08def33ee35ec59ea24e9ece8;
    decBuf[9950] = 256'hebe98debf6eddaf0ccf2dbf32ef4e3f317f35ef2b5f182f154f1d5f062f03ff0;
    decBuf[9951] = 256'h20f0b0f066f10df24ef2ebf1dff086ef41ee17ee8aee7eefdaf0c2f141f21af2;
    decBuf[9952] = 256'hf7f1d8f12ef2e5f2eaf398f479f476f3f6f191f04defceeea8eecbeeebeeceee;
    decBuf[9953] = 256'h7fee38ee4eee3aee70eee2ee49ef11f0c1f168f4e1f66afab5fdb30033048d06;
    decBuf[9954] = 256'h8b090b0d650f3e13d5151f191e1c0f1e8920c822d42438277729182c922e7631;
    decBuf[9955] = 256'h2e34a8368c397e3b8d3cdf3cff3bab3afb3802372635fa32ef307b2d302a3227;
    decBuf[9956] = 256'hb2235821351f0a1efb1ca91c9d1ac1181a16a1130512bb110f13bf142817c318;
    decBuf[9957] = 256'hcf1a231c571de01edf1f2421a2217c218820ea1f5a1f741fa920242289237124;
    decBuf[9958] = 256'h4724d4236b23cd227722c522ad224122b821ac20521f0e1ee71cda1ba01a2519;
    decBuf[9959] = 256'h5a172e152313bf10240fae0de20ca40c6c0c9f0c2a0dfd0d700e1e0f7d0fd40f;
    decBuf[9960] = 256'h22106910d51086112c129812ac12e7115f10660e8a0ce3091f0883063906f505;
    decBuf[9961] = 256'h3206fa0561051d044d029d00a4fe50fd97fc5efc91fc1dfdeffd62fe11ffafff;
    decBuf[9962] = 256'h05008800fe00c101ac02c903d5040f063607f6077609410bf10c5a0ff6106b12;
    decBuf[9963] = 256'h371375133d130a137f1255122e120b12ad119011aa11f111b4129f137c14d314;
    decBuf[9964] = 256'hed14a5149014cb148f15af160818f018c3199c197919db18be180d19b319a11a;
    decBuf[9965] = 256'h3f1b951b131bde190f18e315d813fc114b10520efe0c4e0bc509fa074a065104;
    decBuf[9966] = 256'h750249003efedafb3efac9f885f8cbf704f837f865f83bf87bf741f61af5a7f4;
    decBuf[9967] = 256'hcaf4e7f526f866fa07fd80ffc001a002f403ad045605ef05d706550715083808;
    decBuf[9968] = 256'h9708ed08a4094a0ab60af10a980aa409df072e063504e1022802f0012302f401;
    decBuf[9969] = 256'hca01be000f0032ffdcfec2fed9fe98fe36fe72fd87fce8fb59fb0afb94faa6f9;
    decBuf[9970] = 256'h4af8a8f620f5bbf3d3f2a9f2cff238f3d6f39ff422f569f553f5f1f409f4adf2;
    decBuf[9971] = 256'h68f1edefeeee63ee8dee4def41f01ef1aef131f219f203f217f205f2d4f150f1;
    decBuf[9972] = 256'h67f04bef8bee22eec0ee36f001f22df4a3f5e7f52df5a4f3d9f129f0f1efbeef;
    decBuf[9973] = 256'ha6f021f2ecf39cf525f7f0f825facdfa9afa0ffa3df930f8c7f726f8eff872f9;
    decBuf[9974] = 256'h8af971f831f6f1f3bbf098ee34eedaed2cee0cef50ef12ef4aef17efa3ef75f0;
    decBuf[9975] = 256'h9cf079f0dbef9eee23ed24ec99eb6feb95eb72eb95ea1fe9eee6e3e47fe2e4e0;
    decBuf[9976] = 256'h04e0c0df82dfbadf53e03be10ae3bae4b4e608e8c1e889e88ae7e8e55fe460e3;
    decBuf[9977] = 256'h8fe3b9e3c6e474e594e577e591e5d8e59be6eee733e95aea80ead2e976e831e7;
    decBuf[9978] = 256'h0be697e5bae558e6afe6c9e623e68be529e517e5cae5ffe626e8e5e84ee96ee9;
    decBuf[9979] = 256'h8ae941ea76eb45ed71efe7f03bf279f241f20ef2dff1b5f1dbf1fef11ef201f2;
    decBuf[9980] = 256'hb3f10df175f03af028f039f00cf094efc1eebeed84ec06ec46eb23ebc4ea34ea;
    decBuf[9981] = 256'hb2e96be9abe9abeab6ec56efd0f1b4f4dff5eef69cf6e7f62bf75ff8e8f919fc;
    decBuf[9982] = 256'h8ffde3fe21ff59ff26ff9bfe71fefefd09fdaefbc6fa9ff9dff876f817f8c1f7;
    decBuf[9983] = 256'hd6f67af57cf3a0f1f0ef47efaeee80ee56eec9eeecee8aefc6f041f20cf438f6;
    decBuf[9984] = 256'haef702f9bbf9f3f9c0f9eff9c5f99ef9c1f962f9d2f8e7f7cbf6bef510f5f0f4;
    decBuf[9985] = 256'h46f531f60ff7d8f726f83ef8d2f721f74cf60ff5e9f38ff24bf124f064ef41ef;
    decBuf[9986] = 256'ha0efdcf0abf2d7f478f7f1f931fca7fd83ffb8004102a603470540079408c909;
    decBuf[9987] = 256'h710a0a0b950b140c870c7b0d190ea90ec30e7c0e100ead0d9c0d0d0ecd0eb80f;
    decBuf[9988] = 256'h9610ec109d10980f190e4e0c9d0aa408c80618051f0353029a0142020d043906;
    decBuf[9989] = 256'hd9089e0a390c190dd50c130ddb0c740dff0dd20e920ffa0f9b0f450fc30eda0e;
    decBuf[9990] = 256'h720f7110ab11d21245136813091379128e11b010e70f940e4f0d280c1b0bf90a;
    decBuf[9991] = 256'h970b990c5f0e0f1098119712dc13ae146e15d7157516051753176b1780174517;
    decBuf[9992] = 256'hc8167716d51569150715d114a01491143414c7135f13cc121c12a5113911d710;
    decBuf[9993] = 256'h7d102c108a0f9c0e400d420bde089e062805d4031b0353038603b5033304a604;
    decBuf[9994] = 256'h9a0578062708530af30c221045123714fb154e1603163715f9143115ca150f17;
    decBuf[9995] = 256'h3618f6185e19bd19131a2e1a161aaa19ab18e51635153c1360112b10a20ed70c;
    decBuf[9996] = 256'h270b9e0939080b083508a80811096f098c09db09810a9a0ba70c9b0dfa0d6a0d;
    decBuf[9997] = 256'hb30c7e0b570afe08b9073e06d9044e04cc04d90513078e082709f908d2072c06;
    decBuf[9998] = 256'hc2032702b1005dff20ffe7feb4fe29fe57fd4afc9cfbbbfb4bfc9ffd87fe5cfe;
    decBuf[9999] = 256'h50fd45fb0ef8ebf587f597f6d7f877fb3cfdd7feb7ff8300b801d102d003fe03;
    decBuf[10000] = 256'h80032602e2000f008200bc0137039c042705a90403039a005afe4ffcfbfac6f9;
    decBuf[10001] = 256'h1df9eaf8bcf8e6f8a6f9e0fa5bfc8cfe020056010f02d7013e01b30089006200;
    decBuf[10002] = 256'h3f00e1ff17ff60fe78febdffbb01970347057f058004df0256018bff56feaefd;
    decBuf[10003] = 256'haffc6afb97fa24fa8dfaaafb50fdd9fe3e00c9009f00780010002f004c003200;
    decBuf[10004] = 256'h2dffadfd7cfb71f9a5f867f860fac4fc4d00a702ca042e05d304dc03fc02b802;
    decBuf[10005] = 256'h7103aa03dd0351037f0272010a01a801e4025f045e0530055d0404036201d9ff;
    decBuf[10006] = 256'h0efee3fbd7f973f734f528f3e4f222f33bf43af57ef6a9f682f68ef532f4eef2;
    decBuf[10007] = 256'hc7f154f131f1cff1d2f251f482f623f99cfb38fdadfe79ffc0fe18fe19fd31fc;
    decBuf[10008] = 256'h5efb9efaf0f913f949f85ef7c0f66af650f638f622f6e8f523f538f45af3cbf2;
    decBuf[10009] = 256'hb1f2f8f264f3edf38ef451f570f616f880fa1bfc91fd4dfd18fc1ffabbf77bf5;
    decBuf[10010] = 256'h05f4c1f37bf493f55ef793f81cfa81fbc5fcecfdf9feedff0d00b6ffcbfeeefd;
    decBuf[10011] = 256'h25fda2fc8afca0fcdbfcedfcfdfc29fd87fddcfdfdfda3fdedfc65fbdcf977f8;
    decBuf[10012] = 256'h8ff7bdf649f627f646f663f67df695f6d6f638f7b5f768f80ef9d1f91ffa37fa;
    decBuf[10013] = 256'hcbf91af974f8dcf7c9f746f83af9fffa34fc4cfd19fd8efcbcfb48fb6bfb49fc;
    decBuf[10014] = 256'h4bfdfafd19fe50fd65fcc7fb57fcdffd48002c031e052d063605c103e501b9ff;
    decBuf[10015] = 256'haefdd2fb2af9b1f6cdf314f150effdee73f0d7f2bbf574f838fa2ffbe4fa28fb;
    decBuf[10016] = 256'he2fb4bfe2f01af04090776074c06d203ee00fcfeedfd3ffef4fdb0fd7cfc83fa;
    decBuf[10017] = 256'ha7f872f73af7d3f7bbf88df900faddf9fdf900fb7ffc16ff9001d003db05b707;
    decBuf[10018] = 256'h6709f00a550c9a0d6c0e2c0f4f0ff00e9a0e170e420d780c8d0b710ab1090209;
    decBuf[10019] = 256'h64080e08f4076b085809330b970d7b103413ad15ed1763192f1ae81a201bed1a;
    decBuf[10020] = 256'h621a3b1995172b15ec12b50f920da00bdc09d30a480c240e501030117411bb10;
    decBuf[10021] = 256'ha30f3e0e0f0ee50d580ec10e200f760f95103b12a5148917421a511ba31bc31a;
    decBuf[10022] = 256'he71840167b14e0120012bc11fa11a212a1132c14aa141e1540151e165a178118;
    decBuf[10023] = 256'h4119641908180a16a613c110090e440c050af9071d066d04e402e501b701e101;
    decBuf[10024] = 256'hee026d049e06aa08fe093b0a93099408f3066a056b04e0036103ee0240022301;
    decBuf[10025] = 256'hcaff85fe5efdebfc0efd2bfe1d008102c104cc062008e3073a07d505d703fb01;
    decBuf[10026] = 256'h42019a00670095006b00f8ff8ffff1fe9bfe4cfe64fea5fe7dfff30024035a06;
    decBuf[10027] = 256'h330ad30d1d1141136b14c614cf1359128d115910400fa70ebf0d440c790ad207;
    decBuf[10028] = 256'ha304a501ecfe73fc7cfbc7fb93fcbffe5f018e04b1066a092e0bca0c3f0e830e;
    decBuf[10029] = 256'h460e9d0dd20b220a29084d069d0414037d0003fe1ffb66f8a2f650f69af6eef7;
    decBuf[10030] = 256'h23f9acfa77fc27feb0ff1501b702cf039a05cf06e8078108f50726067f030501;
    decBuf[10031] = 256'hc6fe50fdfcfbc7faaef97df772f596f361f2b9f152f23af3b5f4e6f6f1f8ddfb;
    decBuf[10032] = 256'h96fe0f01ab02200464041e05c6059305ab04330205ff06fc15fa05f9b3f868f8;
    decBuf[10033] = 256'h9cf7ecf563f430f4d1f5abf864fbddfd8bfd15fcc1fa8cf9c4f9c3faabfb81fb;
    decBuf[10034] = 256'hdbf972f732f552f496f44ff5f7f52af69ff524f4f3f152ef24ec4ae8abe460e1;
    decBuf[10035] = 256'h3ddfd9dee9df84e18fe3f3e533e83eea92eb4bec13ece0ebf8eaceea8eeb99ed;
    decBuf[10036] = 256'h3af0fff151f2dbf0ffee58ec48ebf6ea41eb0decc6ec6eed07ee4cef1ff092f0;
    decBuf[10037] = 256'h6ff092ef8feee0ed82ed9eedb8ed71ed30ed1ded9aed8eee0df00cf1def0b7ef;
    decBuf[10038] = 256'h5eeebceca4eba5ea60e991e765e55ae316e353e36ce46be53de5c1e390e185df;
    decBuf[10039] = 256'h31deeade03e0cee17ee397e496e57ee6a5e7b1e8a5e983ead9eabfeae9e9ade8;
    decBuf[10040] = 256'h89e67ee4a2e264e27de3aee5b9e70de9cfe847e77ce5c2e4dbe50ce8adea71ec;
    decBuf[10041] = 256'h68ed48ee14ef40f176f450f8e6fa40fdaefd11fe6cfebefe09ff4dff93fe0afd;
    decBuf[10042] = 256'h3ffb14f99ef74af691f5c9f562f64af771f87df9a0f9c3f886f70bf60cf5def4;
    decBuf[10043] = 256'h5cf51cf685f665f648f663f6d9f645f70bf722f648f4e4f1a4efc4ee08efb8f0;
    decBuf[10044] = 256'hd1f1d0f2fef228f39bf3d5f44df731fbd0fe2a014d0378046803720266008afe;
    decBuf[10045] = 256'h5ffc53faeff7b0f50ff395f0b1edc0ebb0ea5eea3eeb92ecbeeec9f01df25bf2;
    decBuf[10046] = 256'h23f28af1a2f07bef22ee80ec87ea33e9f5e87eea15ed44f042f334f543f6f1f5;
    decBuf[10047] = 256'h3cf690f737fab1fcf0fe3bffe7fdbbfb1bf9a1f606f5bbf477f4acf5c4f68ff8;
    decBuf[10048] = 256'hbbfac6fca2fe5cff24ff8bfea3fd79fdecfde0fefcff090143021603d5038404;
    decBuf[10049] = 256'h64040e04f4036b04af050a084a0a2a0be60ab10998083109300ba40edf12b815;
    decBuf[10050] = 256'h4e18c71834199819f219a019eb19a719601a591ccd1ff9246b288c2bd7294027;
    decBuf[10051] = 256'h1422421d9f17d513c411e40f751003125d143618cd1a361c7e1d701f34211924;
    decBuf[10052] = 256'hd1269628e82847266422c41e791b311acd1973192119d618a219d71ab01d6920;
    decBuf[10053] = 256'h2d22db216520891e5e1ce81aa41a661a9e1ad11aa31a211b941b2c1b4e1a9f18;
    decBuf[10054] = 256'h73166814241462149a1467142213ff10f30eaf0ee40fdd1131136f13c7126211;
    decBuf[10055] = 256'hd710551148132415dd1535150413f8101c0fe80db00d7d0d4e0dd00c430d370e;
    decBuf[10056] = 256'h1110ed1122135a135b12ba10a10f6e0fb310da11e61238125e10720df209a806;
    decBuf[10057] = 256'h5f05c3051d061407f407b00772075a068d0675079809640d0c122e1506188217;
    decBuf[10058] = 256'h28152a12aa0e500c080b16099d066f0273feddfb46fdfa01dd08480f1e15e015;
    decBuf[10059] = 256'h30154f139a1115119d100a11e00f660ddd09930694033103aa0533096e0d4710;
    decBuf[10060] = 256'hd5115c11390f800c070a6c088b0747078507bd0756089b096a0b960d0c0fc80e;
    decBuf[10061] = 256'h9c0c3b0898024afd39fb99fa4efceeff5701c401d3ff59fdbefb9efc7afe2201;
    decBuf[10062] = 256'h9b03ed030d03b9010001a80173039f051507d1069c05a303c701890132029703;
    decBuf[10063] = 256'h7e045404ae02d5ff1cfd58fbaafbb5fda1005a036904720392023e01f7011003;
    decBuf[10064] = 256'hdb0419052003acff70fb97f80af792f6b5f8a7fa6bfc06fe7cffd0008002ea04;
    decBuf[10065] = 256'h85066507210771052702ecfdccf8f9f398efbfec3aecb3ecfbededeffcf0f3f1;
    decBuf[10066] = 256'h69f345f567f841fce9004b0500077c06130514025cffe2fc90fc70fd4cff7801;
    decBuf[10067] = 256'h19047304210416022aff71fc43f91ff767f483f0e4eca8e8f3e66fe6d8e7b1eb;
    decBuf[10068] = 256'h5af0bcf4b8f84efba8fda7009802f302fc01f1ff8dfd4dfbd7f983f84ef7e5f4;
    decBuf[10069] = 256'h01f248ef39ee8bee6bef37f0f1f0b8f01ff04ef020f1c7f2c0f414f648f761f8;
    decBuf[10070] = 256'hc6f921fcbcfd07fe2bfc8df8e4f3c3f00eef89eef2ef60f035ef71ed31ebbbe9;
    decBuf[10071] = 256'h87ea38eca1ee85f13ef46cf76bfa5cfc6cfd75fcfffaabf9e9f952fc37ff2801;
    decBuf[10072] = 256'h830143ff38fde4fb9dfc96fefa004c01d6fffafd4afcf3fc8affb80201040f02;
    decBuf[10073] = 256'h77fd15f919f594f4eef6c7fa67fec1002e01cb002501d3008800bcff0cfe32fb;
    decBuf[10074] = 256'h7af84bf528f3fdf1a3f1f5f16bf3bff4f4f5bcf557f458f204f1c7f0dff176f4;
    decBuf[10075] = 256'h3bf68df617f5b3f2bdf1c8f3c4f707fe3202f402e300c2fda2f891f6b0f442f5;
    decBuf[10076] = 256'hc6f54ef505f4a2f347f33ef449f625f8d6f97efa17fb45fb18fc25fd5efeddfe;
    decBuf[10077] = 256'hb6fe4efe70fd6efcbffba3fa49f94bf7e7f4a7f271ef73ecf3e8a9e585e322e3;
    decBuf[10078] = 256'he6e4cae783eab1edb0f0a1f2d0f5cef84efca8fecb006800a3fe63fceefaaafa;
    decBuf[10079] = 256'h5afce3fd7cfedafc01fa81f618f586f577f7f1f98cfb6cfc28fceafbe4fdd000;
    decBuf[10080] = 256'h4f049a07e2087f08ba06c30579053505f7046e03a3016e00c6fff9ff2700a9ff;
    decBuf[10081] = 256'h69fde1f9a5f5ccf23ff1b7f100f3f1f4b6f6f6f82cfc0500ae041009e80b760d;
    decBuf[10082] = 256'h0d0ce909f8073306e1052c060808330ad40c990e34101411581196113e12d712;
    decBuf[10083] = 256'hbf133e14ca134b121a10790db50b190aa408500796065e065d07b809410d8b10;
    decBuf[10084] = 256'h8a13b4145a1463138312c71205135c12c50f780aa6033bfdbafaf8f96afd8c00;
    decBuf[10085] = 256'h880415069d052f05930557073c0a820e5b11e8125214bf145c14b6146414ee12;
    decBuf[10086] = 256'h0210830c38091407b106c0075c093c0a800a420a0a0aa30aa10c050fe9111413;
    decBuf[10087] = 256'h2314d113f1129d11710f3b0c6108b9039800e2fe67ffc101bf043f08990abc0c;
    decBuf[10088] = 256'h200d7a0d280d870a59077f03d7feb5fb00fa7cf9f4f987f923f9c9f8bff935fb;
    decBuf[10089] = 256'h21feda00e901f2007dffa1fd6cfc14fd45ff7b029f049006eb063d071d08f909;
    decBuf[10090] = 256'ha10c1a0f5a110f11330f950bf507ab046203c6033f06db07e6093a0b6f0c680e;
    decBuf[10091] = 256'hcc10b013da148014f710da0a5a034afcdff50af5ccf53df99ffd54ffd0fe76fc;
    decBuf[10092] = 256'h78f986f796f8d5fa0cfe54ff2afefbfa47f625f394f22af584f782fa74fccefc;
    decBuf[10093] = 256'hc5fdd0ffcc03c9075609cf098608ce050904b703020446041103a700c3fd0bfb;
    decBuf[10094] = 256'h46f94ff89af866f99bfa24fc21ff1f029f05f9078b07610651055a04a504e904;
    decBuf[10095] = 256'hb4036b003efb6cf64bf3b9f234f2bcf173f0bbedf6eb92edf3f116fa1204c80a;
    decBuf[10096] = 256'he210fe11001340106b0fa10b2f080e0535029eff26ff94ff30ffd6fe28ff73ff;
    decBuf[10097] = 256'h4f01f603ba05c404f8003dfad2f3fcedb6eb67ec48eed9ee55eecdee3befbaf2;
    decBuf[10098] = 256'hd7f8adfe7f053f086a07a0038e016dfedbfd57fdeefbeff8a9f466ee3beaf5e7;
    decBuf[10099] = 256'ha5e8c6eb0af2dff72dfd9f00ffff26fd87f92df709f5dff384f3e9f1b3eefee9;
    decBuf[10100] = 256'h9ce5e7e375e5a1ead4f0fff4c1f511f530f3c2f358f684fbb801e305a5063303;
    decBuf[10101] = 256'h50fcbaf78ff3cdf2def4bff62df685f1e3eb11e550e27be145e518ea79ee0bef;
    decBuf[10102] = 256'h7eed24eb00e964e992ec6cf002f37bf357f111ed14e975e50ce479e4a4e5b3e6;
    decBuf[10103] = 256'haae7f5e7b1e76ae8f3e9f0ecc9f069f4c3f630f706f6f6f400f4b5f381f43af5;
    decBuf[10104] = 256'h72f5d9f44ef4ccf4bff6abf964fc73fdd8fb0cf85bf291ee1feb7fea10eba7ed;
    decBuf[10105] = 256'h01f024f2ddf40bf8c0fc22011e05b4072d08e4062c04b201cefe15fc32f880f2;
    decBuf[10106] = 256'h32edc1e9e0e795e93eeee0f3b2fa72fdf2ff30ffe1ff40ffd2ff5700deff96fe;
    decBuf[10107] = 256'hddfb19fac6f911fa75fc59ffa0039c073c0b960dde0eb40def0b0b095206d903;
    decBuf[10108] = 256'h3e02c800ecfeb7fd9efc37fd92ff77026804c304830222fe7ff8b5f4a4f285f4;
    decBuf[10109] = 256'h5ef706fc27ff00028502fd02da00afffebfd3dfe1dff810165041e0778078206;
    decBuf[10110] = 256'h0c05b8037a039304f805e006b5060f051603c2010002a80241035902e2fffefb;
    decBuf[10111] = 256'h5ff8f5f63ef8bdfb17fe60ff35fe52fab2f668f3d5f38ef671fa1aff3b02cd02;
    decBuf[10112] = 256'h3f01f5fdf6faccf926fac1fbf8fef60121037b032903740350057b0787093308;
    decBuf[10113] = 256'h9404d1fc0df502f017ef97f1e5f6b8fb98fd07fd70fa16f8a9f7effb3202b309;
    decBuf[10114] = 256'hba0ca40d240b5a07e8030802bd035306ad08f609590a690ba80d0a12ac17761b;
    decBuf[10115] = 256'he81e881f8c1be31601106b0b4007fa044a046902d70141ffe7fc9efb02fc7bfe;
    decBuf[10116] = 256'ha802a5063b09a40a370a0c096709020b0d0de90e270f9e0d6d0bf7093b0a670c;
    decBuf[10117] = 256'h080f3612a4127911b50fd10ca60b010cf70c6d0ec10f7111bb14e7191b20f025;
    decBuf[10118] = 256'hba296b2a4a272a22571df518f9145a111e0d22098c06220590050f095a0c590f;
    decBuf[10119] = 256'h4a115a1250133114851547152e1497111e0f820dcd0da90f501215140c152b14;
    decBuf[10120] = 256'h4f122410180eb40b2c08e104e301f1ff4c003003af06fa09f80cb10fdf12b916;
    decBuf[10121] = 256'h581aa31d361d7d1a30155e0ef2077205a801f80017ff85fe01fe5b007e023705;
    decBuf[10122] = 256'h46064f054403780231030b068b09d50c1e0e2c0cfe08240597032e029b02c603;
    decBuf[10123] = 256'hd504cc05420796084f09360839056001b7fcd6fa68fbf6fc40003f03f705bc07;
    decBuf[10124] = 256'h5709620bb60c700d370d060bd007d204a70302049d051307df07a10788062305;
    decBuf[10125] = 256'h3b041503550261014400ebfea6fd7ffc72fb0afbabfac8fa16fb8dfb4ffc3bfd;
    decBuf[10126] = 256'h57feb1ff52016b026a033b031402bb001aff01fe02fd77fcf8fb39fb44fa25fa;
    decBuf[10127] = 256'h28fb33fdfe009e040706bf04780058fbe6f706f6bbf763fc0602d005e1074107;
    decBuf[10128] = 256'h8b05fe03950202036603c00312045d04b1056107ea08b7085c062f020ffd9ef9;
    decBuf[10129] = 256'hfdf8b3fa5bff7c025505da058003f0fda2f8d0f3aef01df0a1f00af22ef4e6f6;
    decBuf[10130] = 256'habf846fabcfb88fc4afca2fba3fabbf991f96af9bcf860f7a8f4f0f12bf0d9ef;
    decBuf[10131] = 256'h4ff1c3f4fef81efe900171032605b3063b06f2040103d2ffd4fce2fad3f925fa;
    decBuf[10132] = 256'h70fac4fb74fd8dfe8cff5dff37fef7fb13f921f75df5c1f3e1f28df158f0b0ef;
    decBuf[10133] = 256'haff067f374f847fd28ff96feedf94bf4fdee8bebaae9f5e77ae801e84ae902ec;
    decBuf[10134] = 256'h50f19ef6d1fcfc0042039202f1016001e4015d02ef01feff1afc72f750f49bf2;
    decBuf[10135] = 256'h20f379f578f869fac4fa16fbcbfafff9d4f79df4e9efc8ecefe97cebc7ee57f4;
    decBuf[10136] = 256'ha5f916fdf7fe89ff16019e0056ffd6fbb9f5e4ef96ea84e825e9fdeb8bed03ee;
    decBuf[10137] = 256'hbbec02eaa8e943eba4efc8f78cff920253057d043702c5fee5fc2ffbabfa23fb;
    decBuf[10138] = 256'h6cfc08fcaefb6ef9cdf654f401f477f5dbf776f9c1f96df8bdf615f67af731fa;
    decBuf[10139] = 256'heafcf9fda7fd31fc65fb1efc88fe6c019702d200a5fc62f637f26deebced9def;
    decBuf[10140] = 256'h99f339f783fa82fd73ffceff33fe27fcc3f984f739f7f5f6aef7e6f7b3f785f7;
    decBuf[10141] = 256'hacf8ebfa19ff3804aa074b089506ed014bfcfdf68bf3aaf1f5ef67ee1deb1ee8;
    decBuf[10142] = 256'hf4e603e8d5ec69f479fbb9030d071008250750060a0459033a05cc055006c906;
    decBuf[10143] = 256'h5b06bf0638090a0edc127f18c51ab41892157310a00b7f08a605fd001bfadaf1;
    decBuf[10144] = 256'h4eec43e72de8aeeafcefcef4aff641f7c5f71ffa43fcc2ff1c02ae01bdffd9fb;
    decBuf[10145] = 256'h43f9cbf8eefa6efeb801dc03b102ed00f6ff41002d03ac06f7091a0cb70b3d09;
    decBuf[10146] = 256'ha2075707bb09e90d08137a165b18a6160f14b511b70e530eae0e4910fe0faa0e;
    decBuf[10147] = 256'h880bae070f04a502130376038604eb02df00f3fd02fc11fdf6ff7503b107890a;
    decBuf[10148] = 256'h170c8f0cd80d3b0e4b0f9d0fe80f2c10ee0f460fe10d290ba9076e0395001100;
    decBuf[10149] = 256'h6b024406ed0a0e0ec30f5111ba120214f41503170d16d612220ec009e7066306;
    decBuf[10150] = 256'hcc07ca0af50b4f0cb40a3e09ea07a4089d0a790cae0d560e230ede0c630b9809;
    decBuf[10151] = 256'h6c07f705a304e004690634086909f20a8b0b160ce90ca90dcb0d6d0df70b2c0a;
    decBuf[10152] = 256'h7c08630764067c05ad038a00b0fc11f9b7f64af63bf8b5fa3dfe8801ab036406;
    decBuf[10153] = 256'hdd08c20b410f8c12af1413154e13210f010ace03a3ffd9fb89fc6afe66020606;
    decBuf[10154] = 256'h6008a8094509ea0898087809cc0a860bdd0ae0072c0389fdb7f622f2f7edb1eb;
    decBuf[10155] = 256'ha0e9bfe72de7c4e9ffed42f46dfd87034b0b520e3d0f670e210cb008cf063d06;
    decBuf[10156] = 256'hb004460323016afea6fc54fcc9fdb50035048f06d707ad069d05a704f1044506;
    decBuf[10157] = 256'hf6079e086b08e0070d07e70695073308dd0755060b03fefbf2f65df287f1cdf3;
    decBuf[10158] = 256'h3ff7a1fb7afefefe77ff2efe04fda9fcfbfc46fd7afccafa80f735f412f275f2;
    decBuf[10159] = 256'h85f30ef749fb22fec1012a03730464067407c6077b079f05f802caff81fe1efe;
    decBuf[10160] = 256'he2ff22029803dc03220329014dff18fe51feb6ff5701e0024504d00452044503;
    decBuf[10161] = 256'hc5016000d5ff57ff7dff15ff79fda0fa20f7d6f3d7f0e6ee6cec2cea8ce7c7e5;
    decBuf[10162] = 256'hd0e446e632e979ed75f114f57ef6c6f72af884f81ffa6afaaefafef894f6b0f3;
    decBuf[10163] = 256'hf8f09df0eff0fbf2d7f490f577f4acf278f1b0f17bf39df69cf98dfbe8fba8f9;
    decBuf[10164] = 256'h72f64ef4ebf3faf496f636f9fbfaf2fb3cfc80fcbefc47fe12003e02b4037003;
    decBuf[10165] = 256'hc80030fc4df5e2ee0ce942e531e391e2ffe184e2ede310e61eeb51f1d1f8e1ff;
    decBuf[10166] = 256'h7704f706b9070907a9073b08b6077b035bfec7f6b7ef21eb4cea16eee9f2cbf9;
    decBuf[10167] = 256'h8cfc0cffc6fc54f973f7bef542f68df98cfcd200ab034a07a409c80bf20c980c;
    decBuf[10168] = 256'h580a8c06e40182fda9fa1cf994f9b8fbe2fcf2fd9ffd2afc4efa9df814f715f6;
    decBuf[10169] = 256'h2ef55bf44ef35af23ef131f00ef06af122f42ff902fe63026006f6085f0acd0a;
    decBuf[10170] = 256'hbe0c830e7a0f990e250b080588fd78f60df08ded47eb58ed39ef35f3def73ffc;
    decBuf[10171] = 256'hf5fd82fffaffb2fe87fd0efb73f9fdf7a9f6e7f6fff796fa7afe19027304e104;
    decBuf[10172] = 256'hb603f201b2ff3cfee8fcb3fbbaf9cef688f2afef19eda0ec0eed38eefdefe1f2;
    decBuf[10173] = 256'h27f747fc7b02a5066707b7069603bd0027fe9ffee7ff4b0086fefefac2f6eaf3;
    decBuf[10174] = 256'h53f1cbf139f29cf2acf347f5e8f716fbf0fe7d000500e2fd29fb1afab5fb81ff;
    decBuf[10175] = 256'h20036b06fd05d3045902be009e016a0223039b019efe0ef9c0f34ef0aeef1cef;
    decBuf[10176] = 256'hb3f10df430f6b0f909fc52fd7cfe8cffcc019705400ae20fac13bd155e16ef16;
    decBuf[10177] = 256'h6b16e3169b15e212950d3f057bfd6ff8aff52ff875fae7fd87fef6fd71fd08fc;
    decBuf[10178] = 256'h9bfb8cfd060033042f08d80cf90fae112a11b1108e0e9c0c230a3e078604a200;
    decBuf[10179] = 256'h0cfeb2fb45fb36fd650063038e04e80496044b041705d005e9061c07a7072209;
    decBuf[10180] = 256'h1f0c8a12f518201d661ff41b92174f11cf0e0d0ebd0ede1194131814af124212;
    decBuf[10181] = 256'h171127121d13d3120712e40e0a0b74081a06ac0510066a06bd06dc0500045002;
    decBuf[10182] = 256'h18027d033506090c34107a12ca11e90f100d7a0a1109a308070961090f095a09;
    decBuf[10183] = 256'h9e09d20aeb0b840c0f0de50c720c950c330d6f0e3e106a12e013341572151a16;
    decBuf[10184] = 256'h4d163517b018151afd1a7f1a3f181214f20e1f0abe0508047b02020270020c02;
    decBuf[10185] = 256'h670215025f02a3025d037504da05d8073c0a210dd90f53123715281783178c16;
    decBuf[10186] = 256'h81149511a30fdf0d8d0dd70d1b0e6b0c2109f503c2fd97f9cdf51df5fdf6b3f8;
    decBuf[10187] = 256'h40fab8fa26fb17fdfb00ac067e0d1412ea17ac18fb17da1425138e101610a90f;
    decBuf[10188] = 256'h450f360e9a0cba0b660a280a600a2d0ae9087106230151fae6f311eecbeb1aeb;
    decBuf[10189] = 256'h7cefbff595fb6702fd067d093f0a8e096d067102c8fda7facef753f89dfb77ff;
    decBuf[10190] = 256'h1f044107f608830afc0a690bcd0b080a2407170244fda2f7d8f3c7f167f21cf4;
    decBuf[10191] = 256'hbcf7e8fcba01dc0491060c06a3048002c7ff4efd0efb03f917f65ef39af1a3f0;
    decBuf[10192] = 256'h19f205f5bdf737fa2dfb78fb24fa6bf9c3f82af8fbf7d1f711f71df67ff59cf5;
    decBuf[10193] = 256'heff64af9d3fc1e00f7038e061506f203e4feb1f8dbf211ef9feb7ee8a5e506e2;
    decBuf[10194] = 256'hacdf88ddecddcfe181e753eebef4e9f82ffba1fe8405ef0b6f137b1865193a15;
    decBuf[10195] = 256'h680efd07d20310036002c001a0fc0cf5fced91e711e5d3e545e9a6eda3f14bf6;
    decBuf[10196] = 256'hadfaa9fe520373062808ad082509b708c606970308fe36f7cbf04bee0def7ef2;
    decBuf[10197] = 256'he0f6dcfa61fb07f9bff75bf7d5f95dfdb7ff25006cfd89f9f2f66bf7d8f703f9;
    decBuf[10198] = 256'h3ef7b5f389ee17ebb8eb90ee42f490f962fe84015c04ea054408b1088707c205;
    decBuf[10199] = 256'hde02b401590107012700c3fddefaedf892f81bfc56005304e00586038800cffd;
    decBuf[10200] = 256'hc0fcb7fd57006701150109ffb5fdfcfca4fda3fe75fe51fc86f8e6f49cf12ef1;
    decBuf[10201] = 256'hcbf025f18aef54ec7ae8e4e57ae49ee656e985ec83ef3cf26af544f9dafb34fe;
    decBuf[10202] = 256'h5800820147032b06720a6e0efb0f7410500e430970040e00effa1cf6baf177eb;
    decBuf[10203] = 256'ha1e553e0e1dc82dd5ae003e565e961ed09f26bf667fa1900e3035507f5074006;
    decBuf[10204] = 256'h9701f5fba7f6d4f173edbdeb39eba2ecebeddcef56f24cf32df481f5acf7e3fa;
    decBuf[10205] = 256'hbcfe5c02b504fe05d304c403290248017c003f0096ff31fed6fb97f921f8ddf7;
    decBuf[10206] = 256'h12f97bfbbbfd31fffdff3a00e300480246049a0553063a0509036900a4fe52fe;
    decBuf[10207] = 256'h5d00c1020105e1059d05ed03f401180068fedffcaefa77f79ef3feefc3ebc7e7;
    decBuf[10208] = 256'h30e5b8e425e517e7faeaacf07ef7e9fdbf0389073908d90824078e04340235ff;
    decBuf[10209] = 256'hb6fb5cf938f7d5f62ff76ff910fc3eff1803b706f30aef0e8f12e8147b14c211;
    decBuf[10210] = 256'h2a0dc808cc043e03c60234030902fa00bafe19fc0afbb7fa2dfc81fd43fd2bfc;
    decBuf[10211] = 256'h94f9cff7d8f6e4f8d0fb88fe0201af003affd6fc96fa20f954f816f8fef6cdf4;
    decBuf[10212] = 256'h2cf2b3efbcee5df1aaf600ffc406cf0b900e0f0cc106ef018dfdb4fa39fba2fc;
    decBuf[10213] = 256'h0ffdacfc32faf3f712f7eef88dfc5004140c1f11e01360111a0f470a6608d407;
    decBuf[10214] = 256'h5908d10889070904cefff5fc71fce9fce8ffd9019e034b036b02af026803f104;
    decBuf[10215] = 256'hbc067507ae0715072d065a059a047704d60412068e07f308da095c091c073804;
    decBuf[10216] = 256'h47023701d20209060709f90a530b5c0a7c09480a740c7f0ed30f9e0e550b0a08;
    decBuf[10217] = 256'h0b05a8040205f905ae055a04aa02920191028f04e305a5053c03b3ff68fcfbfb;
    decBuf[10218] = 256'hecfd66004a033b054b06e6071c0bd10f3314c4142e12020d6e055efe9efb1ef9;
    decBuf[10219] = 256'he0f9f1fb91fcfffb7bfbf3fb86fbb0fc75fe10001b020705c007a30b3a0e9310;
    decBuf[10220] = 256'hb712e1133c148e14ae13d211a60f700c9608ee038cff90fbf9f890f723f74df8;
    decBuf[10221] = 256'hc7fa07fd7cfed0ff8a0083025f048107a509960b3c0ba1096a066c03b300a4ff;
    decBuf[10222] = 256'hadfecdfdf1fb4af91bf6f8f3cdf2ddf3c1f607fb2700fa041b08ad081f07d503;
    decBuf[10223] = 256'h20ffbefa09f97cf7e5f808fbc1fd3a00d601b6020a04480480044d041e04a003;
    decBuf[10224] = 256'hc60375049105eb062f0802092809c00864071f065004a0021701180046006d01;
    decBuf[10225] = 256'had03da07d60b7f10e014b9174719dd1704145b0fb909e7027cfca6f6d4ef3feb;
    decBuf[10226] = 256'h14e7cee47ee59fe8bfedf2f373fb7e001405e90ab30e8613a7165d18cf16a311;
    decBuf[10227] = 256'h700b44022bfc9ff693f1a9f07ef140f251f4b3f8affc4f00a8021603eb01dc00;
    decBuf[10228] = 256'h8a006a0136027402cb019aff8ffd4bfdfbfed5015405ae0741078804a500fcfb;
    decBuf[10229] = 256'hdbf826f798f52ff4c2f35ef36ef4adf64ef9c8fb63fd43fe77fdbefca5fba6fa;
    decBuf[10230] = 256'hd5faa7fb01fdfffedb001002480249010400ddfeb7fe65ff43005f00d7fe8efb;
    decBuf[10231] = 256'h61f68ff1aeef1cefb3f1fdf4d7f876fcb200ae045709b80d91101611cb0d3b08;
    decBuf[10232] = 256'hed02bafc8ff849f699f57af752fafbfe5d035907e6086e084a069203630040fe;
    decBuf[10233] = 256'h15fd51fbfffab4fa80fb30fd29ff0501bf011601170076fe0cfc28f9a9f55ef2;
    decBuf[10234] = 256'h60effceec1f0a5f3ebf7c4fa52fcd9fb91fa2dfaf2fbd6fe8e015303a503c502;
    decBuf[10235] = 256'h710133012c0318069809010b6e0b7d09b8071d06fd0651088609be09f307d104;
    decBuf[10236] = 256'hf70058fd0dfac4f861f870f90cfb81fcd5fd13febcfebbffb901a5045d07b807;
    decBuf[10237] = 256'hc1068b038c00d4fd79fd70fe110120027202fd00a9ff7dfd9dfc49fb98f99ff7;
    decBuf[10238] = 256'hb3f4fbf136f040eff5ee49f075f240f6e9fa8b005504c7076708f9086b07f306;
    decBuf[10239] = 256'h860622061305d3029dff79fdddfda1ffce03cb074f08d707d80420025b00ad00;
    decBuf[10240] = 256'hb9020d04cf03f500affcd6f95bfab4fc44020e068009e0082a078b033101e8ff;
    decBuf[10241] = 256'hbefe44fc17f81bf47bf003f04cf159f68cfc62022c069e097f0b340db80d310e;
    decBuf[10242] = 256'hc30d600dba0db10e910fe5109612ce129b12b3118c10e60eed0c890a0007c502;
    decBuf[10243] = 256'ha5fdd2f8b1f51ff5a4f5eef8edfbdefda3fff5ff40009401c0036006da08750a;
    decBuf[10244] = 256'h95093107a8035d0084fcedf994f770f57ff324f3bff4cbf6b7f936fd8100a402;
    decBuf[10245] = 256'h5d052107bc08320afe0a3c0b940a63085706f303fd02470323054f075a09ae0a;
    decBuf[10246] = 256'h710ae808eb05110272fe09fdc0fb24fc33fdcefeda00c6037e06620a010e6a0f;
    decBuf[10247] = 256'hd80fad0e340cf4097e08b20774073c07a306020579031402cf0054ff23fd83fa;
    decBuf[10248] = 256'h09f86ef68ef54af50cf5f3f3c2f14cf080ef31f17bf4a7f919fd3a00cc005001;
    decBuf[10249] = 256'hb902b805c50a980fb9124b13bd11820d8609ef0686051905b5041005bd04dd03;
    decBuf[10250] = 256'h9903e002370238013affd6fcf2f973f619f4d0f234f3adf5daf9d7fd6d00c702;
    decBuf[10251] = 256'h3503d1020d0171fffcfd98fbb3f8fbf581f32ff30ff483f7bffbde00b1059207;
    decBuf[10252] = 256'h4709cc09440a8c0b450ebe105a120f12ab0f220cd808d905760585067c07f208;
    decBuf[10253] = 256'h26087e05500276fee0fb77fa09faa6f900faaef98efa6afc0800c306590b840f;
    decBuf[10254] = 256'hc20e110ef00a17088a061106c904d7023ffe9df84ff37ceedced6dee0df258f5;
    decBuf[10255] = 256'h31f9bffa28fcbafb57fb47fa50f99bf967fa9cfb95fde9fe27ffeffe56fee1fe;
    decBuf[10256] = 256'h0800fb01d7039004e703e802a401250199018d022b03810367034f0312049a05;
    decBuf[10257] = 256'h230788085908de0613056303da014101b600e3ff8afe8cfc38fb03fa5bf9c2f8;
    decBuf[10258] = 256'h93f815f855f7a7f64bf506f48bf2f2f17df2a1f46cf815fdb7028106f309140d;
    decBuf[10259] = 256'hed0f7210f90ffb0c2607fbfd70f5e4efdeecf3eb73eeb9f0caf22af298f11df2;
    decBuf[10260] = 256'h58f69bfc71023b06eb06ca03ceff2efcd4f942fa6cfb31fd28fe72fe2efee8fe;
    decBuf[10261] = 256'h90fff500f30247047c0544057903dbff32fb90f542f031eed1ee86f01df386f4;
    decBuf[10262] = 256'hcef5f9f608f8edfa6cfec600e9028602c10082fe0cfd50fd09feb2fe19fe31fd;
    decBuf[10263] = 256'hb6fbe9fb8afdd4000f050b0987081e074403a5ff4bfdb8fd7100ea022a050a06;
    decBuf[10264] = 256'h3e050a04f10258027001a1fffafc16f96ef44cf174eeefed58ef7cf1fbf446f8;
    decBuf[10265] = 256'h44fb36fd45fe98fee2feaeff6800a0000700c2fe47fdaefc39fdb1ff94033407;
    decBuf[10266] = 256'h7f0ac70b640b540a14080906a5036501c5fe96fbbdf714f3f3ef3eeeb9ed31ee;
    decBuf[10267] = 256'h55f046f275f573f8f3fb3eff61015303ad03ff03b50381043a05e2057b064d06;
    decBuf[10268] = 256'hce05a805cb056906bf060806a404a701cefd37fbcef961f98bfa50fcebfd61ff;
    decBuf[10269] = 256'hb500e9017203d704bf059505ef03a5006afc6df8cef465f3d2f3fdf42bf805fc;
    decBuf[10270] = 256'h9bfef500190343040806a30783084f091109a8061f03d5fffbfb6efaf5f93efb;
    decBuf[10271] = 256'h2ffd8afd37fd57fc8bfbc9fb71fc70fdb5fe33ff0dffeafe49ff1200fd00db01;
    decBuf[10272] = 256'h3102ae017a00a7ffe7fe0affe7ff2401f6011d026e011200cefea4feb0ffbb01;
    decBuf[10273] = 256'h870515078d074406c5026b0023ff4d005d010a0195ff31fd4cfa22f931fabafd;
    decBuf[10274] = 256'h0501030467045703600216026a03950536084609f308e8068404a001e7fe6efc;
    decBuf[10275] = 256'he5f88bf643f5dff459f7e2fa1dff1903a7042e04e602bb01ac00b5ff3ffe63fc;
    decBuf[10276] = 256'hbcf943f7f0f666f862fca5027b08c90d3b11db112610a10f470d6e09c50423ff;
    decBuf[10277] = 256'hd5f963f6c3f555f6e2f75bf8c8f865f855f7a7f788f874fb2cfe5b0159048405;
    decBuf[10278] = 256'h930641068c06c0058b047203a701f7ff6efea3fc6efbc6faf9fae1fb5cfdc1fe;
    decBuf[10279] = 256'h4cffcefec1fd87fc09fcc9fcbdfddafe4dffe4fec4fe1bff6e00100299030003;
    decBuf[10280] = 256'h480001fc05f86ff5e7f530f721f931fadef969f815f7cef7a7fa27fe72019503;
    decBuf[10281] = 256'hf903e9024e010301cf017f037805cc060108aa08dd080b0935095b09c409e409;
    decBuf[10282] = 256'h540900084905c9019dfccaf7a9f4d0f14cf1c4f1c3f442f87efc9d010f053108;
    decBuf[10283] = 256'hc2084709ed06c90411024c0056ffa0ff7c01a803b3058f074908a0073b06e003;
    decBuf[10284] = 256'hfc0044fe7ffc88fb69fcbdfdf1fe9affcdff42ff18ff3eff32008e0176024c02;
    decBuf[10285] = 256'h8c010c00a7fe63fde4fcbefce1fc40fd09fe91ff6a025c042006ce05ee048a02;
    decBuf[10286] = 256'h4a00d4fe08fe4ffd36fc6bfa37f9fff8fef958fc3dfff501ba035505cb061f08;
    decBuf[10287] = 256'hcf09770ade093d086305e40199fe9bfbe2f8d3f7c9f8d5fad1fef003c308e40b;
    decBuf[10288] = 256'h9a0d150dac0b8809d00656047201f3fdb7f9bbf52ef4b5f3d9f558f984fe5703;
    decBuf[10289] = 256'h78062d08a90740061c0464019fff04fe8efcb2fa0bf828f488f03dedd0ecc1ee;
    decBuf[10290] = 256'h5af3fcf8ceff6404e406a607f6065506e7067508de099508a406c00221ffb8fd;
    decBuf[10291] = 256'h4afdaefdbdfeb4ff69ff15fe5cfd24fd23fec4ffbd01110346045f0592050705;
    decBuf[10292] = 256'he0033a024000ecfe33fefbfd2efe16ff3d0049010f03bf044806e106b306e304;
    decBuf[10293] = 256'hc001e7fd47fafdf6b4f551f560f6fcf707fa6bfc06fe1100ed019e032605f106;
    decBuf[10294] = 256'h26083f09d809f00878064a0370ffdafc70fbb9fce3fd5d0054019e014a0016ff;
    decBuf[10295] = 256'hfdfd64fdeffd6aff350161030206c607190838075c05b5023c0045ff65fe21fe;
    decBuf[10296] = 256'hecfc63fb66f842f618f572f557f80ffb3efe86ff23ff5efdc3fb78fbccfc7cfe;
    decBuf[10297] = 256'h0500380050ff2afe6afd18fef2ffde0297055b07ae07f807b4076e081609e308;
    decBuf[10298] = 256'h580889065d045202eeff52fe72fda6fce4fcfcfd2d00ce024805870768083409;
    decBuf[10299] = 256'hed09950ac80a84090c07be0170fc9ef7bdf52bf5b9f603fa27fc18fe28ffc300;
    decBuf[10300] = 256'ha3016f02ad0275021001cbff50feb7fd89fdb3fd73fe21ff7d001e02f804b107;
    decBuf[10301] = 256'hdf0a030df40e4f0ffc0e870d330c070a9108b50605050c03300188fe0ffccff9;
    decBuf[10302] = 256'heff8bbf9e7fb1dff1b02d404e305ed04e1020501d1ff09000801a902a204f605;
    decBuf[10303] = 256'hb006e806b506cd05fa04ee03f902dd018300e2fec9fd64fc36fcb4fc5bfee3ff;
    decBuf[10304] = 256'h48013002b201f200feff9fff2f001a017901e90061ff68fd14fc52fc4bfebf01;
    decBuf[10305] = 256'h0a052d075808fd0706072606e20529051004df013eff7afddffb29fcf5fcaffd;
    decBuf[10306] = 256'he7fde8fc00fcd9fab3fa61fbfcfc85fe1efff0fec9fdd6fb72f932f752f696f6;
    decBuf[10307] = 256'hcbf7c4f928fcc3fda3fe6fffadff550088005a00dcff1cff6dfe4efe17ff6b00;
    decBuf[10308] = 256'haf01d901cd004dff82fdc9fc91fc2afdb5fde2fcd6fbe2fac2fac5fbd0fd7100;
    decBuf[10309] = 256'h8001d2018801340071008a01bb033105fd054c047301f3fda9fa60f98bfa4ffc;
    decBuf[10310] = 256'h8ffe9a006601a401fc0097ff52fed7fc72fb8afab7f9f7f849f8eaf7cdf7edf8;
    decBuf[10311] = 256'he0faccfd4b01a503c9052c06870634067f06c3068e0595033101f1fe11fe55fe;
    decBuf[10312] = 256'h8affa3007000cefef5fb3cf978f725f706f86afaf2fd3d011605ad0716098409;
    decBuf[10313] = 256'h9207190534027cff02fd0cfc2bfb6ffb32fb89fabcfaebfa15fbd5fb83fc21fd;
    decBuf[10314] = 256'h77fd2efe33ff6d00940107029f014300a1fe19fd1afcebfb6dfbadfafff9a0f9;
    decBuf[10315] = 256'ha2faaefc0f013004090796080f09c607d5051004d00130ff01fc03f94af63bf5;
    decBuf[10316] = 256'h8df503f767f94bfc03ff7d011803f8033c04ff03760277018f0065008b006800;
    decBuf[10317] = 256'hcaff54fe89fc55fbacfaabfbf0fc17fed7feb4fe55fe72fefafff30157044d05;
    decBuf[10318] = 256'h6d04090280fe27fcdefa42fb06fd46ffbc008801bc026503fe0389045f040503;
    decBuf[10319] = 256'h6401dbff42ff70ffefff1500dbfeb8fcacfa58f912fa0bfcf7feaf0174036b04;
    decBuf[10320] = 256'h4b05170655068d065a067205f7032c027b0082fe2efdfafbc1fbf4fb96fd8fff;
    decBuf[10321] = 256'h6b0124025c025d01d200a80068012d03de04860553056b04f0028b01460074ff;
    decBuf[10322] = 256'hb4fe7afdfffb9afa0ffae1fa87fcf1fe8c000202be010501ecff53ff25fff7ff;
    decBuf[10323] = 256'h9d0126038b0416059804f202f90095fef9fc19fc5dfc92fd3afed3fe48fecafd;
    decBuf[10324] = 256'hbdfc0ffc71fb1afb98fa51fa66fa65fb70fd11008b02ca044006840646062e05;
    decBuf[10325] = 256'h2f04ea026f01a4fff4fd6bfc6cfb3efb68fb8efb3cfc9bfcb8fc06fd7dfd15fe;
    decBuf[10326] = 256'h14ff0800a600c300d8fffdfd99fb59f979f8adf766f80ff90efa3cfa12faecf9;
    decBuf[10327] = 256'he0fabafca6ff5f022304750495033101a8fd4ffb2bf901f85bf852f9c8faa4fc;
    decBuf[10328] = 256'h4bff0f014f035a05ae066807bf06f404c802bd00e1fea3fedcfedbff66009000;
    decBuf[10329] = 256'h1d00b4ff13004f011f034a05c006040754057a02c2ff48fdadfbf8fb4cfdf3ff;
    decBuf[10330] = 256'hb701f7034204860451033902d40048001e00910040015f0196000eff15fdc1fb;
    decBuf[10331] = 256'h83fb2cfc5dfe6800cc0267047306d708160b220d660db50b6b08300434009dfd;
    decBuf[10332] = 256'h34fcc7fb63fb54fa14f89ef65af68ff788f974fc2dff3c0033017e01c201f602;
    decBuf[10333] = 256'h7f044a06fa078309820a540ad6092f0836064a03920018fed9fb63fa1ffa5dfa;
    decBuf[10334] = 256'he5fbe2fe9703f907d10a5f0c050a2c067a00b0fc3ef9def970fafefb58fea0ff;
    decBuf[10335] = 256'h9201560396053708460998092308bf057f0374012000ebfed2fd39fdaefc84fc;
    decBuf[10336] = 256'h11fc34fc53fce3fc37fe3500110246030d0342019bfe22fc86fa3cfa80fa42fa;
    decBuf[10337] = 256'hb9f822f6f4f2f5ef92ef56f1dff41af916fdb6001f026803cb03db0476065607;
    decBuf[10338] = 256'h9a075c076305ff021b0062fd9efb03fa22f966f9a4f94dfab2fbf6fcc6fe7600;
    decBuf[10339] = 256'hff016403920368035b022101fbffa1fe16fe43fdd0fc22fc84fb2efb48fb7cfc;
    decBuf[10340] = 256'ha0fed601d5045408bd092b0a39085604adff4cfb73f8e5f66df6dbf63ef74ef8;
    decBuf[10341] = 256'he9f9f4fbe0fe9901c704eb06dc08ec09870b670cab0cf20bf9090d078d034300;
    decBuf[10342] = 256'h1ffe2efc69fa72f992f8c6f70df745f7def723f99efa03fca4fd2dff2c00b700;
    decBuf[10343] = 256'h8d0080ffd2fef2fef4ffba016a03a203a302ebff6cfc12facaf866f8c1f813f9;
    decBuf[10344] = 256'hc8f8fcf7bef7b7f9b3fdd302a6078709f5085e0623024affbdfd35fe7effa800;
    decBuf[10345] = 256'h4e00fbff46009a014a039406ee08120b750b660a26088505c1032502db011f02;
    decBuf[10346] = 256'he101a901aa0008ff7ffde6fc15fd90fe5b0014016c00a1fef1fcb8fcb7fd1200;
    decBuf[10347] = 256'hf702e8044305a7033202de009701af02e004c1057d05cc0363017ffe54fdfafc;
    decBuf[10348] = 256'h4cfd2cfee8fd2ffd87fc54fc3cfd5fff0002c4031704a1023d0059fd67fb77fc;
    decBuf[10349] = 256'h12fe480147047105cc05d5048a04ce0403063b0608060a041e0165fea1fc98fd;
    decBuf[10350] = 256'h380067038a05b506a505af04ce031204470560062d064505cd02540014fe9efc;
    decBuf[10351] = 256'hd2fb10fcb8fc83fe2a0159045707100a890c800d350de10b310ae7069d03c3ff;
    decBuf[10352] = 256'h2dfdd3fa8af9eef9b2fbf2fdfdff51018602be02f102c30244023801b8ffedfd;
    decBuf[10353] = 256'h3dfc95fb2efc72fdedfeb8007201aa017701ec00c1009b007800daff9efecefc;
    decBuf[10354] = 256'h1efb25f9d1f793f7acf8ddfa7efdf7ff9201dd01990164004cff4dfe1efe49fe;
    decBuf[10355] = 256'hbcfe24ffc2ff8c00df0181030a05090637061005d00248fffdfbdaf921f75df5;
    decBuf[10356] = 256'h0af5c0f48cf5c0f69af919fd55015105fa09da0b6c0cdf0a85088605ce029fff;
    decBuf[10357] = 256'h7cfdc3fafff863f719f76df80bfcb3001505ee077b090309e006270418032102;
    decBuf[10358] = 256'h6c0228026e01e5ff1afee6fcaefcadfd4eff670000017400a2ffe2febffe9cff;
    decBuf[10359] = 256'hd900000273020a02ed0094fff3fddafcdbfbf3fa21fa61f96df88ff739f71ff7;
    decBuf[10360] = 256'h66f7fdf7d5f8d8f912fb39fc45fd3afe95ffda0055025403df03b503f5020102;
    decBuf[10361] = 256'h24015b000c00f4ffdfffa4ff27fff6fe22ffebff610192039d0579073208fa07;
    decBuf[10362] = 256'h9506dd03250141fdabfa51f809f7a5f600f79bf83cfbb5fd3e018804ac060f07;
    decBuf[10363] = 256'h4b056702aeff80fc37fb62fc26fe66007102c50303045b03c2027d01560049ff;
    decBuf[10364] = 256'h10fe94fc95fbaefa2ffa6ff9c1f8a1f8f8f84bfa49fcadfeed00f802d4041205;
    decBuf[10365] = 256'h6a049f02f7ffc9fccaf9d9f7e8f828fb5efe3802d7054107ae074b073b06a004;
    decBuf[10366] = 256'h9502a9fff0fcc2f99ef774f6cef669f875fad9fc74febffe7bfe46fd0efda7fd;
    decBuf[10367] = 256'h48ff2202da04ea05e0060006bc057e05b70550067e06ab05b8035401b9ffd9fe;
    decBuf[10368] = 256'h1dffcd00560255032703fd02d602ca03a50581073109f9082e07870458015afe;
    decBuf[10369] = 256'h68fc59fb06fbbcfa00fbb9fb42fd0dffbd00d60109027d01ab009eff36ff16ff;
    decBuf[10370] = 256'hf9feabfed5fdd2fc24fc83fcbffd8eff3f01570224023c016a00f7ff5f003d01;
    decBuf[10371] = 256'h93017901d300e5ff86ffdcffc700e401a402c702aa015100affe26fd27fc3ffb;
    decBuf[10372] = 256'h15fb88fb7dfcd8fd7aff030102028d025f03d3033b041c04df02670039fd15fb;
    decBuf[10373] = 256'h24f97ef9befbc9fda5ff5f00970064009200650171029402780138ff54fc9bf9;
    decBuf[10374] = 256'h8cf8def854fa30fc5cfed1ff2501d6025e04c305080786076007260657042b02;
    decBuf[10375] = 256'h2000bcfd21fc40fbfcfaadfca6fe82003b01030138ff88fdfffb66fb4efc74fd;
    decBuf[10376] = 256'hcefe59ff2fff22fe2efd51fc6dfcf0fcc6fd56fea4febcfe7bfeb6fe57ffeeff;
    decBuf[10377] = 256'h50001a0027ffedfd6efd95fdcffe9e00d301eb0252026b01efff8afea3fd24fd;
    decBuf[10378] = 256'h64fcb6fb18fbfbfae6fbc1fdbd01b9055809a30ceb0d880d780cdd0ad2085e05;
    decBuf[10379] = 256'h230126fd7ef81cf467f2ebf254f478f669f8c4f816f9cbf897f9c3fb64fe9201;
    decBuf[10380] = 256'hb6031904bf03c8027d02c1027204fb0560078e07bb06af052f0464022f01a6ff;
    decBuf[10381] = 256'hdbfd2bfc13fb14fa2cf9adf83af817f876f8ecf983fcfcfee1010b0366031303;
    decBuf[10382] = 256'hc90285023e0376034303fe0187ffc2fd27fc72fc3efd72fe1bffe8fe5dfedefd;
    decBuf[10383] = 256'h05fe6dfe0bff62ff7cff93ff2b002a0164023603c302fe0057feddfb42faf7f9;
    decBuf[10384] = 256'h3bfa70fb18fce5fbb7fb35fc42fd4dff830282053a08ff09510a71091d086d06;
    decBuf[10385] = 256'h73049702de0136010301d4005600e3ffeffed2fd12fdeffc4efd51fe8bffb200;
    decBuf[10386] = 256'h0b02f302710398037503980295015b00e0fe7bfd36fc64fba4fa3bfad9fadcfb;
    decBuf[10387] = 256'he7fd8800010341054c07a0085a0992095f097708fc069705f5034d031a03ec02;
    decBuf[10388] = 256'hc10202023c0010fedafab7f88cf7e7f7ddf8e9fad5fd8d005202ed03cd041105;
    decBuf[10389] = 256'hd3040c057304a104770450042e04cf033f03bc021602d5019a0141018e0089ff;
    decBuf[10390] = 256'h09fe3efc8efa75f976f848f81ef8def85dfa8efc2fffa9018d0445070a09010a;
    decBuf[10391] = 256'hb6097209c207c9056503c901e9001d0064ff4bfee6fc8bfa4cf801f855f9fcfb;
    decBuf[10392] = 256'he0ff7602df034d042203c8027502eb03c7058006d8050d046601ecfeadfca1fa;
    decBuf[10393] = 256'h3df8fef5c7f2a4f040f005f232f652fbc4fee5019a031f049704e0050a07cf08;
    decBuf[10394] = 256'h7c080707930357ff7efce8f970f902f92dfaf1fbe8fc5efe2aff5e009600c900;
    decBuf[10395] = 256'h3e0017ff0bfe8bfc8cfba4fa26fa33fbf8fc9fffce02f1041c06c10526044603;
    decBuf[10396] = 256'h02033f0358048b040004dc01a6fea8fbeff8e0f732f812f9def997fa40fbd9fb;
    decBuf[10397] = 256'h64fcdffd10001b02f703b004e9045004c4034603b90322044104b203c7026b01;
    decBuf[10398] = 256'h8300590019010d02ab025502350142ff66fd32fc6afc03fd47fec2ffc100f000;
    decBuf[10399] = 256'hc600060012ff74fe57fed9feafff3f008d004600daffc6ff4300370171029803;
    decBuf[10400] = 256'h5804350497034103f2027b020f02e9001affeefc78fbacfa65fb7efc7dfd65fe;
    decBuf[10401] = 256'h8ffe69fe46fee4fe93004302cc03ff037403a501f4ffdcfe0ffff7ff7201d702;
    decBuf[10402] = 256'h1b0446041f04b7031803c202a80290027b02f1012d014200a3ff87ff6dff84ff;
    decBuf[10403] = 256'h43ff44fec5fc60fbd5fafffa0bfc45fd18fef1fd43fda5fcc2fce1fdd4ff3802;
    decBuf[10404] = 256'h1c050e071d086f088f07c3061305fa0395020a023801c4005c00beff67ffeaff;
    decBuf[10405] = 256'hc000fc01cf025c022201fefef3fc9ffb61fb7afcdffdc7fef1fe7efe15fef5fd;
    decBuf[10406] = 256'hf8febd00e9028a054e07a10756070206d603cb01efffbafef2fe25ffb0ff86ff;
    decBuf[10407] = 256'h13ff65fe84fe4effa10043025b038e030303880123003bffbdfee3fec0fe61fe;
    decBuf[10408] = 256'h0bfebdfd04fef2fecfffd2003b015a010401b6006e0059006c00a20034013302;
    decBuf[10409] = 256'h6d0394040705e404c8036e022a010001730121028002630244019effa5fdc9fb;
    decBuf[10410] = 256'h94faecf985fac9fb44fd0fffc000d801d702bf033d04170469038b0216011700;
    decBuf[10411] = 256'h8bff0dff33ff11fff1fe0eff28ff9fff0b00f7ff0fff74fdebfb86fafbf979fa;
    decBuf[10412] = 256'h39fbe7fb07fc24fc3efce4fcfdfd0afffeff9c00b9009f00b6002201ac01e101;
    decBuf[10413] = 256'hf201c501680113018400acff70fe49fd3cfcd4fb33fc35fd29fe88fe6cfeb5fd;
    decBuf[10414] = 256'h6dfd05fe2bff4f015a0326046404bb03bc0231025b023502cc012e01f2ffcbfe;
    decBuf[10415] = 256'h0bfe5dfd3dfd5afdddfdb2feefff6a01cf0213043e046404fb03dc03bf03a503;
    decBuf[10416] = 256'h5e039b02e4010e0145008eff89fe09fd3efb8ef9e6f8b3f83ef910fa84fa32fb;
    decBuf[10417] = 256'h8efc8cfe00024b0549087409190922084207fe063c079306c804a601f1fcd0f9;
    decBuf[10418] = 256'h1bf89ff808fa07fd6afd10fd19fca3fa5ffa19fb12fd66fe1fff77fe78fd90fc;
    decBuf[10419] = 256'hbafc7afd6efecdfe76fe57fd97fcbafcd7fd1600fb02ec0466075c08d209160a;
    decBuf[10420] = 256'hd8094f081e065302b3fe69fb6af879f669f572f4bdf489f539f7a3f92bfd7600;
    decBuf[10421] = 256'h7503660576066c07b70773073e062605f502e90095ffe5fd3dfda4fc19fc9afb;
    decBuf[10422] = 256'h0dfcbcfc57fee0ff4501d001520192009effc0fe30feaefda9fce3fab7f8acf6;
    decBuf[10423] = 256'h68f69df706faebfca3ff1d0213035e032a04e304fc052f0647052303edffeffc;
    decBuf[10424] = 256'h36fa27f930f850f794f7d1f7eaf81bfbe7fe8f03b106ad0a310bb90a9508dd05;
    decBuf[10425] = 256'hae02b0ffbefdfafb5ffa7ef93af978f991faf6fbf4fdd0ff8001990298032304;
    decBuf[10426] = 256'h4d0473045104730370023701100003ffe0fe3fff080028013402e30202031f03;
    decBuf[10427] = 256'h3903df03a2045905a0050905e2036b01f1fe56fde0fb9cfb5efb26fbbffba7fc;
    decBuf[10428] = 256'h22fe5300f4026d05ad07f807b407fb06e2051704eb014bff1cfc1ef92cf71df6;
    decBuf[10429] = 256'h6ff6e5f739f96dfaf6fb5bfda0fe6f001f02a803410470049d0390029c013d01;
    decBuf[10430] = 256'h94011602bd022903ee0229020a01b0ff25fffbfe6eff1d00fdfffafeeffc4efa;
    decBuf[10431] = 256'hd5f783f7f8f8e4fb9dfe16010d02c201f6003401bd02880438060006cf032e01;
    decBuf[10432] = 256'h00fedcfb40fc4ffd46febcff78ff43febafc21fc50fc77fd1dff16016a029f03;
    decBuf[10433] = 256'h47047a044c042104ae03ba021f0126ffc2fc27fb46fa02fa40fa59fb58fce3fc;
    decBuf[10434] = 256'h0dfd33fde2fd3eff3c01a0033b05b106e505b00427035c0127007fff80fe3bfd;
    decBuf[10435] = 256'hc0fbc1faf0fac2fb02fe42004d02a1036303da010f005ffe46fd47fc19fceffb;
    decBuf[10436] = 256'h7cfbcdfaaefa04fbeffb8afd13ff7800600136015c013901d801da02ce036d04;
    decBuf[10437] = 256'h890407046003c902dd027e034004f704df04c603d3016fff30fd24fb58fa1bfa;
    decBuf[10438] = 256'he2f97bfa07fb85fbabfb5afc37fde6fe1201b3032c066c084c098008d006d704;
    decBuf[10439] = 256'hfb02c6011e01eb00600039ff93fd9afb46fa8cf9c4f9c3faabfbd2fc92fd86fe;
    decBuf[10440] = 256'ha3ff4901d2026b033c0316026f0076feaafde8fd90fe29fffbfed4fd2efca5fa;
    decBuf[10441] = 256'h72fafdfa78fca9feb5000902c202fa022d035b03860312031e02c20021ff08fe;
    decBuf[10442] = 256'h6ffdfbfd76ffdb007c022403f1026602eb0086ff42fe6ffdfcfc93fcf5fb9ffb;
    decBuf[10443] = 256'h85fbfbfb15fdbbfeb40008023d03e5031804ea03bf0333049b04fa0417056004;
    decBuf[10444] = 256'h5b039501e5ff5cfec3fd95fdbffd32fe55fef6fdd9fdf3fd6afe58ff75003501;
    decBuf[10445] = 256'h5701b9002a000f0086009f014503ce046705dc04b5030f02860087fffcfed2fe;
    decBuf[10446] = 256'hf8fe1bff3bffe5fe96fe20fedffd7dfd47fdf6fc8efcfbfb99fb64fbf6fb1cfd;
    decBuf[10447] = 256'h40ff4b0127035c0494046104d6030004da03fc035e03e901b8ffacfdd0fb17fb;
    decBuf[10448] = 256'h4ffbb4fc56fe6eff07003600b7ffdeff00009f002e01480101013f0088ffe1fe;
    decBuf[10449] = 256'hccfe55ffd2ff65005100d4ffe0fea6fdd4fcadfcd0fc6efdfefd4cfe64fea5fe;
    decBuf[10450] = 256'ha4ffaf015004c9060909e909a5097a07d904aa0187ffcefc55fabaf8d9f70df7;
    decBuf[10451] = 256'h4bf7f4f7bff96ffbf8fcc3feee006402400475058e065b06cf05a9049c03a802;
    decBuf[10452] = 256'h0a027a01c3001d00b1ffc4ff1e008f00d900b100fbff44fffdfe94ffbb00de02;
    decBuf[10453] = 256'h54049804df035602f100c3009501550278029b01ebff44fd35fc87fc28ffa101;
    decBuf[10454] = 256'h8504b0050a0614053304ef032d0465043204a703d502c8015f017f014802ff02;
    decBuf[10455] = 256'h460305032e02f100caff0bffe8fe47ffd6ff8d00d40094000a0046fff7fe3eff;
    decBuf[10456] = 256'h2c00880170029a02270233011600f0ff590036013902a10242027901f700af00;
    decBuf[10457] = 256'h9a00ad00540081ff44fe1efdaafccdfcabfde7fe6200c701af022d035403eb02;
    decBuf[10458] = 256'hce0128002ffe53fc1efb76fa43facefa4dfbc0fbb4fc10fe54ff7b008801f001;
    decBuf[10459] = 256'h920102014b00a5ff0dff5dfe87fdbefc3bfc82fc45fd64fe71ff650085006800;
    decBuf[10460] = 256'h4e00360020000d0090ff9cfe91fc86faaaf875f7adf712f910fbfcfdb5002e03;
    decBuf[10461] = 256'hc9041405480413031a01c6ff16fefdfc98fbb0fa32fabff96dfa8afb30fdb9fe;
    decBuf[10462] = 256'hb8ff43006d00e000d4017003f804f7056c05f103c001b5ffd9fd9bfdd3fdd2fe;
    decBuf[10463] = 256'h5dff33ff0dff5ffe00fe1cfed3fea9ff7200f5000d0122013601d701c502a203;
    decBuf[10464] = 256'hf803de03d9029f01cc0059007c00db006b01ed0105021b027d021e03e0039704;
    decBuf[10465] = 256'h0e05f8042104ab02e000abff03ffd0fe5bff82004201f0011002660251036e04;
    decBuf[10466] = 256'h2d059605b9040903e7ffc3fdd2fb77fb6efcb9fcfdfc3afd73fd0cfeadff1602;
    decBuf[10467] = 256'h56046106a506ec05d304d403a603d003f70319047b03ec029d02e4027c030504;
    decBuf[10468] = 256'hd003dc021601ebfedffc8bfbd2fa2afa5dfaa1fb71fd9dff3d02020454049f04;
    decBuf[10469] = 256'hd30395035d0390036203e3028a014500c7ff3a0074019b025b0366028c00b0fe;
    decBuf[10470] = 256'h84fc3afc7efc37fd4ffe1cfeeefd70fd96fdd0fe4b001602cf0227025c0030fe;
    decBuf[10471] = 256'h25fc59fb97fb20fd85fec9ff9c000f013201910120020c03e90306041b037f01;
    decBuf[10472] = 256'h86ffaafdf1fcb9fc86fcb4fc8afccafba7fbc7fbcafc49fe48ffd4ff55fffcfd;
    decBuf[10473] = 256'h14fdeafcaafd29ff8e007601a0012d01c5002301ed010c031904810422042003;
    decBuf[10474] = 256'ha001d5ff25fe9cfc37fb4ffa25fa4bfafafad7fba0fcc0fdccfe06008101e602;
    decBuf[10475] = 256'hce034d048d03530283004fffc6fd61fc79fb52fa92f92af9c8f93dfb6efd7aff;
    decBuf[10476] = 256'hce0087014f011c014a011d02dd028b032c0329021e0013feaffbb8fa6efab2fa;
    decBuf[10477] = 256'h6bfb13fc78fd60fe33ffa6ff0e00efff99ff7eff67ffd3ff8300fa0066012b01;
    decBuf[10478] = 256'hae00dbff12ff5bfee4fda3fd90fd5afd4afd59fdb6fd6cfe57ff740080012f02;
    decBuf[10479] = 256'hcd02ea02380350033a03270386026d01130072fec9fd96fd7efef9ff5e01a302;
    decBuf[10480] = 256'hcd02f4024502e6015701a000f9ffe0fed4fd25fd06fd95fde9fe8a0013021203;
    decBuf[10481] = 256'he402ba024702980179015c01aa01f2015e0271023c02ca010a011f0042ffb2fe;
    decBuf[10482] = 256'h98feb0fef0fe2bff85ff37000d01490270033004530436039001070008ff37ff;
    decBuf[10483] = 256'h09006301a7022603ff0251027401aa002800b1ff70ffc0feeafd5afd0cfd53fd;
    decBuf[10484] = 256'h97fe3900c201c1024c0322036202f901d901bd01d7019001230173009dff0dff;
    decBuf[10485] = 256'hf3fedbfe1cffcdffa300a501df02b203d8037003140216003afe89fc01fb02fa;
    decBuf[10486] = 256'h76f94cf973f967fac3fbc1fd9dff4d01660233024b01240017ff69fe0afe60fe;
    decBuf[10487] = 256'he3feb9ff82006d010b0228020e029701a9008dffe6fdedfb11fa61f848f715f7;
    decBuf[10488] = 256'hfdf7cdf9f8fb04fe58ff1100d9ff40ffb5fe8bfe64fe41fe22fe92fd44fdfcfc;
    decBuf[10489] = 256'h12fdc3fdf7fec700770200046505930515056f03760112ffd2fc5cfb08fad3f8;
    decBuf[10490] = 256'h2bf8f8f783f8aaf99dfb01fe4100b6018202c0028802ef016401e5007200c4ff;
    decBuf[10491] = 256'h26ff09ffc0ffc500ff01d2024503dc027d027b01cc00b0ffa3fe69fd42fc82fb;
    decBuf[10492] = 256'h5ffb3dfc40fd34fe93fe76fe27fe3ffe2dffc800c1029d0457051e05b9037502;
    decBuf[10493] = 256'hfa00fbff59fed0fc6bfb84faaefaedfc7600b1048a071809900948088f05cb03;
    decBuf[10494] = 256'h8b0180ffa4fdf3fb6afa6bf9e0f8b3f9a6fb0afea5ff1b01e701a90171010a02;
    decBuf[10495] = 256'h9502bc03c904310512050f04d502ae018801ab0149026502e301de005efff9fd;
    decBuf[10496] = 256'h6efd98fd58fe4cffeaffcdff4bffa4fe38fe9afea7ff4d01d6026f034003c202;
    decBuf[10497] = 256'hb5014d01ee000a01590141010001ed002201d5010a03dc034f045b03810195fe;
    decBuf[10498] = 256'hdcfb18fac6f910fadcfa96fbaefcadfdf2fe6d003802e8039104f80310039501;
    decBuf[10499] = 256'h300048ffc9fea3fec6fea6fec3fe11ff88ff4b000201d7012e027c026402cd01;
    decBuf[10500] = 256'h1c01170023ff06fe93fde5fc86fc30fcadfb95fb01fc01fd80feb100bc029804;
    decBuf[10501] = 256'hcd0576064306b705e8033802ceffeafcf9fae9f93bfa86fa52fb87fc2ffd2efe;
    decBuf[10502] = 256'h16ff3d0096017e02fd028a025001d5ff70fe2bfdadfcd3fc3cfddafda3fec2ff;
    decBuf[10503] = 256'h1c0160023303a6033d032102c70026ff0dfedafd66fe38ff4500f30013018300;
    decBuf[10504] = 256'h64ffa4fe3bfedcfdf9fdabfd04fd42fcf3fb6afc83fd76ff52018702a003d303;
    decBuf[10505] = 256'h0104d70364037002140116ff3afd05fc5cfb8ffbd4fc4ffeb4ff9c006f01e201;
    decBuf[10506] = 256'h0502e501c80146019f000800cdffdfff920097014502a402c1023e02c8013001;
    decBuf[10507] = 256'ha7002a0098ffc0febdfd83fc5cfb9cfa79fa99fa62fb82fc28feb1ff7c01b002;
    decBuf[10508] = 256'h39043805c305ee05c70519057b04b103fb0225022201e8ff16ff09fea0fd81fd;
    decBuf[10509] = 256'hd7fd25fe6dfe82fe96feeffea2ff78007a012902090279018e0072ffb2fe49fe;
    decBuf[10510] = 256'h2afe46fec9fe10ff7cff2d00d3006b01f4012a023a020e02e5010a0257028902;
    decBuf[10511] = 256'h8002140237015a0091ff42ff5aff70ff83ff71ff41ff32ff75ffe2ff49008c00;
    decBuf[10512] = 256'h4f00ecff8fff6aff75ffa7ff7afffefef2fde5fc37fc17fc1afd54fecfffce00;
    decBuf[10513] = 256'hb6018802950389046705bd056e050a043f0213009efed2fd18fde0fcadfc7ffc;
    decBuf[10514] = 256'ha9fc1cfdcbfd29fe46fef8fd22fd92fc44fc5cfc4afd66fec0ff04017f02e403;
    decBuf[10515] = 256'h29055006c306a006c30586040b030c02c80049003dff49fe2cfd1ffce5fa13fa;
    decBuf[10516] = 256'ha0f97df95df9b3f99ffa3afca3fee3008403fd05f406a906dd05a8040004cd03;
    decBuf[10517] = 256'h9f03c90356036102060107ffb3fd7ffc47fc14fc42fcc0fce7fc4ffdaefd77fe;
    decBuf[10518] = 256'h2eff0400cd005001f6016202ec026903db032404fc0377036b02110170ff57fe;
    decBuf[10519] = 256'h58fd87fd59fe66ff5a0037018e017401fd000f00f2fee6fd37fd99fceffcdbfd;
    decBuf[10520] = 256'h36ffd8006102c603ae042c059f057c051d058e04d703010338028101db00edff;
    decBuf[10521] = 256'h0fffd3fdacfc39fc16fc75fccbfce5fc9efc32fc6dfc55fdf0feea00c602fa03;
    decBuf[10522] = 256'ha3047004410417048a04ad048e04c403a5024c01070034ff74fe0cfeadfd1dfd;
    decBuf[10523] = 256'hcffcb7fc23fd22fe5cff2f00ef001201b300b0ff76fe4ffddcfcb9fc97fd0cff;
    decBuf[10524] = 256'hd7000c022503f2020a0237012b000800e8ffcbff7dff06ff18fe7afd24fd3efd;
    decBuf[10525] = 256'he4fda7fe2aff71ff5bff48ff59ffabff2f00ad00dd009400000050ff09ff75ff;
    decBuf[10526] = 256'h7400ae01d502fb0207026c0002fec3fb4dfa81f943f9ebf950fbf2fc7bfeac00;
    decBuf[10527] = 256'hb70293044c058405eb044a03c1015c00d1ff53ff79ff56ffb8feeffd04fd26fc;
    decBuf[10528] = 256'h96fbb1fb27fceafca1fd47feb3fe64ff3a003c013002cf02eb02690293019000;
    decBuf[10529] = 256'he2ff83ff66ffb5ffccffe2ffceff99ffa9ffd5ff4e0000017701e301d0017601;
    decBuf[10530] = 256'he4005b000100d0ffa4ffb2ffa5ff84ff52ff13fffafe1fff6bffedff6a00dc00;
    decBuf[10531] = 256'h43018601db015402e6026f03a5033303560239017a0011003100c0000f01f700;
    decBuf[10532] = 256'h340049ffabfe55fea3fe49ff0c008f00a60091007d006b007c00a800b500da00;
    decBuf[10533] = 256'h11016b01f0016d02ff0213030103b00249020602b1017a010c014c0095ff90fe;
    decBuf[10534] = 256'he2fd43fd27fd0dfd24fd65fdc7fdb0fe8dffc9009c015c027f022002ca01af01;
    decBuf[10535] = 256'h9801ad01c101d30182011a016c00c6ff2fffcdfebbfecbfef7fe3aff5fff6aff;
    decBuf[10536] = 256'h4cff30ff17ff01ffd1fe73fefbfd68fd2efd3ffdf2fdf7fe31000401c4012c02;
    decBuf[10537] = 256'h8b02a802c202da026e02bd01880062ff55fe61fd02fde5fcfffca6fd68fe53ff;
    decBuf[10538] = 256'hf1ff81006700c1fffefe47fed1fd90fda3fdb5fda5fdb4fdf7fdacfe00004501;
    decBuf[10539] = 256'h6c02df027602d8010f0158001100d0ff6effcdfe35feacfd9afdcbfd32fe90fe;
    decBuf[10540] = 256'h84fe4dfef3fdb6fd95fdb3fdf3fd5efee3fe84ff1b00a400fe002f015b018301;
    decBuf[10541] = 256'hd80125026b023d02c101b5000fff86fdedfc62fc8cfcb3fc61fdfffdc8fee8ff;
    decBuf[10542] = 256'hf400a30141022402d60130014200a4ff14ffc5fe7efe69fe7cfeb2fee3fe0fff;
    decBuf[10543] = 256'h1cff10ff47ffa1ff3f000101b8012f0245023102d80145019500eeff2cffa9fe;
    decBuf[10544] = 256'h62fecefe7fff84007801d701ba0138016200d2ff84ffcbff8e00100187017101;
    decBuf[10545] = 256'h0f016e000200a0ff6aff3affb5fe14fea8fd6dfd0efe27ff3400e200c200c0ff;
    decBuf[10546] = 256'h40fe41fd6ffd96fed60016038b0457051a0571043e04b30389037c02430173ff;
    decBuf[10547] = 256'hc3fd3afc07fc92fc0dfe72ffb7008a016301b5001700c0ffa6ffbeffd4ffe7ff;
    decBuf[10548] = 256'hb2ff40fff6fe04ff71ff4e006b017702e002c00230027a010301c200d6000b01;
    decBuf[10549] = 256'hda005600b5ff49ff35ff8eff2100aa00e000f000c40081004400f7ff9dff30ff;
    decBuf[10550] = 256'hc9fe86fe7afeddfe8bff3100c8005201870198014e01bb00e3ff1aff2efed0fd;
    decBuf[10551] = 256'h26fea8fe1fff8bff78ff42ff52ff9cff65002e01e501fd01bc015a01dc00ed00;
    decBuf[10552] = 256'hfb00ee008100c1ffd6fe38fe55fed7feadff3d005700b1ffeefe03fe65fd0ffd;
    decBuf[10553] = 256'hf4fc3cfd7dfddffda3fe8effab00b801ac020b0327030d039702a9018c0033ff;
    decBuf[10554] = 256'heefd1bfda8fccbfc2afdbafd3cfe42ff3600d1015a035904e4041104b8025d00;
    decBuf[10555] = 256'h1dfea8fcdcfb9efbd6fb09fc94fc12fd1ffe59ff2801d902f103240499037202;
    decBuf[10556] = 256'h6601710094ff77ff29ff11ffd0fe47fe11fe22fea6fe8fffab001e01fc001e00;
    decBuf[10557] = 256'ha8fea9fd7bfdf9fd53ff97006a01dd01ba019b01f1013f02b602cc02f401b800;
    decBuf[10558] = 256'he8feb3fd9bfccefc59fd2cfeebfe54ff34ff8bff0d0013014c021f03df03bc03;
    decBuf[10559] = 256'hdf0215022a01cb00af00c900e1002101e7008d001b0079ffe2fe58feb8fd20fd;
    decBuf[10560] = 256'h70fcf9fbb8fb1afcdffc32fed4ff5d015c024303c2033504580477049404ae04;
    decBuf[10561] = 256'h9704d403b5020e0115ffc1fd8dfc54fc87fc6ffd42feb5fed8fef8fea1febbfe;
    decBuf[10562] = 256'hd3fee9fefcfe0efffefeeffe17ff85ff4400fb00d1019a02e9020003eb02b002;
    decBuf[10563] = 256'h9e02ae029f0242028c013800f4fecdfd5afd37fd56fde6fd35fe1dfedcfdc8fd;
    decBuf[10564] = 256'hfefd70fe4dffebff7b0061001900d9ff9eff8cffbdffe9ffdbff9fff7eff88ff;
    decBuf[10565] = 256'hdaff7f00250191017e014801d6006f00470053005e007c006100480031000f00;
    decBuf[10566] = 256'h09000e00280052008400a700b9007c00000083ff11ffe5fef2fe2fff3afff4fe;
    decBuf[10567] = 256'h7dfe0bfe1afeadfe85ff8800ab008b0088ffdafe7bfe98fe4fff2400b4000301;
    decBuf[10568] = 256'heb00d50010016901db012502fd017701b300fcff26ff5dfedafd34fdc8fcb4fc;
    decBuf[10569] = 256'h0efdc0fd96fe5fffe2ffb8008101a002ad035b04ba046404ad033603ca02de02;
    decBuf[10570] = 256'ha8021602f000ccfec1fc6dfb38fa70fa09fbf1fb18fdd8fd86fe64ff2d001801;
    decBuf[10571] = 256'hb6010c02f201ab013f012b01190109011801f000b3005000bdff0cff66fefafd;
    decBuf[10572] = 256'h35fef9fee5ff0101740197013801a9005a004200020078ff6cfe13fdcefba4fb;
    decBuf[10573] = 256'h64fc6ffe100189032405050649060b06d30506067b055404ae02440060fd6ffb;
    decBuf[10574] = 256'haaf9b3f869f8adf8eaf803fa02fba3fc9cfe78002902b203b1043c056605a604;
    decBuf[10575] = 256'h2603c1017d0056ff96fe73fe53fe37fe1dfe64fed0fe81ff2700be00d2009c00;
    decBuf[10576] = 256'h2a00e1ffb9ffddfffefff4ffd9ffafffa8ffe6ff610002019a01ad0178012601;
    decBuf[10577] = 256'hbf00b200d600230155012801cd006000160023007800af00a5001c001dff29fe;
    decBuf[10578] = 256'h4cfdf5fc44fdeafd03ffc3ff2c004b00f5ff72ff2bff16ff29ff83ffd4ffe3ff;
    decBuf[10579] = 256'hd5ffb1ff7aff84ffb1ff0c00490054000e00ceffc6ff36002a0164028b03fe03;
    decBuf[10580] = 256'hdb033d037402bd014601300144010e015c0086ffbdfe6efeb5fe22ffabff99ff;
    decBuf[10581] = 256'h27ff68fee5fd9efddffd41fe9afe8afe23fee0fdecfd91fef5ffc001f5029d03;
    decBuf[10582] = 256'h6a03df02b8015f0077ffa4fe31fec9fd6afd13fdf9fc41fdadfd85fec1ffe800;
    decBuf[10583] = 256'ha8011002f1016101de006700fbffe8ffd6ffa5ff5bfffefe0aff83ff7700f601;
    decBuf[10584] = 256'h5b03e60310049d03a902cc01030180003900cdff1cff76feb3fd30fde9fcfffc;
    decBuf[10585] = 256'h3afd93fde4fd69fec2fe34ff7effc1ffcdffd8ffbaff7aff0fffc5fe82fe8efe;
    decBuf[10586] = 256'hf1fe84ff3500ac00c1005f00e2ff50ff3cff4eff9fffe9ffdcff9fff52ff48ff;
    decBuf[10587] = 256'hbfffb300a701c302360359033a031d0337034f033903b002c701ab00ebff3dff;
    decBuf[10588] = 256'h1dff3aff20ffd8fe41fe42fd4efceffbd2fb55fcfbfce9fdc6fe56ffd9ff4f00;
    decBuf[10589] = 256'hbb0045019e0110025a0267022a029b01c400c1ffcdfeeffd99fd4bfd62fd78fd;
    decBuf[10590] = 256'h01fe7ffe31ffd8ff6f00aa00bc008b0041004f00a3001c01af01110223023302;
    decBuf[10591] = 256'h42026a02bf020c032a030e03c4026a021502de01840117013a001dffc4fddcfc;
    decBuf[10592] = 256'hb5fb42fb1ffbbdfbc0fcfafdccfe8cfff5ffd5ffb9ff9effe6fffbff5d006f00;
    decBuf[10593] = 256'h5f0033000b002f00660098008f0013004fff63fec5fda9fd2bfed1fe69ffa4ff;
    decBuf[10594] = 256'h92ff61ff52ffcbff9e00da010103c1032a0449042c04de0367032603c4024702;
    decBuf[10595] = 256'hd50133017100baff13ffa7fe6cfe5bfe4afe1efef6fda1fd80fd9efd02fe96fe;
    decBuf[10596] = 256'h1fff9cffcdffa1ff5eff21ff00ffe2feebfed2fe9efe45febffd42fdf1fc3bfd;
    decBuf[10597] = 256'h03fe3fff66007301dc01fb01a50157013f0129013d012b01fa00b0006e007a00;
    decBuf[10598] = 256'hdd00a501a8025603b5039903e2023b02cf016d015b012b01e1006800d6ff4dff;
    decBuf[10599] = 256'h17ff27ff36ff44ff07ff8efefcfd72fd3dfd4dfd97fdf4fd49fe96feb4fef4fe;
    decBuf[10600] = 256'h3eff98ff050032003f00eaff71fffffe98fe8bfe97fea2fe98fe7dfe43fe3bfe;
    decBuf[10601] = 256'h50feaefe76ff40002b0147020703b6031404a404f3046905aa059705f604dd03;
    decBuf[10602] = 256'h83023f01180058ffeffe90fe3afe4ffdb1fc21fc3bfc11fd4dfec8ffc7005201;
    decBuf[10603] = 256'h2801b500920033001700fdffb5ff1eff6dfe98fdcefc4cfc04fc1afc55fcf6fc;
    decBuf[10604] = 256'h8dfd17fe70fea1feeafe63ff1600eb00b5016b02b3029d028902780288029702;
    decBuf[10605] = 256'h6e0201025f019c001a0032009e0076013f028d02a50264020202a90157010e01;
    decBuf[10606] = 256'hcb004500c8ff77ff4bff8efffbff7f00b5008400e2ffc9febcfdc8fc2afcd4fb;
    decBuf[10607] = 256'heefb06fcf0fbb5fb80fb6ffbb9fb82fcbefd39ff9e00860159027f02a202c102;
    decBuf[10608] = 256'hde02c4027d02e5010e01440059fffafe17ffceffa4006d01f001a8013c016400;
    decBuf[10609] = 256'hd5ffefff65007f013e02ed02cd027702f401ad01c301fe01330202027e019500;
    decBuf[10610] = 256'hb8ff28ffdafec2fe81fe46fe82fd97fcb9fbf0faa2fa18fbdbfbfafc07fe70fe;
    decBuf[10611] = 256'h8ffe39feb6fd9ffddffd69fe2dffe4ff8b00cb002e01ce0166023e03cd031c04;
    decBuf[10612] = 256'hd5033d036502d60153013b0151011601e0008f00450053008f00f20035014101;
    decBuf[10613] = 256'h0a01ec00f5002f018201e5010d021902cc014a01a900e6fffbfe1efe55fdd2fc;
    decBuf[10614] = 256'h5bfc46fc32fcfcfbecfbddfbebfb40fcb9fc4bfdfcfda2fe0eff97ff1400a700;
    decBuf[10615] = 256'h3001ad01fe01d2017501ef009600a6000d01a0012a025f0270022602e301d701;
    decBuf[10616] = 256'hf8012a026a0283024e02f50188010301cd00bd00e9006201d3013b0248020b02;
    decBuf[10617] = 256'h9201e00039004bffadfeabfdb6fc9afbdafa2cfa4bfaa1fac1fbcdfc4dfe4cff;
    decBuf[10618] = 256'h3400b200d900410122010501eb0074000800a6ff4cff1cffd2feaafe85fe90fe;
    decBuf[10619] = 256'h9afedafe25ff7fff0400a5006701870247033b045a043e04bb03440303033e03;
    decBuf[10620] = 256'h9803e9031504d20335034702690167002dff5afe9afd32fdd3fc7dfc62fc7afc;
    decBuf[10621] = 256'h39fc26fcf0fb00fc4afcc2fc75fd1bfeb3fe15ff6effc0ff09004c0058003700;
    decBuf[10622] = 256'hddff88ff51ff83fffaff8c00ee002401d3003100c4ff62ff74ffc5ff2d008a00;
    decBuf[10623] = 256'haf00d000ee001b017601fb017902ea02340341033503e8028e02520231024f02;
    decBuf[10624] = 256'h6a0283025d02f60136014b002fff22fe2efd51fc87fb05fb8efa4dfa61fa02fb;
    decBuf[10625] = 256'heffb0cfd19fe0dffabff010084002a019601f801c30110010b008bfe8cfda4fc;
    decBuf[10626] = 256'h7afcedfc9cfdf7fe3c00630170026403020458043e04c7033003a6024d023d02;
    decBuf[10627] = 256'h6902ac02d002c5026b02fe0179012001ae0082002400d0ff57ffc4fe62fee5fd;
    decBuf[10628] = 256'h94fd4afd07fde3fceefc0cfd4cfda6fdfbfd48fe66fe5dfe55fe3efe45fe8afe;
    decBuf[10629] = 256'h01ff93ff4400ba00d0009500180045ffb5fe67feaefe45ff4400f30091012102;
    decBuf[10630] = 256'h3b0252029302a702b902a9027c0254021802f701c50172010f01b2005d003c00;
    decBuf[10631] = 256'h5a009a00d400db009d00210081ffe9fe60fe06fed6fda9fdb7fddbfd12fe58fe;
    decBuf[10632] = 256'haafef7fe01ffe6fe9cfe56fe28fe51fec2fe75ff1b0087009b001d004aff81fe;
    decBuf[10633] = 256'hcafdb2fd1efecffe75ffe1ff1c000a00faff090067000401c7014902c0020103;
    decBuf[10634] = 256'h3c039503070451044304d6031703f701eb00f6ff98ff08ffb9fe72fe06fea4fd;
    decBuf[10635] = 256'h6efd3efd87fde5fd6afe0bffa3ff2c00cd000e012101c80015003fff76febffd;
    decBuf[10636] = 256'ha8fd92fdcdfd02fe13fe21fe14fe20fe41fe87fed9fe26ff80ffd5ff7a002001;
    decBuf[10637] = 256'h0e02ec024203900379030c03aa02750244021802d5018001070195001000b7ff;
    decBuf[10638] = 256'h66ff57ff4aff6effbbff3d00ba002c013b0113018d00ecff55ff1aff08ff18ff;
    decBuf[10639] = 256'h27ff4fff74ffabffc9fff6ffeeffc9ff61ffbffe28fe9efdfefc91fc2ffcfafb;
    decBuf[10640] = 256'he9fb16fc73fc29fd49fe55ff8f00b601c30271039103ad035f031803ac027102;
    decBuf[10641] = 256'h5f026f0260026e0262022b02f90194013701c90062001f00e3ffacff8eff72ff;
    decBuf[10642] = 256'h39fff5fe91fe18fee8fdd9fd36febcfe80ff03004a003500faffc4ff93ffa2ff;
    decBuf[10643] = 256'h95ff89ff52ffd0fe53fec0fd5efd29fd18fd0afd32fd6efde7fd9afe40ff0300;
    decBuf[10644] = 256'hba0090011f02a202e9022a0316032803390365038d0399030a030b028b0026ff;
    decBuf[10645] = 256'h3efe14fe87fe36ff130069001b00a4ff0dffd2fe08ff79fffeff340065003800;
    decBuf[10646] = 256'h1000ecffcbffadff7fff24ffd0fe6dfe2afe36fe6dfedbfe60ffb9ffeaffdbff;
    decBuf[10647] = 256'h7dfff8fe7bfe6bfeb4fe47ff1f00af00fd00e600a5001b00c2ffd2ffffff7700;
    decBuf[10648] = 256'hc80012013a015e0169018701a301ab01a4018f0157011301c100740006009fff;
    decBuf[10649] = 256'h41ffecfee1fe13ff9cff4d002301ec013a0252023c02da018101ef003e0039ff;
    decBuf[10650] = 256'hfffdd8fccbfb63fb82fb12fc95fcdcfcf2fcdefcccfcfdfc82fd6afe47ff4a00;
    decBuf[10651] = 256'h3e011c02ab02fa027003dd033f04740485045804c503c6028c01110012ff87fe;
    decBuf[10652] = 256'h09fe2ffe0cfeecfd96fd7cfdf3fde1fe3d00de01f702900361038f021b026d01;
    decBuf[10653] = 256'h4d01f7007500feff3bff84fe0efecdfd08fe19fe2afee0fd68fdd5fc73fc61fc;
    decBuf[10654] = 256'hb3fc90fdecfe30005701170280029f02bc026e022602640179009bffd2fe84fe;
    decBuf[10655] = 256'h9bfe08ff6aff7cff6bff3fff4cffbaff9700f3013703b6032904c00322035902;
    decBuf[10656] = 256'ha201fc00390082ffdcfe70fe35fe6bfefdfed5ff9e0021013801cc004300a2ff;
    decBuf[10657] = 256'h0bffa8fe73fe42fe33fef0fd9cfd0dfd83fc4efc5efc00fd19fe73ffb700de01;
    decBuf[10658] = 256'h51022e02cf01b301cd01e501250239020302b20168015b019801e501ef017801;
    decBuf[10659] = 256'h840005ffa0fd15fd96fc09fdfdfddbfedeff8c0069013302e90231034603e402;
    decBuf[10660] = 256'h20026901c2002b00a2ff01ff3efe87fd40fd2afd3efd97fda8fd99fd8cfd98fd;
    decBuf[10661] = 256'he5fd67fe08ff74ffafffe4fff4ff5c00ef00c701900213035a03440309038c02;
    decBuf[10662] = 256'hfa0149017400aafff3fe4dfee1fd7ffd91fde2fd84fe1cffccff1400feffeaff;
    decBuf[10663] = 256'hfcff6e002e011902b7029a0218024201b2009800df0077010002ee017c01bd00;
    decBuf[10664] = 256'h06005fff1fffbcfe3ffe8dfde6fc24fca1fb89fb21fcf9fcfbfd35ff08002e00;
    decBuf[10665] = 256'h0b00acff56ff3cffb3ff750095015502bd029e0247026202d8029b0352046a04;
    decBuf[10666] = 256'hfd03d7020801d3ff2bff92fe63fee5fd25fd31fc93fbe9fbd4fc6ffe6800bc01;
    decBuf[10667] = 256'h76023d02700242021802f2018901eb00e8ffaefe87fd14fdf1fc8ffd1ffed6fe;
    decBuf[10668] = 256'h4dff37ff24ffeefefefe48fff6ff9c005f01ad01c501af014d01d0007f005200;
    decBuf[10669] = 256'h2a000600cfffc5ffceff180086000b0141013001c9001b00a5ff64ff77ffadff;
    decBuf[10670] = 256'hdeffb1ff39ffc7fe7efea6fe43ff3100cf005f01ad01240290024103b803f903;
    decBuf[10671] = 256'h96038a02e4005bfff6fd0efd3cfcc9fba6fb86fbdcfb93fc99fdd2fea5ff6500;
    decBuf[10672] = 256'h8800680012002c001400ffff9dff43ff33ff9aff63009f01c9015601d6ff71fe;
    decBuf[10673] = 256'ha0fe6f00920390068208720733056701d0fe67fdd5fd38fe48ff9aff4fff0bff;
    decBuf[10674] = 256'h49ff81ffb4ffe3ff64ffa4fe6afdecfc5ffddffe10011b036f043a03f0ffb5fb;
    decBuf[10675] = 256'hb9f722f58bf665fa160064057607d506fd035d0012fdcafb2dfc3dfd7dffb302;
    decBuf[10676] = 256'hd6045608b00af80bce0aea063000c5f9eff3a9f1baf39dfade026a086c09d604;
    decBuf[10677] = 256'h00ff2ef86ef544f60efae0fe82044c085e0abd09080869041e0169fc08f852f6;
    decBuf[10678] = 256'hd7f612fb5601d608e10da110770c2104edf7cdef6be8c3e9ddefd9f9ed050d0e;
    decBuf[10679] = 256'h7b12d213b80dbc0357faccf178ee7befe6f566fd7f08e10fe813b012240d1406;
    decBuf[10680] = 256'hd3fd0ff608f31ef29ef4ecf91f00f505bf096f0a4e072e02fbfb25f6dff38ff4;
    decBuf[10681] = 256'hf1f858006c09860fda12d30f6809e801dcfc47f871f733f8e4f884f916faa3fb;
    decBuf[10682] = 256'hfdfdfc00ed0248036300e4fc99f92cf9e4fb3201fc040d076d067002c8fde7fb;
    decBuf[10683] = 256'h9cfd3c0177052c07b107570559022e018901c803a904dd033e0096fb34f77ff5;
    decBuf[10684] = 256'h03f64ef971fb9cfcf6fc5bfb7bfabffaebfcb6005604a107c409280acd093208;
    decBuf[10685] = 256'h5207860651053804a10173fe74fbbcf8acf7a3f819faf5fb29fd62fd2ffd5dfd;
    decBuf[10686] = 256'hdbfd35ff7900f4018d025f02e1016e0179009cffd3fe1cfe76fd8bfdedfdfafe;
    decBuf[10687] = 256'h53009801be02320354033503a50222027c018e00f0ff27ffd9fef0fe31ff6cff;
    decBuf[10688] = 256'ha2ffb2ffa3ff1c000f014902c403c3049504c203cf016bffd0fd5afc8efb51fb;
    decBuf[10689] = 256'h19fbe6fa14fb92fb52fcd2fd37ff7b00fa00870093ff37fe4ffdcdfdc0ff2402;
    decBuf[10690] = 256'h080533068d06f2047c03a001e700af004801d301a9018301d40036001900ffff;
    decBuf[10691] = 256'he7ff7bffa3fe2efdc9fb84fa06fa12fb1dfd54007702a203fc03610256007afe;
    decBuf[10692] = 256'h45fd7dfd16feb7ffd000cf01b70235030f03a6028a013000ecfec5fd9efd07fe;
    decBuf[10693] = 256'h24ff30002401c30119023302ec01fe00e1ff88fe43fd19fd8cfdc6feedffad00;
    decBuf[10694] = 256'hd000320068ffb1fe3bfe50fe8bfee5fe36ff9dff1500a8000a011c01ca002800;
    decBuf[10695] = 256'hbcfff7ffdf007a0203046805f30575051c047a028100a5fef5fc6cfb6dfa85f9;
    decBuf[10696] = 256'h5bf91bfa55fb24fdd4fe5d00c2014d02cc02f202cf02b0025902d70131011700;
    decBuf[10697] = 256'h0bff5cfebefda2fd24fefafec3ff4600bd00d200e600d400c4000d0186011802;
    decBuf[10698] = 256'hc902e00249022301fffef4fca0fbe7fa8ffb5afd0aff930092017a02a4027e02;
    decBuf[10699] = 256'ha10202023901e6ffa1fe26fd8dfc18fd93fef8ff990142020f02ca00a3ff97fe;
    decBuf[10700] = 256'h74fe51ffc7002c02140392036c03030365026201280002ff5bfd43fc44fbb9fa;
    decBuf[10701] = 256'h37fbf7fbebfc08fec8febcff5a002301da015102660204026301cc00b8003501;
    decBuf[10702] = 256'hc80151021b0248010c0039ffc6fe2fff8b00cf01a202c80260024301360042ff;
    decBuf[10703] = 256'h65fe0ffec0fd79fd38fdfdfc33fda5fd82fe9fffab005a017901e900caff0aff;
    decBuf[10704] = 256'ha2fe00ff0300f700560100011500f8fe38fe5bfe78ff8400790117023302e501;
    decBuf[10705] = 256'hcd01e30145029e02af0247027f01b600caff6cff4fff9dff1400feff4eff19fe;
    decBuf[10706] = 256'h9efc39fbaefa84fa43fbc3fc28fe6dff3f00ff00ae018b021b03d203e9037d03;
    decBuf[10707] = 256'ha502a301ae00500033008100c8000901ce007500e3ff59ffdcfe4afee8fdd6fd;
    decBuf[10708] = 256'he6fd4efe16ff19000d01ab01c8017a01a400dbff24ffadfe6cfe58fe23fe13fe;
    decBuf[10709] = 256'h5cfe0affe0ffe3004b016b01db0059001100270089002a019601d1019b014a01;
    decBuf[10710] = 256'h0001a3001d007cffe5fe34febefdfffdaffee4ff0b011702c602e5028f020d02;
    decBuf[10711] = 256'h07011300b7fe73fd4cfc3ffb1cfb7bfb7efcfefd63ff4a0071013102e002ff02;
    decBuf[10712] = 256'he2026002ba014d01eb00fd004e0198017001eb002600a3ff2dff17ff2bff3dff;
    decBuf[10713] = 256'h0cffa5fe47fe0afe15fe6ffedcfe44ffa1ffadffa2ff84ff45fffafedcfef8fe;
    decBuf[10714] = 256'h52fff0ffb3006a01e00121028302b9020a03fb02b9020302e300d7ffe3fe84fe;
    decBuf[10715] = 256'ha0feeffe66ffa6ff93ff39ffc8fe7efe71fe95fee2fe50ff1000fb00d8012e02;
    decBuf[10716] = 256'h14026e012a0088fe70fd71fc42fc6cfce0fc8efd6bfea8ff23018802cc034b04;
    decBuf[10717] = 256'h2404760399020902ef01d701ed01b2013501a200f2ff4bff5efebffd30fd4afd;
    decBuf[10718] = 256'h91fd54fe0bff81ff6cffe2fe1efe9bfd83fdeffdc7fecaffbe005c01b3010102;
    decBuf[10719] = 256'h480289029d0267021602af011b0192005c002c003a002d002100eaff90ff3bff;
    decBuf[10720] = 256'h04ff22ff74ffd7ff35002900b0ffbcfec8fdeafc5bfca9fcaefda2febfffcc00;
    decBuf[10721] = 256'h34019301e90104021b02af01ff00f9ff4bffecfe42ff2d00cc00220108019100;
    decBuf[10722] = 256'hfaff97ffa9ff3c00c5004201730182015901350114010a01dc00b30070003000;
    decBuf[10723] = 256'he6ffa0ff3bffdefe58feb7fd4bfde9fcd7fc28fdadfd4efe11ffc8ff3e00aa00;
    decBuf[10724] = 256'h97003d00ecff67ff0eff1eff86ff33000901d201be025c03b203980380031403;
    decBuf[10725] = 256'h8b020d029c013401bc00090034ff31fef7fcd0fb10fba8fa88fadefac9fb64fd;
    decBuf[10726] = 256'h5eff3a01ea0202049b0410043e037e021502b601600112016b00a9fff2fe4cfe;
    decBuf[10727] = 256'he0fd1afe74fe06ff68ff9effefff3900cc0055018b013a015c00c1fe38fd39fc;
    decBuf[10728] = 256'haefbd8fbe5fc1ffe46ff9f008701050279029b02bb029e025002380223020f02;
    decBuf[10729] = 256'hb6014401bf001e0087fffdfe80feeefd8cfd56fda8fd67fe87ffe0002502f702;
    decBuf[10730] = 256'hb7039403350333023f01e3fffbfe28feb5fd4cfdeefc97fc49fc31fc9dfc75fd;
    decBuf[10731] = 256'hb1fed8ff9800bb009b007f00990010017c01de01f0019e013701da00e6003301;
    decBuf[10732] = 256'hc9016002110358034203b902f401d500c8ff1aff3dfeadfd2afd54fc8bfbd4fa;
    decBuf[10733] = 256'h8dfaf9fa20fceffd1b009001e4029e03660399036a0340036603fe029f020f02;
    decBuf[10734] = 256'h8d011601d5007300f6ff22ff20fe2cfd8dfc71fcbffc36fda2fd04fe5dfecffe;
    decBuf[10735] = 256'h71ff3400b700fe00e80086002d00fcffd0ffddffd1ffc6ffbcffd7ff11005500;
    decBuf[10736] = 256'ha700f4003a018c01d9010b021402ca0134017100efffa7ffbdff1f0078008900;
    decBuf[10737] = 256'h5c001a00c5ffd0ff2a00c7005f019a016401d200faff31ffaefe37fecbfd42fd;
    decBuf[10738] = 256'ha1fc09fca7fb95fbe7fba6fc92fdaefebbff690007015e01ac01c4013002b902;
    decBuf[10739] = 256'h3603a8030f0437042b04f4038603e402cb0172002dffb2fd4dfcc2fb98fb57fc;
    decBuf[10740] = 256'h06fd22fee2fe4bff6bff4eff68ffafff1b007d00fb002b011d012a0136018301;
    decBuf[10741] = 256'hc901f701cd016c01d900770041005100430000007affb6fe33feecfd01fe3cfe;
    decBuf[10742] = 256'h96fea6fe7afe37fe12fe33fec9fe8cffab00b80121024002ea01cb00beffcafe;
    decBuf[10743] = 256'h2cfe49fefffea6ff3d009f00b100c100ee0030018501bc01c601ab01b3010602;
    decBuf[10744] = 256'h7f02d002c1021302df0063ff64fe36feb4fe28ffd6fff6ffd9ff8aff43ff02ff;
    decBuf[10745] = 256'hc7fe27fe39fd5bfc05fc88fcbcfd38ffd1ffffff81ff27fe9cfdc6fd86fec0ff;
    decBuf[10746] = 256'h3b013a022203a003c703a4038403f4027202cc013401f900e700d700ab003300;
    decBuf[10747] = 256'h5fff96feabfd4cfd2ffd7efd53fe56ff4a0028017e01980180019601aa01df01;
    decBuf[10748] = 256'hcf018501bd00baff0bff6dfe17fe31fe49fe33fef8fdc3fdb3fdfcfdaafeafff;
    decBuf[10749] = 256'h5e00fc0052016c0155016a01a501fe012f02030270019800cfffe4fe45feb6fd;
    decBuf[10750] = 256'h9cfd84fdc5fd4efe13ffcaff7000b1009d008b007b00c500080144017b015d01;
    decBuf[10751] = 256'h42014a017f01ca01100207028b01c700dcff3dff21ff6fff1500ad000f01fd00;
    decBuf[10752] = 256'h8b00e9ff52ffeffebafe89fe3ffec7fd55fd29fd51fd07fef2fe90ffadff5fff;
    decBuf[10753] = 256'hb8fe4cfe60fe01ffefffcc005c017601ff00be008300b9002b0174019d017801;
    decBuf[10754] = 256'h2b01e500ca00d200da00ee00e800c100920067003f001100d9ff95ff56ff4dff;
    decBuf[10755] = 256'h73ffdaff9a005101c701b2015001af00c1ff23ff93fe10fec9fdb3fda0fdd5fd;
    decBuf[10756] = 256'h47feaefef1fee5fe82fe25fe18fea7feceff9d01d2027a0347035f0239017900;
    decBuf[10757] = 256'hcaff2cff9cfe1afe74fd5efdc0fda8fec5ff3800a10081002b0045008c002401;
    decBuf[10758] = 256'hd4011c025c0249021302e201b601a9019d0192016001fb00680090ff8efedffd;
    decBuf[10759] = 256'hc0fd16fe01ffdeffe1004a016901da0023004dff84fecdfd56fdeafcd6fc0cfd;
    decBuf[10760] = 256'h3dfd86fdfffd91fe42ff1700a700c100aa003d00b4ffa2ffd3ff75000d019601;
    decBuf[10761] = 256'ha80198016b0193010102680290025302ae01a9004000600029014902a2032d04;
    decBuf[10762] = 256'h0304aa024f000ffe6efb5ffa68f948fa9cfb4dfd46ff9a0053011b0182009aff;
    decBuf[10763] = 256'h73fe00fe69fe46ffbc00bb014602c7010801ceff4fff29ff92ff6f00ff008101;
    decBuf[10764] = 256'hf801bb023d03b40373037402f40029fff5fd4cfd7ffdaefd84fd10fd1cfc00fb;
    decBuf[10765] = 256'h8dfaf5fa12fcb8fdb1ff8d013d035604ef04c104420482038e02f001d301ed01;
    decBuf[10766] = 256'h3502760213024f012f0023ff74fe55fe1eff720013029c030105d3045703c000;
    decBuf[10767] = 256'h92fd93fa69f959f8acf88cf9d0f90efad6f909fa94fabbfb61fdeafe4f009301;
    decBuf[10768] = 256'hba021304b5053e07d7074c072506e5034a02d4009000ce00060139010b018c00;
    decBuf[10769] = 256'h6600430063007f009900b100c700da00ec009b00beff62fec1fc38fb9ffacdfa;
    decBuf[10770] = 256'ha0fbf9fce1fdb4fedafeb7fe97fe7bfec9fe6fffb400f80173037204a1042204;
    decBuf[10771] = 256'h1603dc010901960073005400fdff7bffd5fe68fe2efe1cfeebfda1fd44fd07fd;
    decBuf[10772] = 256'h80fd74fe39006e01860253022502a70134011101f1009b00180042ffb3fe99fe;
    decBuf[10773] = 256'he0fe4cffaeff9cff8cff9bff1300070141021303d303f603970307038502df01;
    decBuf[10774] = 256'h7201e9006c0099ff96fe5cfd89fc7dfb14fb34fb51fb6bfb53fb12fb26fb7ffb;
    decBuf[10775] = 256'h52fc8ffdb5fe75ff240001013d02b8031d0505062f06bc050e0570041a04ff03;
    decBuf[10776] = 256'hb803f602a2015d0036ff77fe54fe73fe57fe71fe29fe3ffe53fe65fe95fea4fe;
    decBuf[10777] = 256'h97fe8bfe96fedcfe2eff91ffb9ffadffa2ff70ff30fff6fec2fed6fe34fffdff;
    decBuf[10778] = 256'h7201d70262038d031903250287013101e300fa00b90030006bff80fea3fddafc;
    decBuf[10779] = 256'h23fc7dfb10fb24fba1fb95fc15fee0ff9001a802a70333045d043604ce036f03;
    decBuf[10780] = 256'h19039602f0010201a6ff61fe8ffd68fd17fe33ff400034019301760128014001;
    decBuf[10781] = 256'h5501df015c028c026002b201ad0073ff4cfe40fd91fcb4fb24fbd6faeefa2efb;
    decBuf[10782] = 256'h91fb31fcc9fc04fd39fd6afdd1fd9afe1000db0106047c05d0060e0746074706;
    decBuf[10783] = 256'h020533038301faff61ff33ff5dffd0ff7e009e004800f9ffb2ff71ff5dff93ff;
    decBuf[10784] = 256'he4ff4c0074004f00c0ff9afe73fd1afc32fb08fb7bfb6ffccbfdb3fedaff9900;
    decBuf[10785] = 256'h8e012c0282029c02b40273021102db018a012301aa0018008fff59ff69ffd1ff;
    decBuf[10786] = 256'h49009a00a9006600f9ff92ff6aff76ff81ff9fffa8ffb0ff8bff23ff81fe93fd;
    decBuf[10787] = 256'hb6fc26fc0cfce2fc1efe99ff98008001fe0172022003be034e049c0484041804;
    decBuf[10788] = 256'hb6033903c702250237015a0057ffa9fe4afe2dfe47fe2ffe45fe80feb6fec6fe;
    decBuf[10789] = 256'hb7fe74fed7fd3ffdddfccbfc1cfd66fd74fd1ffd7afc74fb0cfb2bfb68fc8bfe;
    decBuf[10790] = 256'h2c01a603410521066506ac05740541056f05990573057f046203550261010201;
    decBuf[10791] = 256'hac002a0024ff30fe53fdc3fcddfc83fdf0fd03feaafd59fd0ffd37fdbcfd81fe;
    decBuf[10792] = 256'h04ff4bff35ffacfee7fd65fdeefc03fdb4fdb9fef3ff1a0127028f02af02cc02;
    decBuf[10793] = 256'hb202f90265033d040605bd0534061e066d053904150274fffbfcbbfab0f86cf8;
    decBuf[10794] = 256'haaf852f9ebf9d3fa51fb11fcbffcdcfd35ffd700ef0154033c040f058205a505;
    decBuf[10795] = 256'hc80418036801dfff46ff18ff96ff09007200d100ee007001e7017e022f037603;
    decBuf[10796] = 256'h350385025001d5ff70fecefcb6fbb7fa2cfaadf987f9f0f98efa90fbcafcf1fd;
    decBuf[10797] = 256'hfefe66ff86ffdcffc700e4013d032504a4047d045a04bc032d03de026702fb01;
    decBuf[10798] = 256'h990187019801a601990175011201b4005f006a008800b600be007a00f2fff2fe;
    decBuf[10799] = 256'hb9fd92fc38fbadfa2ffaa2fa50fb2efcbdfc0cfd83fd45fe99ff97017303a804;
    decBuf[10800] = 256'h500551040c03e60126014901e7017602c5024e02b7012d01d400e400d5009300;
    decBuf[10801] = 256'hf5ff07ff2afe9afd17fd00fd15fd02fd13fde3fcd4fcfcfc51fdf6fd2bffa600;
    decBuf[10802] = 256'h0b024f032204fc03d903fb026c02e901d101e701fb01c5015301b1001a00dfff;
    decBuf[10803] = 256'hf1ff42008c006300f6ff37ffb4fe6dfe82febdfef3fec2fe20fe5dfd0ffdf7fc;
    decBuf[10804] = 256'h38fdc1fdf7fde7fd9dfd3ffd03fd3afdd0fd14ffb500af028b043b06e3061607;
    decBuf[10805] = 256'h8b060d06000552043503dc019700c8fe93fdebfc52fc80fcaafc1dfdccfda9fe;
    decBuf[10806] = 256'hacff5a0037018e017401fd009100e0ff0affcefda7fc4efb66fae8f9a7fae1fb;
    decBuf[10807] = 256'h5cfd27ffd800f00155039a04c1051a07a507cf075c07ae0652050d049202c700;
    decBuf[10808] = 256'h9cfe90fcb4fa80f9d7f8a4f82ff9aef9bafaaefbcbfcd8fd57ffbc0001022803;
    decBuf[10809] = 256'he80350047004e003f5029901550082ff75fe0dfeedfd7dfe68ffc40065027e03;
    decBuf[10810] = 256'hb10382035803e502c202e202ff027c027701f7ff92fe4efd7bfc08fc59fbbbfa;
    decBuf[10811] = 256'h2cfa11fa59fa47fb63fc70fd1efebcfe13ff95ff0c00fa00d701a0028c032a04;
    decBuf[10812] = 256'h80046604ef032c0341026401d4001d0077ff0bffd0fee2fe74ff730067014502;
    decBuf[10813] = 256'h9b0281023a02f90197013d01ab00acffb8fe9bfddbfcb8fcd8fcbbfc6dfc97fb;
    decBuf[10814] = 256'h5bfa34f974f897f8f3f9f1fb55fe9500a002f403ad04e5041805470571059705;
    decBuf[10815] = 256'h000620063c062206ab05be04e3027f003ffe34fce0faa2fadbfa74fb5bfc86fc;
    decBuf[10816] = 256'h5ffc3cfc9efb81fbd0fb47fc09fdc0fd66fed2fe0dff1fff50ff9aff2d00dd00;
    decBuf[10817] = 256'he301d702b4030a045904410457046a04a004d104df049d04170453039c022502;
    decBuf[10818] = 256'h8e01b60040ff75fd49fb3ef962f7a9f6e1f614f7fcf77af8edf89cf9f7faf6fc;
    decBuf[10819] = 256'h5aff3e02f6040606fd06b206e6052d05140415032d0206019300e5ffc5ffa8ff;
    decBuf[10820] = 256'h8eff05009c0074017702b1038304aa048704aa036d024601edffa8fed6fd16fd;
    decBuf[10821] = 256'h68fcc9fb3afb83faddf91af963f8ecf7d7f787f8bcf98bfb3cfda5ff4001b602;
    decBuf[10822] = 256'h0a04c3046c059f05cd054b060b07ff075e08420822072f05cb02300125ff59fe;
    decBuf[10823] = 256'ha0fd67fdcefca0fc76fc50fc2dfc4cfcf6fba8fb31fbf0fa2bfb84fb17fca0fc;
    decBuf[10824] = 256'hf9fc2afd56fd7efd04feecfe4800e90172033d05f7059f06d206a406d1055e05;
    decBuf[10825] = 256'h3b05dc04bf04a5042e046c03180277007efea2fcf1fa69f9d0f844f81af841f8;
    decBuf[10826] = 256'ha9f808f998f94ffaf5fab8fb6ffc74fdaefe29005a026504b905ee0626078d06;
    decBuf[10827] = 256'h02062f05230474039702ce014b010401980084007200620071007e008a003d00;
    decBuf[10828] = 256'ha7ff8efe35fd4dfc7afba0fb09fc26fde6fd08feaafde0fcc1fbb4fa4cfa2cfa;
    decBuf[10829] = 256'hf5fa15fcbbfd44ff7501ea023e04f804a0053906c40643071c0728060b05b203;
    decBuf[10830] = 256'h1102f80093fff2fd69fc04fbbff941f9b4f9a8fac5fb1efda9fd28fe9bfe03ff;
    decBuf[10831] = 256'ha1ff6b00560175015901a2006dff9afedbfdb8fdd7fd2efeb0fe56ff19000401;
    decBuf[10832] = 256'he201ab022d034503300343037903aa0311040304af030a03a501daff2afe31fc;
    decBuf[10833] = 256'hddfaa8f990f8f7f76bf796f709f8b7f8d4f92dfbcefc57fe2200d3013c047c06;
    decBuf[10834] = 256'hf107450983096b08a006740469028d00dcfec4fd2bfda0fc1efddefdd2feefff;
    decBuf[10835] = 256'hfb00aa01c9017301f0007a003900afffebfecbfd25fc9cfa9df9b5f88bf8fef8;
    decBuf[10836] = 256'hf3f90ffb69fc0afe0300df0114039d0436056405e2055606be06de06c1063e06;
    decBuf[10837] = 256'h0a058f03c4018f0006ffa1fd5cfc35fb76fa0dfa2dfabcfadcfb35fd1dfe44ff;
    decBuf[10838] = 256'h0400b2008f015902db025203e602e70167009cfeecfcd3fba0fbcffba1fcaefd;
    decBuf[10839] = 256'he8fe0f001b019b020004e8046605d905b60558053b0521056805520517052f04;
    decBuf[10840] = 256'h94029b0037fe53fb61f99df7a6f6f1f6bdf76df9f6fac1fc71fefafff9008401;
    decBuf[10841] = 256'h020229024c02aa023a03bd033404f30342033d020301dcff69ff46ffe4ffad00;
    decBuf[10842] = 256'h010246036d04c605ae06d806fe065006f40453035a01f6feb6fcabfa57f919f9;
    decBuf[10843] = 256'h51f984f90ffa39fa13fa36fa95fa5efbe6fc4fff3302250434052b06e0051405;
    decBuf[10844] = 256'h5b04b3038003510327034e037003cf03260440049903ac0250010b00e4fe24fe;
    decBuf[10845] = 256'h8dfeaaff03014802c602a002ab0150000bffe4fdbefde1fd3ffe23fe6cfd67fc;
    decBuf[10846] = 256'h2dfb06fa93f941fa5efb51fda5fe5500fd00960121024803ee04e706c308740a;
    decBuf[10847] = 256'h1c0bb50b870b080baf09b107c50445010afd31faa4f82bf899f8fcf80cfa03fb;
    decBuf[10848] = 256'h4dfb91fbcffbe8fce7fd2bff52005f010d02ee019701e0003a004cffedfe97fe;
    decBuf[10849] = 256'hb1fef9febbff0f010d0371055508470aa10a4f0a6f090b076f05fa032e037402;
    decBuf[10850] = 256'hcc01cd0088ff0dfea8fcc0fbeefae1f9a7f880f774f651f66ef714f97dfb61fe;
    decBuf[10851] = 256'h1a01de027a045a059e05dc0533059a040f04e5037203950375035803d6028e02;
    decBuf[10852] = 256'h4e02880206039803fa0330041f04b8034003ce024902850199007dff23fedffc;
    decBuf[10853] = 256'hb8fbf8fa4afaebf9cef9e8f92ffa9cfa73fb76fc6afd87fee0ffc8004302a803;
    decBuf[10854] = 256'hed0414066d07550828099b09be099e094809c50890071506e403d90175ffdafd;
    decBuf[10855] = 256'hfafc2efc74fbccfa33faa8f929f950f9fef91bfb74fcb9fde0feecff9b003901;
    decBuf[10856] = 256'hc9014b02c202030316034c037d03e4035c04ef042a053b05a904d10308038502;
    decBuf[10857] = 256'h9d02b6035c05e5064a087908a607b3054f036b00b2fd39fbf9f8eef612f5ddf3;
    decBuf[10858] = 256'ha5f33ef483f5fef695f90efc97ffe202e00599085d0a540b9f0b5b0ba10af909;
    decBuf[10859] = 256'h94089606ba048e0283002ffffafdc2fdf5fd80fe53ffac004e02d603d5040405;
    decBuf[10860] = 256'h85042c038b0102009dfefbfce3fb18fae3f8caf731f7bdf7e3f88afa83fc5ffe;
    decBuf[10861] = 256'h8a000002dc038c058607da088a0aa20b3b0c0d0ce30bd60a57098c07e4046b02;
    decBuf[10862] = 256'h87ffcefc55fa5ef97ef8c2f87bf923fabcfa47fbc6fb86fcc0fd3bff0601b602;
    decBuf[10863] = 256'hcf0368043904bb03fb02070229016000deff37ffcbfe90fec6fe58ff57004b01;
    decBuf[10864] = 256'ha70249046105c60668088009190a480a7509cf07d60572038e00d5fd5cfbc0f9;
    decBuf[10865] = 256'h4bf87ff7c5f6adf57af505f6d7f6caf82efb6efd0f00d301ca0240040c05c505;
    decBuf[10866] = 256'h6d06060792076707a8066e054704ed026202e401be019b01fa0150023b031804;
    decBuf[10867] = 256'he2046405ed04a90308029eff03fe8dfc39fb80fa67f902f81bf7f4f59af4dff5;
    decBuf[10868] = 256'h57f8a4fd66fe17ffb7ff4900c4ff3d00cfff3300d8ff2a00e0ff2400e6ff1e00;
    decBuf[10869] = 256'hebff1900efff1600f3ff1200f6ffdbfff3ffdefff1ff0300f3ff02000f000300;
    decBuf[10870] = 256'h0e001800fcff0500fdfff6ff09000300feff0300fffffbfffefffbfffeff0100;
    decBuf[10871] = 256'h03000e001400150011000000f5fff3ffebfff0fffafff6fff5fff8fff3fff4ff;
    decBuf[10872] = 256'hf7fff4fff7fffbfffcff04000300040011001700150020002200180017001100;
    decBuf[10873] = 256'h08000700fffffafff8ffeeffe7ffe3ffe0ffe5ffe6ffe3ffe9ffeefff6ff0600;
    decBuf[10874] = 256'h0e001000120013000f00130012000e000d000600faffefffe5ffe9fff6ffffff;
    decBuf[10875] = 256'h01000200feff02000a000f001000110010000300f9fff7fffcfffdff04000a00;
    decBuf[10876] = 256'h0b000a0008000200fcfffbfffdfffefff8fff7fffcff00000300050006000c00;
    decBuf[10877] = 256'h0a00fcfff6fff5fff3fff5fff6fff7fff6fff3fff4fff7fff4fff7fff9fff5ff;
    decBuf[10878] = 256'hf2fff8ff000006000d000c000d0015001d0020001f001e001d0012000300fdff;
    decBuf[10879] = 256'hf8fff3fff1ffeaffe4ffe3ffe6ffeaffedfff5ff01000d000b00150016000e00;




    $display("Done initializing");

  end

  //---------------------------------------------------------------------------------------
  // test bench implementation
  // global signals generation
  always @(posedge clk) begin
    mCtr <= mCtr + 1;

    if (testCount >= TESTS_TO_RUN) $finish(1);

    case (mainState)
      MAIN0: begin
        rst <= 1;

        inDone <= 0;
        encDone <= 0;
        decDone <= 0;

        if (mCtr >= 2) begin
          $display("");
          $display("IMA ADPCM encoder & decoder simulation");
          $display("--------------------------------------");
          mCtr <= 0;
          mainState <= MAIN1;
        end
      end

      MAIN1: begin
        rst <= 0;

        mCtr <= 0;
        mainState <= MAIN2;
      end // case: MAIN1

      MAIN2: begin
        if (inDone && encDone && decDone) begin
          $display("Test %d done!. mCtr: %d", testCount , mCtr);

          testCount <= testCount + 1;
          mCtr <= 0;
          mainState <= MAIN0;
        end
      end

    endcase // case (mainState)
  end

  //------------------------------------------------------------------
  // encoder input samples read process
  always @(posedge clk) begin
    iCtr <= iCtr + 1;
    if (rst) inState <= IN1;

    case (inState)
      IN0: begin
        iCtr <= 0;
      end

      IN1: begin
        // clear encoder input signal
        inSamp <= 16'b0;
        inValid <= 1'b0;
        // clear samples counter
        sampCount <= 0;
        inBytesRead <= 0;

        // binary input file
        inIdx <= 0;

        if (!rst) begin
          iCtr <= 0;
          inState <= IN2;
        end
      end // case: IN1

      IN2: begin
        if (iCtr >= 50) begin
          // read input samples file
          intmp <= inBuf[inIdx][(BUFFER_BYTES << 3) - 1:(BUFFER_BYTES << 3) - 8];
          inBytesRead <= inBytesRead + 1;

          $display("inBuf[%d] = %h%h%h%h%h%h%h%h", inIdx,
                   inBuf[inIdx][255:224],
                   inBuf[inIdx][223:192],
                   inBuf[inIdx][191:160],
                   inBuf[inIdx][159:128],
                   inBuf[inIdx][127:96],
                   inBuf[inIdx][95:64],
                   inBuf[inIdx][63:32],
                   inBuf[inIdx][31:0]);


          iCtr <= 0;
          inState <= IN3;
        end
      end // case: IN2

      IN3: begin
        // Stop looping through inputs if eof
        if (inBytesRead >= TOTAL_IN_BYTES) begin
          $display("Reached eof of input");

          iCtr <= 0;
          inState <= IN5;
        end

        else begin
          if (iCtr == 0) begin
            // read the next character to form the new input sample
            // Note that first byte is used as the low byte of the sample
            inSamp[7:0] <= intmp;

            case (inBytesRead % BUFFER_BYTES)
              1:  inSamp[15:8] <= inBuf[inIdx][247:240];
              3:  inSamp[15:8] <= inBuf[inIdx][231:224];
              5:  inSamp[15:8] <= inBuf[inIdx][215:208];
              7:  inSamp[15:8] <= inBuf[inIdx][199:192];
              9:  inSamp[15:8] <= inBuf[inIdx][183:176];
              11: inSamp[15:8] <= inBuf[inIdx][167:160];
              13: inSamp[15:8] <= inBuf[inIdx][151:144];
              15: inSamp[15:8] <= inBuf[inIdx][135:128];
              17: inSamp[15:8] <= inBuf[inIdx][119:112];
              19: inSamp[15:8] <= inBuf[inIdx][103:96];
              21: inSamp[15:8] <= inBuf[inIdx][87:80];
              23: inSamp[15:8] <= inBuf[inIdx][71:64];
              25: inSamp[15:8] <= inBuf[inIdx][55:48];
              27: inSamp[15:8] <= inBuf[inIdx][39:32];
              29: inSamp[15:8] <= inBuf[inIdx][23:16];
              31: inSamp[15:8] <= inBuf[inIdx][7:0];
              default: $display("Unexpected number of bytes read for inSamp");

            endcase // case (inBytesRead % BUFFER_BYTES)

            // until next clock tick, inBytesRead is still previous value
            inBytesRead <= inBytesRead + 1;
          end // if (iCtr == 0)

          if (iCtr == 1) begin
            // sign input sample is valid
            inValid <= 1'b1;

            if ((inBytesRead % BUFFER_BYTES) == 0) begin
              inIdx <= inIdx + 1;

              $display("inBuf[%d] = %h%h%h%h%h%h%h%h", inIdx + 1,
                   inBuf[inIdx][255:224],
                   inBuf[inIdx][223:192],
                   inBuf[inIdx][191:160],
                   inBuf[inIdx][159:128],
                   inBuf[inIdx][127:96],
                   inBuf[inIdx][95:64],
                   inBuf[inIdx][63:32],
                   inBuf[inIdx][31:0]);

            end // if ((inBytesRead % BUFFER_BYTES) == 0)

            // Prepare for next state
            iCtr <= 0;
            inState <= IN4;

          end // if (iCtr >= 1)

        end // else: !if($eof(instream))

      end // case: IN3


      IN4: begin
        // update the sample counter
        if (iCtr == 0) begin
          sampCount <= sampCount + 1;
        end


        // wait for encoder input ready assertion to confirm the new sample was read
        // by the encoder.
        if (inReady) begin
          //$display("Sample count: %d, iCtr: %d", sampCount, iCtr);

          // read next character from the input file
          case (inBytesRead % BUFFER_BYTES)
            0:  intmp <= inBuf[inIdx][255:248];
            2:  intmp <= inBuf[inIdx][239:232];
            4:  intmp <= inBuf[inIdx][223:216];
            6:  intmp <= inBuf[inIdx][207:200];
            8:  intmp <= inBuf[inIdx][191:184];
            10: intmp <= inBuf[inIdx][175:168];
            12: intmp <= inBuf[inIdx][159:152];
            14: intmp <= inBuf[inIdx][143:136];
            16: intmp <= inBuf[inIdx][127:120];
            18: intmp <= inBuf[inIdx][111:104];
            20: intmp <= inBuf[inIdx][95:88];
            22: intmp <= inBuf[inIdx][79:72];
            24: intmp <= inBuf[inIdx][63:56];
            26: intmp <= inBuf[inIdx][47:40];
            28: intmp <= inBuf[inIdx][31:24];
            30: intmp <= inBuf[inIdx][15:8];
            default: $display("Unexpected value");

          endcase // case (inBytesRead % BUFFER_BYTES)


          // use sampCount because you inReady occurs at an unknown time count
          inBytesRead <= (sampCount << 1) + 1;

          iCtr <= 0;
          inState <= IN3;
        end

      end // case: IN4

      IN5: begin
        // sign input is not valid
        inValid <= 1'b0;

        if (iCtr >= 1) begin
          inDone <= 1;

          iCtr <= 0;
          inState <= IN0;
        end
      end // case: IN5

      default: inState <= IN0;
    endcase // case (inState)

  end // always @ (posedge clk)


  // encoder output checker - the encoder output is compared to the value read from
  // the ADPCM coded samples file.
  always @(posedge clk) begin
    eCtr <= eCtr + 1;
    if (rst) encState <= ENC1;

    case(encState)
      ENC0: begin
        eCtr <= 0;
      end

      ENC1: begin
        // clear encoded sample value
        encCount <= 0;
        encBytesRead <= 0;

        // open input file
        encIdx <= 0;


        // wait for reset release
        if (!rst) begin
          enctmp <= encBuf[encIdx][(BUFFER_BYTES << 3) - 1:(BUFFER_BYTES << 3) - 8];
          encBytesRead <= encBytesRead + 1;

          $display("encBuf[%d] = %h%h%h%h%h%h%h%h", encIdx,
                   encBuf[encIdx][255:224],
                   encBuf[encIdx][223:192],
                   encBuf[encIdx][191:160],
                   encBuf[encIdx][159:128],
                   encBuf[encIdx][127:96],
                   encBuf[encIdx][95:64],
                   encBuf[encIdx][63:32],
                   encBuf[encIdx][31:0]);


          eCtr <= 0;
          encState <= ENC2;
        end
      end // case: ENC1

      // encoder output compare loop
      ENC2: begin
        if (encBytesRead >= TOTAL_ENC_BYTES) begin
          $display("Reached eof of encryption file");
          eCtr <= 0;
          encState <= ENC4;
        end

        else begin
          encExpVal <= enctmp;

          // wait for encoder output valid
          if (encValid) begin
            if (!decReady) $display("Encoder output too quickly into decoder!!!");


            eCtr <= 0;
            encState <= ENC3;
          end
        end // else: !if($eof(encstream))

      end // case: ENC2

      ENC3: begin
        // compare the encoded value with the value read from the input file
        if (encPcm != encExpVal) begin
          // announce error detection and exit simulation
          if (eCtr == 0) begin
            $display(" Error!");
            $display("Error found in encoder output index %d.", encCount + 1);
            $display("   (expected value 'h%h, got value 'h%h). encIdx: %d, inIdx: %d, decIdx: %d", encExpVal, encPcm, encIdx, inIdx, decIdx);            

          end

          // wait for a few clock cycles before ending simulation
          if (eCtr >= 20) $finish();
        end // if (encPcm != encExpVal)

        else begin
          //$display("encoder output correct. expected %h, got %h", encExpVal, encPcm);

          // update the encoded sample counter
          if (eCtr == 0) encCount <= encCount + 1;

          // delay for a clock cycle after comparison
          if (eCtr == 1) begin
            // read next char from input file
            case (encBytesRead % BUFFER_BYTES)
              0:  enctmp <= encBuf[encIdx][255:248];
              1:  enctmp <= encBuf[encIdx][247:240];
              2:  enctmp <= encBuf[encIdx][239:232];
              3:  enctmp <= encBuf[encIdx][231:224];
              4:  enctmp <= encBuf[encIdx][223:216];
              5:  enctmp <= encBuf[encIdx][215:208];
              6:  enctmp <= encBuf[encIdx][207:200];
              7:  enctmp <= encBuf[encIdx][199:192];
              8:  enctmp <= encBuf[encIdx][191:184];
              9:  enctmp <= encBuf[encIdx][183:176];
              10: enctmp <= encBuf[encIdx][175:168];
              11: enctmp <= encBuf[encIdx][167:160];
              12: enctmp <= encBuf[encIdx][159:152];
              13: enctmp <= encBuf[encIdx][151:144];
              14: enctmp <= encBuf[encIdx][143:136];
              15: enctmp <= encBuf[encIdx][135:128];
              16: enctmp <= encBuf[encIdx][127:120];
              17: enctmp <= encBuf[encIdx][119:112];
              18: enctmp <= encBuf[encIdx][111:104];
              19: enctmp <= encBuf[encIdx][103:96];
              20: enctmp <= encBuf[encIdx][95:88];
              21: enctmp <= encBuf[encIdx][87:80];
              22: enctmp <= encBuf[encIdx][79:72];
              23: enctmp <= encBuf[encIdx][71:64];
              24: enctmp <= encBuf[encIdx][63:56];
              25: enctmp <= encBuf[encIdx][55:48];
              26: enctmp <= encBuf[encIdx][47:40];
              27: enctmp <= encBuf[encIdx][39:32];
              28: enctmp <= encBuf[encIdx][31:24];
              29: enctmp <= encBuf[encIdx][23:16];
              30: enctmp <= encBuf[encIdx][15:8];
              31: enctmp <= encBuf[encIdx][7:0];
              default: $display("Unexpected value when filling in enctmp");

            endcase // case (encBytesRead % BUFFER_BYTES)

            encBytesRead <= encBytesRead + 1;

          end // if (eCtr == 1)

          if (eCtr == 2) begin
            // This only happens because encBytesRead 
            if ((encBytesRead % BUFFER_BYTES) == 0) begin
              $display("Reading more enc bytes");
              encIdx <= encIdx + 1;

              $display("encBuf[%d] = %h%h%h%h%h%h%h%h", encIdx + 1,
                   encBuf[encIdx][255:224],
                   encBuf[encIdx][223:192],
                   encBuf[encIdx][191:160],
                   encBuf[encIdx][159:128],
                   encBuf[encIdx][127:96],
                   encBuf[encIdx][95:64],
                   encBuf[encIdx][63:32],
                   encBuf[encIdx][31:0]);

            end

            // Prepare next state
            eCtr <= 0;
            encState <= ENC2;

          end // if (eCtr == 2)
        end // else: !if(encPcm != encExpVal)
        
      end // case: ENC3

      ENC4: begin
        encDone <= 1;

        eCtr <= 0;
        encState <= ENC0;

      end

      default: encState <= ENC0;

    endcase // case (encState)

  end // always @ (posedge clk)


  // decoder output checker - the decoder output is compared to the value read from
  // the ADPCM decoded samples file.
  always @(posedge clk) begin
    dCtr <= dCtr + 1;

    if (rst) decState <= DEC1;

    case (decState)
      DEC0: begin
        dCtr <= 0;
      end

      DEC1: begin
        // clear decoded sample value
        decCount <= 0;
        dispCount <= 0;

        decBytesRead <= 0;

        // "open" input file
        decIdx <= 0;

        // wait for reset release
        if (!rst) begin

          // decoder output compare loop
          dectmp <= decBuf[decIdx][(BUFFER_BYTES << 3) - 1:(BUFFER_BYTES << 3) - 8];
          decBytesRead <= decBytesRead + 1;
          
          $display("decBuf[%d] = %h%h%h%h%h%h%h%h", decIdx,
                   decBuf[decIdx][255:224],
                   decBuf[decIdx][223:192],
                   decBuf[decIdx][191:160],
                   decBuf[decIdx][159:128],
                   decBuf[decIdx][127:96],
                   decBuf[decIdx][95:64],
                   decBuf[decIdx][63:32],
                   decBuf[decIdx][31:0]);


          dCtr <= 0;
          decState <= DEC2;
        end
      end // case: DEC1

      DEC2: begin
        if (decBytesRead >= TOTAL_DEC_BYTES) begin
          $display("Reached eof of dec file");
          dCtr <= 0;
          decState <= DEC4;
        end

        else begin
          // read the next char to form the expected 16 bit sample value
          if (dCtr == 0) begin
            // display simulation progress bar title
            //$display("Simulation progress: ");
            
            decExpVal[7:0] <= dectmp;

            case (decBytesRead % BUFFER_BYTES)
              1:  decExpVal[15:8] <= decBuf[decIdx][247:240];
              3:  decExpVal[15:8] <= decBuf[decIdx][231:224];
              5:  decExpVal[15:8] <= decBuf[decIdx][215:208];
              7:  decExpVal[15:8] <= decBuf[decIdx][199:192];
              9:  decExpVal[15:8] <= decBuf[decIdx][183:176];
              11: decExpVal[15:8] <= decBuf[decIdx][167:160];
              13: decExpVal[15:8] <= decBuf[decIdx][151:144];
              15: decExpVal[15:8] <= decBuf[decIdx][135:128];
              17: decExpVal[15:8] <= decBuf[decIdx][119:112];
              19: decExpVal[15:8] <= decBuf[decIdx][103:96];
              21: decExpVal[15:8] <= decBuf[decIdx][87:80];
              23: decExpVal[15:8] <= decBuf[decIdx][71:64];
              25: decExpVal[15:8] <= decBuf[decIdx][55:48];
              27: decExpVal[15:8] <= decBuf[decIdx][39:32];
              29: decExpVal[15:8] <= decBuf[decIdx][23:16];
              31: decExpVal[15:8] <= decBuf[decIdx][7:0];
              default: $display("Unexpected number of bytes read for decExpVal");

            endcase // case (inBytesRead % BUFFER_BYTES)

            decBytesRead <= decBytesRead + 1;
          end // if (dCtr == 0)

          // This could be problematic bc what if decValid happens at dCtr 0?
          if (dCtr == 1) begin
            if ((decBytesRead % BUFFER_BYTES) == 0) begin
              decIdx <= decIdx + 1;

              $display("decBuf[%d] = %h%h%h%h%h%h%h%h", decIdx + 1,
                   decBuf[decIdx][255:224],
                   decBuf[decIdx][223:192],
                   decBuf[decIdx][191:160],
                   decBuf[decIdx][159:128],
                   decBuf[decIdx][127:96],
                   decBuf[decIdx][95:64],
                   decBuf[decIdx][63:32],
                   decBuf[decIdx][31:0]);
            end
          end

          // wait for decoder output valid
          if (decValid && dCtr >= 1) begin

            dCtr <= 0;
            decState <= DEC3;

          end
        end // else: !if($eof(decstream))

      end // case: DEC2

      DEC3: begin
        // compare the decoded value with the value read from the input file
        if (decSamp != decExpVal) begin
          if (dCtr == 0) begin
            // announce error detection and exit simulation
            $display(" Error!");
            $display("Error found in decoder output index %d.", decCount+1);
            $display("   (expected value 'h%h, got value 'h%h)", decExpVal, decSamp);
          end

          
          // wait for a few clock cycles before ending simulation
          if (dCtr >= 20) $finish();

        end // if (decSamp != decExpVal)

        else begin
          //$display("Dec correct! expected: %h, got: %h", decExpVal, decSamp);

          // delay for a clock cycle after comparison
          if (dCtr == 1) begin
            // update the decoded sample counter
            decCount <= decCount + 1;

            //// check if simulation progress should be displayed
            //if (dispCount[31:13] != (decCount >> 13))
            //  $write(".");
            // update the display counter
            //dispCount <= decCount;

            // read next char from input file
            case (decBytesRead % BUFFER_BYTES)
              0:  dectmp <= decBuf[decIdx][255:248];
              2:  dectmp <= decBuf[decIdx][239:232];
              4:  dectmp <= decBuf[decIdx][223:216];
              6:  dectmp <= decBuf[decIdx][207:200];
              8:  dectmp <= decBuf[decIdx][191:184];
              10: dectmp <= decBuf[decIdx][175:168];
              12: dectmp <= decBuf[decIdx][159:152];
              14: dectmp <= decBuf[decIdx][143:136];
              16: dectmp <= decBuf[decIdx][127:120];
              18: dectmp <= decBuf[decIdx][111:104];
              20: dectmp <= decBuf[decIdx][95:88];
              22: dectmp <= decBuf[decIdx][79:72];
              24: dectmp <= decBuf[decIdx][63:56];
              26: dectmp <= decBuf[decIdx][47:40];
              28: dectmp <= decBuf[decIdx][31:24];
              30: dectmp <= decBuf[decIdx][15:8];
              default: $display("Unexpected value");

            endcase // case (inBytesRead % BUFFER_BYTES)


            decBytesRead <= decBytesRead + 1;

          end // if (dCtr == 1)

          if (dCtr == 2) begin
            dCtr <= 0;
            decState <= DEC2;
          end // if (dCtr == 2)
        end // else: !if(decSamp != decExpVal)
      end // case: DEC3

      DEC4: begin
        // "close" input file

        // when decoder output is done announce simulation was successful
        $display(" Done");
        $display("Simulation ended successfully after %d samples", decCount);

        decDone <= 1;

        dCtr <= 0;
        decState <= 0;
      end // case: DEC4

      default: decState <= DEC0;

    endcase // case (decState)
  end // always @ (posedge clk)

/* */
  //------------------------------------------------------------------
  // device under test
  // Encoder instance


  ima_adpcm_enc enc
    (
     .clock(clk),
     .reset(rst),
     .inSamp(inSamp),
     .inValid(inValid),
     .inReady(inReady),
     .outPCM(encPcm),
     .outValid(encValid),
     .outPredictSamp(/* not used */),
     .outStepIndex(/* not used */)
     );



  // Decoder instance
  ima_adpcm_dec dec
    (
     .clock(clk),
     .reset(rst),
     .inPCM(encPcm),
     .inValid(encValid),
     .inReady(decReady),
     .inPredictSamp(16'b0),
     .inStepIndex(7'b0),
     .inStateLoad(1'b0),
     .outSamp(decSamp),
     .outValid(decValid)
     );

endmodule

test t(clock.val);
