module flushbuffer#( bytes )();
  parameter bytes = 2048;
  input wire[31:0] in_ld_bfr;


  output wire[31:0] out_ld_bfr;

  integer incnt;



endmodule
