module flushbuffer#(
  parameter BYTES = 2048
)(
  clk, 
  rst,
  N,
  in_valid,
  //in_incnt,
  in_bfr, 
  out_ld_bfr, 
  out_incnt,
  done
);
  localparam BITS = BYTES << 3;

  input wire clk;
  input wire rst;

  input wire [31:0] N;
  input wire in_valid;
  //input wire [31:0] in_incnt;
  input wire[BITS - 1:0] in_bfr;

  output reg[31:0] out_ld_bfr;
  output reg[31:0] out_incnt;
  output reg done;

  
  reg [31:0] ld_bfr;
  reg signed [31:0] incnt;
  integer bytes_read;
  reg loading_bfr;
  //reg [7:0] byte0, byte1, byte2, byte3;


  // Create byte array from input
  genvar i;
  for (i = 0; i < BYTES; i = i + 1) begin : BYTE
    wire [7:0] bi;

    assign bi = in_bfr[((BYTES - i) << 3) - 1:((BYTES - i) << 3) - 8];
    $display("BYTE[i].bi: %d", BYTE[i].bi);

  end
 
 
  always @(posedge clk) begin
    if (rst) begin
      $display("rst");
      ld_bfr <= 32'h4100000;
      incnt <= 32'b0;
      out_incnt <= 32'b0;
      done <= 1'b0;
      out_ld_bfr <= 0;  // TODO: something reasonable

      //temp_incnt <= 0;
      bytes_read <= 0;
      loading_bfr <= 1'b0;

      //byte0 <= 8'b0;
      //byte1 <= 8'b0;
      //byte2 <= 8'b0;
      //byte3 <= 8'b0;

    end
    else if (loading_bfr) begin
      $display("loading_bfr");
      if (incnt > 24) begin
        out_ld_bfr <= ld_bfr;
        out_incnt <= incnt;
        done <= 1'b1;
        loading_bfr <= 1'b0;

      end

      if (incnt <= 0) begin
        ld_bfr <= ld_bfr;
      end
      else if (incnt <= 8) begin
      end
           else if (incnt <= 16) begin
           end

                else if (incnt <= 24) begin
                end




    end
    else if (in_valid) begin // this should be last
      $display("starting new flush");

      // TODO: figure out how to mark inCnt as invalid
      // also deal with clock cycle delay between assigning incnt and getting incnt...
      $display("incnt: %d", incnt);
      ld_bfr <= (ld_bfr << (N % 32));
      incnt <= incnt - N;
      loading_bfr <= 1'b1;

      // TODO: deal with potential index out of bounds errors
      //byte0 <= in_bfr[(BYTES - bytes_read) - 1 : (BYTES - bytes_read) - 8];
      //byte1 <= in_bfr[(BYTES - bytes_read) - 9 : (BYTES - bytes_read) - 16];
      //byte2 <= in_bfr[(BYTES - bytes_read) - 17 : (BYTES - bytes_read) - 24];
      //byte2 <= in_bfr[(BYTES - bytes_read) - 25 : (BYTES - bytes_read) - 32];
      

    end

    //assign incnt = out_incnt - N;
    

  end

  


endmodule


// INITIALIZE FLUSH_BUFFER WITH IN_INCNT AS 0.
// in_incnt should be a reg that gets set to out_incnt from top module whenever
// flushbuffer = done
module test_flush_buf(input wire clk);

localparam in_bfr = {
  8'd0, 8'd104, 8'd120, 8'd48, 8'd72, 8'd32, 8'd160, 8'd192, 8'd192, 8'd64, 8'd56, 8'd248, 8'd248, 8'd88, 8'd136, 8'd224, 8'd200,
  8'd208, 8'd176, 8'd72, 8'd96, 8'd40, 8'd184, 8'd160, 8'd32, 8'd32, 8'd120, 8'd168, 8'd64, 8'd32, 8'd72, 8'd184,
  8'd216, 8'd240, 8'd0, 8'd216, 8'd192, 8'd64, 8'd112, 8'd48, 8'd160, 8'd152, 8'd40, 8'd176, 8'd32, 8'd32, 8'd248, 8'd200,
  8'd104, 8'd24, 8'd216, 8'd240, 8'd128, 8'd176, 8'd72, 8'd232, 8'd240, 8'd184, 8'd48, 8'd120, 8'd48, 8'd192, 8'd64, 8'd168,
  8'd160, 8'd128, 8'd160, 8'd160, 8'd232, 8'd208, 8'd104, 8'd120, 8'd232, 8'd120, 8'd8, 8'd184, 8'd120, 8'd200, 8'd64, 8'd160,
  8'd200, 8'd224, 8'd64, 8'd168, 8'd40, 8'd120, 8'd80, 8'd104, 8'd16, 8'd0, 8'd8, 8'd120, 8'd144, 8'd136, 8'd80, 8'd144,
  8'd72, 8'd24, 8'd128, 8'd216, 8'd216, 8'd24, 8'd80, 8'd16, 8'd64, 8'd32, 8'd200, 8'd112, 8'd128, 8'd144, 8'd88, 8'd24, 8'd112,
  8'd120, 8'd32, 8'd104, 8'd72, 8'd176, 8'd24, 8'd16, 8'd184, 8'd56, 8'd24, 8'd200, 8'd152, 8'd152, 8'd48, 8'd48,
  8'd136, 8'd80, 8'd240, 8'd8, 8'd216, 8'd200, 8'd240, 8'd32, 8'd168, 8'd112, 8'd48, 8'd56, 8'd40, 8'd192, 8'd232, 8'd32, 8'd48,
  8'd232, 8'd232, 8'd32, 8'd0, 8'd88, 8'd208, 8'd24, 8'd240, 8'd72, 8'd120, 8'd96, 8'd248, 8'd136, 8'd224, 8'd208,
  8'd8, 8'd184, 8'd192, 8'd144, 8'd88, 8'd48, 8'd144, 8'd136, 8'd112, 8'd192, 8'd96, 8'd240, 8'd200, 8'd160, 8'd184, 8'd160,
  8'd24, 8'd48, 8'd208, 8'd152, 8'd128, 8'd184, 8'd184, 8'd144, 8'd144, 8'd168, 8'd240, 8'd144, 8'd160, 8'd168, 8'd48,
  8'd48,
  8'd24, 8'd200, 8'd144, 8'd120, 8'd208, 8'd56, 8'd96, 8'd72, 8'd48, 8'd88, 8'd80, 8'd200, 8'd248, 8'd208, 8'd248, 8'd40, 8'd136,
  8'd112, 8'd32, 8'd8, 8'd8, 8'd80, 8'd192, 8'd40, 8'd32, 8'd224, 8'd56, 8'd192, 8'd200, 8'd56, 8'd56, 8'd232,
  8'd200, 8'd80, 8'd120, 8'd8, 8'd184, 8'd216, 8'd232, 8'd80, 8'd168, 8'd128, 8'd32, 8'd216, 8'd136, 8'd104, 8'd248, 8'd168,
  8'd248, 8'd8, 8'd192, 8'd168, 8'd192, 8'd56, 8'd240, 8'd192, 8'd208, 8'd136, 8'd120, 8'd48, 8'd224, 8'd112, 8'd168, 8'd80,
  8'd192, 8'd96, 8'd80, 8'd120, 8'd120, 8'd16, 8'd120, 8'd48, 8'd168, 8'd168, 8'd160, 8'd224, 8'd128, 8'd24, 8'd72, 8'd24,
  8'd248, 8'd240, 8'd152, 8'd160, 8'd208, 8'd56, 8'd192, 8'd56, 8'd88, 8'd128, 8'd192, 8'd136, 8'd128, 8'd208, 8'd112,
  8'd40,
  8'd64, 8'd192, 8'd32, 8'd176, 8'd80, 8'd56, 8'd168, 8'd208, 8'd24, 8'd168, 8'd168, 8'd248, 8'd240, 8'd136, 8'd96, 8'd32, 8'd56,
  8'd184, 8'd8, 8'd136, 8'd16, 8'd0, 8'd176, 8'd40, 8'd0, 8'd32, 8'd104, 8'd160, 8'd56, 8'd88, 8'd232, 8'd56,
  8'd0, 8'd240, 8'd184, 8'd232, 8'd88, 8'd32, 8'd176, 8'd0, 8'd216, 8'd248, 8'd184, 8'd40, 8'd16, 8'd80, 8'd8, 8'd208, 8'd64,
  8'd224, 8'd72, 8'd40, 8'd72, 8'd72, 8'd144, 8'd80, 8'd144, 8'd120, 8'd136, 8'd64, 8'd184, 8'd160, 8'd136, 8'd16,
  8'd48, 8'd104, 8'd232, 8'd104, 8'd104, 8'd72, 8'd208, 8'd72, 8'd192, 8'd184, 8'd40, 8'd56, 8'd232, 8'd72, 8'd160, 8'd80,
  8'd152, 8'd232, 8'd248, 8'd32, 8'd224, 8'd40, 8'd0, 8'd168, 8'd24, 8'd96, 8'd112, 8'd160, 8'd152, 8'd8, 8'd32, 8'd160,
  8'd104, 8'd208, 8'd32, 8'd24, 8'd248, 8'd8, 8'd248, 8'd144, 8'd120, 8'd16, 8'd192, 8'd88, 8'd152, 8'd176, 8'd200, 8'd160,
  8'd152, 8'd160, 8'd96, 8'd168, 8'd240, 8'd16, 8'd248, 8'd176, 8'd24, 8'd216, 8'd0, 8'd56, 8'd80, 8'd248, 8'd96, 8'd8,
  8'd128, 8'd32, 8'd192, 8'd104, 8'd48, 8'd208, 8'd240, 8'd184, 8'd128, 8'd80, 8'd56, 8'd192, 8'd0, 8'd112, 8'd176, 8'd48, 8'd96,
  8'd56, 8'd24, 8'd56, 8'd24, 8'd32, 8'd24, 8'd96, 8'd80, 8'd0, 8'd64, 8'd112, 8'd48, 8'd24, 8'd88, 8'd56,
  8'd152, 8'd224, 8'd160, 8'd192, 8'd184, 8'd72, 8'd248, 8'd128, 8'd8, 8'd8, 8'd104, 8'd104, 8'd200, 8'd48, 8'd136, 8'd136,
  8'd208, 8'd144, 8'd80, 8'd40, 8'd136, 8'd96, 8'd8, 8'd208, 8'd160, 8'd104, 8'd160, 8'd80, 8'd64, 8'd96, 8'd176, 8'd144,
  8'd8, 8'd56, 8'd88, 8'd88, 8'd208, 8'd120, 8'd48, 8'd240, 8'd240, 8'd96, 8'd248, 8'd192, 8'd104, 8'd128, 8'd248, 8'd24, 8'd104,
  8'd72, 8'd64, 8'd120, 8'd248, 8'd192, 8'd48, 8'd192, 8'd32, 8'd80, 8'd144, 8'd16, 8'd80, 8'd96, 8'd112, 8'd184,
  8'd56, 8'd80, 8'd248, 8'd232, 8'd0, 8'd40, 8'd248, 8'd56, 8'd192, 8'd32, 8'd192, 8'd96, 8'd248, 8'd48, 8'd136, 8'd224, 8'd80,
  8'd0, 8'd192, 8'd128, 8'd104, 8'd120, 8'd208, 8'd128, 8'd0, 8'd176, 8'd216, 8'd8, 8'd192, 8'd96, 8'd16, 8'd40,
  8'd184, 8'd96, 8'd32, 8'd72, 8'd80, 8'd192, 8'd104, 8'd104, 8'd136, 8'd0, 8'd16, 8'd160, 8'd24, 8'd104, 8'd48, 8'd8, 8'd24,
  8'd152, 8'd120, 8'd128, 8'd72, 8'd32, 8'd176, 8'd112, 8'd104, 8'd120, 8'd16, 8'd32, 8'd144, 8'd160, 8'd56, 8'd240,
  8'd0, 8'd232, 8'd184, 8'd24, 8'd16, 8'd208, 8'd200, 8'd240, 8'd200, 8'd200, 8'd104, 8'd112, 8'd24, 8'd208, 8'd128, 8'd168,
  8'd248, 8'd64, 8'd152, 8'd120, 8'd64, 8'd224, 8'd128, 8'd208, 8'd120, 8'd216, 8'd16, 8'd152, 8'd48, 8'd144, 8'd240, 8'd80,
  8'd144, 8'd224, 8'd48, 8'd160, 8'd192, 8'd248, 8'd0, 8'd128, 8'd120, 8'd128, 8'd160, 8'd232, 8'd168, 8'd208, 8'd112, 8'd112,
  8'd104, 8'd184, 8'd8, 8'd192, 8'd56, 8'd176, 8'd40, 8'd96, 8'd64, 8'd72, 8'd104, 8'd216, 8'd152, 8'd216, 8'd80, 8'd152,
  8'd184, 8'd216, 8'd32, 8'd56, 8'd32, 8'd64, 8'd240, 8'd152, 8'd240, 8'd168, 8'd136, 8'd8, 8'd232, 8'd168, 8'd128, 8'd88, 8'd72,
  8'd128, 8'd8, 8'd192, 8'd48, 8'd120, 8'd112, 8'd32, 8'd144, 8'd208, 8'd192, 8'd216, 8'd16, 8'd176, 8'd168, 8'd160,
  8'd168, 8'd88, 8'd136, 8'd56, 8'd8, 8'd64, 8'd0, 8'd80, 8'd216, 8'd104, 8'd64, 8'd80, 8'd88, 8'd208, 8'd64, 8'd80, 8'd200, 8'd24,
  8'd120, 8'd160, 8'd80, 8'd72, 8'd56, 8'd216, 8'd24, 8'd56, 8'd72, 8'd40, 8'd72, 8'd0, 8'd56, 8'd136,
  8'd56, 8'd200, 8'd72, 8'd136, 8'd88, 8'd72, 8'd136, 8'd240, 8'd0, 8'd176, 8'd176, 8'd152, 8'd192, 8'd248, 8'd224, 8'd240,
  8'd72, 8'd8, 8'd112, 8'd232, 8'd200, 8'd120, 8'd16, 8'd0, 8'd40, 8'd48, 8'd64, 8'd72, 8'd32, 8'd136, 8'd104, 8'd152,
  8'd16, 8'd240, 8'd184, 8'd80, 8'd0, 8'd152, 8'd32, 8'd176, 8'd128, 8'd120, 8'd0, 8'd160, 8'd40, 8'd64, 8'd112, 8'd40, 8'd80,
  8'd48, 8'd144, 8'd96, 8'd168, 8'd0, 8'd152, 8'd72, 8'd184, 8'd136, 8'd88, 8'd152, 8'd184, 8'd48, 8'd88, 8'd152,
  8'd96, 8'd216, 8'd240, 8'd184, 8'd200, 8'd136, 8'd64, 8'd104, 8'd112, 8'd232, 8'd0, 8'd208, 8'd176, 8'd128, 8'd112, 8'd248,
  8'd144, 8'd248, 8'd120, 8'd112, 8'd0, 8'd120, 8'd240, 8'd88, 8'd88, 8'd88, 8'd8, 8'd248, 8'd80, 8'd8, 8'd64, 8'd216,
  8'd240, 8'd56, 8'd56, 8'd144, 8'd112, 8'd208, 8'd144, 8'd72, 8'd16, 8'd160, 8'd136, 8'd216, 8'd176, 8'd112, 8'd56, 8'd8,
  8'd168, 8'd104, 8'd72, 8'd40, 8'd176, 8'd88, 8'd40, 8'd120, 8'd24, 8'd40, 8'd56, 8'd104, 8'd40, 8'd160, 8'd232, 8'd160,
  8'd24, 8'd144, 8'd144, 8'd232, 8'd120, 8'd144, 8'd112, 8'd96, 8'd136, 8'd176, 8'd8, 8'd128, 8'd112, 8'd184, 8'd96, 8'd120,
  8'd64, 8'd112, 8'd0, 8'd184, 8'd80, 8'd72, 8'd184, 8'd80, 8'd144, 8'd72, 8'd120, 8'd200, 8'd168, 8'd32, 8'd24, 8'd0,
  8'd144, 8'd72, 8'd24, 8'd248, 8'd24, 8'd152, 8'd72, 8'd128, 8'd0, 8'd8, 8'd224, 8'd32, 8'd72, 8'd72, 8'd48, 8'd112, 8'd232, 8'd16,
  8'd240, 8'd24, 8'd64, 8'd32, 8'd232, 8'd120, 8'd168, 8'd200, 8'd152, 8'd112, 8'd8, 8'd144, 8'd0, 8'd120,
  8'd112, 8'd0, 8'd112, 8'd144, 8'd72, 8'd160, 8'd24, 8'd216, 8'd112, 8'd128, 8'd224, 8'd152, 8'd104, 8'd136, 8'd40, 8'd0, 8'd16,
  8'd144, 8'd48, 8'd248, 8'd136, 8'd48, 8'd64, 8'd88, 8'd152, 8'd208, 8'd248, 8'd16, 8'd112, 8'd224, 8'd184, 8'd168,
  8'd40, 8'd168, 8'd64, 8'd248, 8'd144, 8'd104, 8'd200, 8'd144, 8'd152, 8'd16, 8'd168, 8'd192, 8'd240, 8'd96, 8'd72, 8'd136,
  8'd216, 8'd136, 8'd0, 8'd32, 8'd192, 8'd112, 8'd240, 8'd160, 8'd248, 8'd184, 8'd16, 8'd48, 8'd232, 8'd88, 8'd160, 8'd16,
  8'd104, 8'd176, 8'd144, 8'd136, 8'd24, 8'd240, 8'd184, 8'd160, 8'd8, 8'd16, 8'd32, 8'd56, 8'd176, 8'd144, 8'd168, 8'd168,
  8'd56, 8'd88, 8'd88, 8'd104, 8'd248, 8'd184, 8'd96, 8'd32, 8'd128, 8'd88, 8'd224, 8'd240, 8'd32, 8'd120, 8'd216, 8'd136,
  8'd8, 8'd72, 8'd80, 8'd104, 8'd120, 8'd152, 8'd32, 8'd96, 8'd232, 8'd80, 8'd232, 8'd24, 8'd80, 8'd200, 8'd208, 8'd216, 8'd184,
  8'd16, 8'd56, 8'd40, 8'd216, 8'd208, 8'd128, 8'd120, 8'd16, 8'd16, 8'd80, 8'd200, 8'd144, 8'd104, 8'd160, 8'd72,
  8'd24, 8'd136, 8'd176, 8'd32, 8'd192, 8'd120, 8'd136, 8'd80, 8'd16, 8'd88, 8'd208, 8'd160, 8'd16, 8'd232, 8'd40, 8'd24, 8'd144,
  8'd208, 8'd32, 8'd16, 8'd88, 8'd192, 8'd48, 8'd176, 8'd152, 8'd24, 8'd160, 8'd32, 8'd80, 8'd24, 8'd240, 8'd80,
  8'd160, 8'd152, 8'd160, 8'd128, 8'd80, 8'd88, 8'd40, 8'd184, 8'd208, 8'd144, 8'd48, 8'd200, 8'd200, 8'd48, 8'd112, 8'd144,
  8'd104, 8'd224, 8'd144, 8'd224, 8'd200, 8'd8, 8'd224, 8'd240, 8'd32, 8'd152, 8'd232, 8'd16, 8'd8, 8'd80, 8'd184, 8'd40,
  8'd184, 8'd248, 8'd64, 8'd8, 8'd232, 8'd16, 8'd88, 8'd88, 8'd8, 8'd120, 8'd128, 8'd48, 8'd240, 8'd88, 8'd64, 8'd104, 8'd104,
  8'd248, 8'd96, 8'd240, 8'd192, 8'd152, 8'd208, 8'd56, 8'd152, 8'd240, 8'd136, 8'd8, 8'd216, 8'd24, 8'd112, 8'd168,
  8'd88, 8'd136, 8'd80, 8'd224, 8'd136, 8'd152, 8'd40, 8'd24, 8'd248, 8'd216, 8'd152, 8'd136, 8'd96, 8'd224, 8'd64, 8'd80, 8'd56,
  8'd56, 8'd72, 8'd8, 8'd24, 8'd64, 8'd144, 8'd24, 8'd208, 8'd216, 8'd128, 8'd120, 8'd96, 8'd168, 8'd120, 8'd152,
  8'd112, 8'd232, 8'd136, 8'd80, 8'd72, 8'd96, 8'd152, 8'd208, 8'd72, 8'd216, 8'd64, 8'd120, 8'd120, 8'd48, 8'd232, 8'd72,
  8'd184, 8'd176, 8'd48, 8'd232, 8'd200, 8'd184, 8'd120, 8'd72, 8'd112, 8'd128, 8'd248, 8'd160, 8'd168, 8'd216, 8'd152,
  8'd80,
  8'd176, 8'd112, 8'd48, 8'd152, 8'd112, 8'd64, 8'd40, 8'd200, 8'd232, 8'd80, 8'd160, 8'd56, 8'd216, 8'd192, 8'd168, 8'd72,
  8'd40, 8'd64, 8'd208, 8'd32, 8'd224, 8'd240, 8'd24, 8'd104, 8'd232, 8'd240, 8'd168, 8'd24, 8'd248, 8'd32, 8'd80, 8'd152,
  8'd144, 8'd160, 8'd112, 8'd120, 8'd96, 8'd240, 8'd64, 8'd160, 8'd248, 8'd248, 8'd152, 8'd48, 8'd112, 8'd88, 8'd128, 8'd232,
  8'd240, 8'd240, 8'd232, 8'd168, 8'd120, 8'd32, 8'd152, 8'd176, 8'd104, 8'd16, 8'd80, 8'd152, 8'd240, 8'd224, 8'd128,
  8'd16,
  8'd48, 8'd32, 8'd216, 8'd8, 8'd104, 8'd248, 8'd184, 8'd208, 8'd216, 8'd120, 8'd80, 8'd208, 8'd128, 8'd56, 8'd112, 8'd40,
  8'd184, 8'd16, 8'd224, 8'd168, 8'd152, 8'd248, 8'd56, 8'd144, 8'd168, 8'd224, 8'd8, 8'd168, 8'd80, 8'd136, 8'd152, 8'd48,
  8'd96, 8'd0, 8'd184, 8'd88, 8'd192, 8'd24, 8'd16, 8'd128, 8'd0, 8'd176, 8'd152, 8'd40, 8'd96, 8'd72, 8'd192, 8'd0, 8'd32, 8'd128,
  8'd24, 8'd240, 8'd48, 8'd248, 8'd176, 8'd120, 8'd16, 8'd168, 8'd224, 8'd72, 8'd8, 8'd200, 8'd48, 8'd176,
  8'd112, 8'd224, 8'd160, 8'd8, 8'd152, 8'd64, 8'd16, 8'd16, 8'd240, 8'd224, 8'd64, 8'd144, 8'd128, 8'd80, 8'd184, 8'd40, 8'd232,
  8'd200, 8'd112, 8'd248, 8'd24, 8'd112, 8'd176, 8'd128, 8'd128, 8'd56, 8'd40, 8'd152, 8'd24, 8'd184, 8'd120, 8'd104,
  8'd72, 8'd64, 8'd200, 8'd48, 8'd224, 8'd0, 8'd56, 8'd232, 8'd32, 8'd240, 8'd184, 8'd104, 8'd104, 8'd32, 8'd192, 8'd200, 8'd200,
  8'd64, 8'd152, 8'd72, 8'd216, 8'd216, 8'd80, 8'd0, 8'd80, 8'd0, 8'd0, 8'd160, 8'd120, 8'd40, 8'd136, 8'd240,
  8'd32, 8'd120, 8'd152, 8'd216, 8'd56, 8'd112, 8'd16, 8'd24, 8'd8, 8'd120, 8'd104, 8'd192, 8'd144, 8'd176, 8'd8, 8'd16, 8'd96,
  8'd104, 8'd168, 8'd80, 8'd192, 8'd232, 8'd112, 8'd112, 8'd56, 8'd88, 8'd176, 8'd240, 8'd32, 8'd176, 8'd248, 8'd80,
  8'd176, 8'd24, 8'd224, 8'd192, 8'd8, 8'd176, 8'd168, 8'd16, 8'd232, 8'd248, 8'd16, 8'd16, 8'd104, 8'd128, 8'd232, 8'd0, 8'd32,
  8'd240, 8'd112, 8'd32, 8'd184, 8'd184, 8'd56, 8'd232, 8'd80, 8'd144, 8'd16, 8'd72, 8'd240, 8'd208, 8'd64, 8'd176,
  8'd240, 8'd16, 8'd136, 8'd16, 8'd80, 8'd192, 8'd24, 8'd72, 8'd216, 8'd56, 8'd80, 8'd216, 8'd32, 8'd144, 8'd72, 8'd24, 8'd64,
  8'd248, 8'd0, 8'd224, 8'd72, 8'd32, 8'd136, 8'd232, 8'd240, 8'd72, 8'd32, 8'd88, 8'd128, 8'd104, 8'd16, 8'd8,
  8'd32, 8'd192, 8'd224, 8'd8, 8'd152, 8'd248, 8'd224, 8'd0, 8'd176, 8'd48, 8'd16, 8'd104, 8'd216, 8'd176, 8'd24, 8'd240, 8'd200,
  8'd80, 8'd248, 8'd208, 8'd128, 8'd200, 8'd72, 8'd8, 8'd152, 8'd128, 8'd80, 8'd120, 8'd80, 8'd152, 8'd232, 8'd200,
  8'd168, 8'd88, 8'd16, 8'd176, 8'd232, 8'd40, 8'd72, 8'd208, 8'd232, 8'd112, 8'd240, 8'd112, 8'd80, 8'd176, 8'd176, 8'd16,
  8'd72, 8'd120, 8'd32, 8'd184, 8'd224, 8'd80, 8'd24, 8'd176, 8'd0, 8'd208, 8'd16, 8'd56, 8'd112, 8'd16, 8'd120, 8'd160,
  8'd24, 8'd216, 8'd128, 8'd136, 8'd192, 8'd152, 8'd248, 8'd120, 8'd160, 8'd56, 8'd192, 8'd224, 8'd0, 8'd136, 8'd112, 8'd112,
  8'd8, 8'd8, 8'd184, 8'd168, 8'd88, 8'd160, 8'd120, 8'd160, 8'd240, 8'd168, 8'd32, 8'd40, 8'd168, 8'd88, 8'd8, 8'd16,
  8'd24, 8'd104, 8'd104, 8'd48, 8'd248, 8'd136, 8'd72, 8'd144, 8'd128, 8'd160, 8'd216, 8'd88, 8'd240, 8'd120, 8'd232, 8'd72,
  8'd192, 8'd200, 8'd248, 8'd192, 8'd48, 8'd240, 8'd104, 8'd208, 8'd40, 8'd104, 8'd16, 8'd128, 8'd80, 8'd224, 8'd224, 8'd56,
  8'd56, 8'd120, 8'd40, 8'd24, 8'd176, 8'd16, 8'd184, 8'd24, 8'd176, 8'd224, 8'd168, 8'd16, 8'd184, 8'd104, 8'd136, 8'd200,
  8'd168, 8'd208, 8'd120, 8'd200, 8'd224, 8'd40, 8'd208, 8'd16, 8'd112, 8'd160, 8'd192, 8'd224, 8'd64, 8'd40, 8'd232,
  8'd120,
  8'd24, 8'd232, 8'd168, 8'd80, 8'd88, 8'd144, 8'd104, 8'd72, 8'd192, 8'd112, 8'd0, 8'd112, 8'd104, 8'd224, 8'd232, 8'd160,
  8'd112, 8'd208, 8'd176, 8'd216, 8'd56, 8'd224, 8'd224, 8'd160, 8'd104, 8'd56, 8'd176, 8'd216, 8'd192, 8'd24, 8'd208, 8'd8,
  8'd40, 8'd56, 8'd248, 8'd8, 8'd120, 8'd184, 8'd128, 8'd40, 8'd168, 8'd56, 8'd184, 8'd192, 8'd136, 8'd96, 8'd72, 8'd216, 8'd8,
  8'd64, 8'd72, 8'd56, 8'd16, 8'd176, 8'd144, 8'd16, 8'd128, 8'd176, 8'd136, 8'd208, 8'd120, 8'd16, 8'd184, 8'd224,
  8'd160, 8'd216, 8'd144, 8'd88, 8'd208, 8'd200, 8'd144, 8'd96, 8'd152, 8'd200, 8'd224, 8'd208, 8'd240, 8'd120, 8'd8, 8'd104,
  8'd184, 8'd112, 8'd168, 8'd200, 8'd112, 8'd72, 8'd0, 8'd192, 8'd0, 8'd40, 8'd120, 8'd136, 8'd112, 8'd40, 8'd152, 8'd56,
  8'd144, 8'd32, 8'd224, 8'd240, 8'd32, 8'd192, 8'd56, 8'd200, 8'd16, 8'd136, 8'd104, 8'd192, 8'd192, 8'd0, 8'd0, 8'd0, 8'd8,
  8'd232, 8'd104, 8'd240, 8'd88, 8'd192, 8'd8, 8'd168, 8'd216, 8'd208, 8'd184, 8'd224, 8'd240, 8'd72, 8'd152, 8'd72,
  8'd168, 8'd184, 8'd176, 8'd216, 8'd48, 8'd144, 8'd80, 8'd32, 8'd184, 8'd208, 8'd112, 8'd160, 8'd88, 8'd88, 8'd8, 8'd144,
  8'd144, 8'd120, 8'd152, 8'd48, 8'd200, 8'd168, 8'd112, 8'd8, 8'd160, 8'd216, 8'd240, 8'd128, 8'd104, 8'd128, 8'd144,
  8'd248,
  8'd64, 8'd168, 8'd136, 8'd240, 8'd160, 8'd56, 8'd136, 8'd216, 8'd80, 8'd56, 8'd192, 8'd32, 8'd64, 8'd128, 8'd80, 8'd32, 8'd32,
  8'd96, 8'd88, 8'd200, 8'd152, 8'd72, 8'd160, 8'd16, 8'd128, 8'd200, 8'd160, 8'd144, 8'd112, 8'd16, 8'd112, 8'd152,
  8'd56, 8'd136, 8'd56, 8'd216, 8'd8, 8'd24, 8'd192, 8'd144, 8'd176, 8'd200, 8'd48, 8'd72, 8'd40, 8'd72, 8'd240, 8'd120, 8'd120,
  8'd160, 8'd80, 8'd152, 8'd144, 8'd216, 8'd224, 8'd152, 8'd40, 8'd144, 8'd160, 8'd88, 8'd184, 8'd184, 8'd192, 8'd128,
  8'd0, 8'd200, 8'd72, 8'd112, 8'd208, 8'd248, 8'd152, 8'd0, 8'd152, 8'd8, 8'd40, 8'd16, 8'd168, 8'd152, 8'd64, 8'd176, 8'd88,
  8'd24, 8'd232, 8'd136, 8'd32, 8'd152, 8'd232, 8'd208, 8'd192, 8'd240, 8'd136, 8'd0, 8'd232, 8'd200, 8'd8, 8'd216,
  8'd104, 8'd184, 8'd64, 8'd192, 8'd8, 8'd96, 8'd184, 8'd120, 8'd208, 8'd80, 8'd16, 8'd64, 8'd136, 8'd136, 8'd72, 8'd8, 8'd112,
  8'd184, 8'd248, 8'd120, 8'd136, 8'd8, 8'd56, 8'd232, 8'd208, 8'd96, 8'd16, 8'd64, 8'd168, 8'd112, 8'd48, 8'd32,
  8'd184, 8'd224, 8'd72, 8'd88, 8'd128, 8'd184, 8'd72, 8'd168, 8'd224, 8'd216, 8'd160, 8'd232, 8'd64, 8'd168, 8'd48, 8'd152,
  8'd64, 8'd152, 8'd16, 8'd200, 8'd168, 8'd56, 8'd144, 8'd192, 8'd64, 8'd120, 8'd168, 8'd8, 8'd128, 8'd216, 8'd16, 8'd8,
  8'd104, 8'd32, 8'd128, 8'd96, 8'd160, 8'd88, 8'd136, 8'd96, 8'd56, 8'd16, 8'd128, 8'd56, 8'd88, 8'd16, 8'd208, 8'd200, 8'd24,
  8'd96, 8'd240, 8'd32, 8'd232, 8'd192, 8'd104, 8'd168, 8'd40, 8'd0, 8'd192, 8'd40, 8'd200, 8'd96, 8'd184, 8'd8,
  8'd72, 8'd216, 8'd104, 8'd232, 8'd112, 8'd248, 8'd8, 8'd8, 8'd248, 8'd192, 8'd152, 8'd32, 8'd0, 8'd168, 8'd232, 8'd80, 8'd248,
  8'd64, 8'd8, 8'd24, 8'd80, 8'd32, 8'd96, 8'd240, 8'd232, 8'd48, 8'd80, 8'd16, 8'd144, 8'd200, 8'd16, 8'd48,
  8'd88, 8'd40, 8'd112, 8'd232, 8'd88, 8'd168, 8'd56, 8'd160, 8'd232, 8'd16, 8'd128, 8'd248, 8'd48, 8'd80, 8'd200, 8'd168,
  8'd152, 8'd72, 8'd216, 8'd224, 8'd72, 8'd208, 8'd152, 8'd192, 8'd0, 8'd224, 8'd48, 8'd136, 8'd168, 8'd96, 8'd16, 8'd152
};

const unsigned char out_ld_Rdptr[Num] = {
  8'72, 8'd184, 8'd216, 8'd240, 8'd0, 8'd216, 8'd192, 8'd64, 8'd112, 8'd48, 8'd160, 8'd152, 8'd40, 8'd176, 8'd32, 8'd32, 8'd248,
  8'd200, 8'd104, 8'd24, 8'd216, 8'd240, 8'd128, 8'd176, 8'd72, 8'd232, 8'd240, 8'd184, 8'd48, 8'd120, 8'd48, 8'd192,
  8'd64, 8'd168, 8'd160, 8'd128, 8'd160, 8'd160, 8'd232, 8'd208, 8'd104, 8'd120, 8'd232, 8'd120, 8'd8, 8'd184, 8'd120, 8'd200,
  8'd64, 8'd160, 8'd200, 8'd224, 8'd64, 8'd168, 8'd40, 8'd120, 8'd80, 8'd104, 8'd16, 8'd0, 8'd8, 8'd120, 8'd144, 8'd136,
  8'd80, 8'd144, 8'd72, 8'd24, 8'd128, 8'd216, 8'd216, 8'd24, 8'd80, 8'd16, 8'd64, 8'd32, 8'd200, 8'd112, 8'd128, 8'd144, 8'd88,
  8'd24, 8'd112, 8'd120, 8'd32, 8'd104, 8'd72, 8'd176, 8'd24, 8'd16, 8'd184, 8'd56, 8'd24, 8'd200, 8'd152, 8'd152,
  8'd48, 8'd48, 8'd136, 8'd80, 8'd240, 8'd8, 8'd216, 8'd200, 8'd240, 8'd32, 8'd168, 8'd112, 8'd48, 8'd56, 8'd40, 8'd192, 8'd232,
  8'd32, 8'd48, 8'd232, 8'd232, 8'd32, 8'd0, 8'd88, 8'd208, 8'd24, 8'd240, 8'd72, 8'd120, 8'd96, 8'd248, 8'd136,
  8'd224, 8'd208, 8'd8, 8'd184, 8'd192, 8'd144, 8'd88, 8'd48, 8'd144, 8'd136, 8'd112, 8'd192, 8'd96, 8'd240, 8'd200, 8'd160,
  8'd184, 8'd160, 8'd24, 8'd48, 8'd208, 8'd152, 8'd128, 8'd184, 8'd184, 8'd144, 8'd144, 8'd168, 8'd240, 8'd144, 8'd160,
  8'd168,
  8'd48, 8'd48, 8'd24, 8'd200, 8'd144, 8'd120, 8'd208, 8'd56, 8'd96, 8'd72, 8'd48, 8'd88, 8'd80, 8'd200, 8'd248, 8'd208, 8'd248,
  8'd40, 8'd136, 8'd112, 8'd32, 8'd8, 8'd8, 8'd80, 8'd192, 8'd40, 8'd32, 8'd224, 8'd56, 8'd192, 8'd200, 8'd56,
  8'd56, 8'd232, 8'd200, 8'd80, 8'd120, 8'd8, 8'd184, 8'd216, 8'd232, 8'd80, 8'd168, 8'd128, 8'd32, 8'd216, 8'd136, 8'd104,
  8'd248, 8'd168, 8'd248, 8'd8, 8'd192, 8'd168, 8'd192, 8'd56, 8'd240, 8'd192, 8'd208, 8'd136, 8'd120, 8'd48, 8'd224,
  8'd112,
  8'd168, 8'd80, 8'd192, 8'd96, 8'd80, 8'd120, 8'd120, 8'd16, 8'd120, 8'd48, 8'd168, 8'd168, 8'd160, 8'd224, 8'd128, 8'd24,
  8'd72, 8'd24, 8'd248, 8'd240, 8'd152, 8'd160, 8'd208, 8'd56, 8'd192, 8'd56, 8'd88, 8'd128, 8'd192, 8'd136, 8'd128, 8'd208,
  8'd112, 8'd40, 8'd64, 8'd192, 8'd32, 8'd176, 8'd80, 8'd56, 8'd168, 8'd208, 8'd24, 8'd168, 8'd168, 8'd248, 8'd240, 8'd136,
  8'd96, 8'd32, 8'd56, 8'd184, 8'd8, 8'd136, 8'd16, 8'd0, 8'd176, 8'd40, 8'd0, 8'd32, 8'd104, 8'd160, 8'd56, 8'd88,
  8'd232, 8'd56, 8'd0, 8'd240, 8'd184, 8'd232, 8'd88, 8'd32, 8'd176, 8'd0, 8'd216, 8'd248, 8'd184, 8'd40, 8'd16, 8'd80, 8'd8,
  8'd208, 8'd64, 8'd224, 8'd72, 8'd40, 8'd72, 8'd72, 8'd144, 8'd80, 8'd144, 8'd120, 8'd136, 8'd64, 8'd184, 8'd160,
  8'd136, 8'd16, 8'd48, 8'd104, 8'd232, 8'd104, 8'd104, 8'd72, 8'd208, 8'd72, 8'd192, 8'd184, 8'd40, 8'd56, 8'd232, 8'd72,
  8'd160, 8'd80, 8'd152, 8'd232, 8'd248, 8'd32, 8'd224, 8'd40, 8'd0, 8'd168, 8'd24, 8'd96, 8'd112, 8'd160, 8'd152, 8'd8,
  8'd32, 8'd160, 8'd104, 8'd208, 8'd32, 8'd24, 8'd248, 8'd8, 8'd248, 8'd144, 8'd120, 8'd16, 8'd192, 8'd88, 8'd152, 8'd176,
  8'd200, 8'd160, 8'd152, 8'd160, 8'd96, 8'd168, 8'd240, 8'd16, 8'd248, 8'd176, 8'd24, 8'd216, 8'd0, 8'd56, 8'd80, 8'd248,
  8'd96, 8'd8, 8'd128, 8'd32, 8'd192, 8'd104, 8'd48, 8'd208, 8'd240, 8'd184, 8'd128, 8'd80, 8'd56, 8'd192, 8'd0, 8'd112, 8'd176,
  8'd48, 8'd96, 8'd56, 8'd24, 8'd56, 8'd24, 8'd32, 8'd24, 8'd96, 8'd80, 8'd0, 8'd64, 8'd112, 8'd48, 8'd24,
  8'd88, 8'd56, 8'd152, 8'd224, 8'd160, 8'd192, 8'd184, 8'd72, 8'd248, 8'd128, 8'd8, 8'd8, 8'd104, 8'd104, 8'd200, 8'd48, 8'd136,
  8'd136, 8'd208, 8'd144, 8'd80, 8'd40, 8'd136, 8'd96, 8'd8, 8'd208, 8'd160, 8'd104, 8'd160, 8'd80, 8'd64, 8'd96,
  8'd176, 8'd144, 8'd8, 8'd56, 8'd88, 8'd88, 8'd208, 8'd120, 8'd48, 8'd240, 8'd240, 8'd96, 8'd248, 8'd192, 8'd104, 8'd128,
  8'd248, 8'd24, 8'd104, 8'd72, 8'd64, 8'd120, 8'd248, 8'd192, 8'd48, 8'd192, 8'd32, 8'd80, 8'd144, 8'd16, 8'd80, 8'd96,
  8'd112, 8'd184, 8'd56, 8'd80, 8'd248, 8'd232, 8'd0, 8'd40, 8'd248, 8'd56, 8'd192, 8'd32, 8'd192, 8'd96, 8'd248, 8'd48, 8'd136,
  8'd224, 8'd80, 8'd0, 8'd192, 8'd128, 8'd104, 8'd120, 8'd208, 8'd128, 8'd0, 8'd176, 8'd216, 8'd8, 8'd192, 8'd96,
  8'd16, 8'd40, 8'd184, 8'd96, 8'd32, 8'd72, 8'd80, 8'd192, 8'd104, 8'd104, 8'd136, 8'd0, 8'd16, 8'd160, 8'd24, 8'd104, 8'd48, 8'd8,
  8'd24, 8'd152, 8'd120, 8'd128, 8'd72, 8'd32, 8'd176, 8'd112, 8'd104, 8'd120, 8'd16, 8'd32, 8'd144, 8'd160,
  8'd56, 8'd240, 8'd0, 8'd232, 8'd184, 8'd24, 8'd16, 8'd208, 8'd200, 8'd240, 8'd200, 8'd200, 8'd104, 8'd112, 8'd24, 8'd208,
  8'd128, 8'd168, 8'd248, 8'd64, 8'd152, 8'd120, 8'd64, 8'd224, 8'd128, 8'd208, 8'd120, 8'd216, 8'd16, 8'd152, 8'd48,
  8'd144,
  8'd240, 8'd80, 8'd144, 8'd224, 8'd48, 8'd160, 8'd192, 8'd248, 8'd0, 8'd128, 8'd120, 8'd128, 8'd160, 8'd232, 8'd168, 8'd208,
  8'd112, 8'd112, 8'd104, 8'd184, 8'd8, 8'd192, 8'd56, 8'd176, 8'd40, 8'd96, 8'd64, 8'd72, 8'd104, 8'd216, 8'd152, 8'd216,
  8'd80, 8'd152, 8'd184, 8'd216, 8'd32, 8'd56, 8'd32, 8'd64, 8'd240, 8'd152, 8'd240, 8'd168, 8'd136, 8'd8, 8'd232, 8'd168,
  8'd128, 8'd88, 8'd72, 8'd128, 8'd8, 8'd192, 8'd48, 8'd120, 8'd112, 8'd32, 8'd144, 8'd208, 8'd192, 8'd216, 8'd16, 8'd176,
  8'd168, 8'd160, 8'd168, 8'd88, 8'd136, 8'd56, 8'd8, 8'd64, 8'd0, 8'd80, 8'd216, 8'd104, 8'd64, 8'd80, 8'd88, 8'd208, 8'd64, 8'd80,
  8'd200, 8'd24, 8'd120, 8'd160, 8'd80, 8'd72, 8'd56, 8'd216, 8'd24, 8'd56, 8'd72, 8'd40, 8'd72, 8'd0,
  8'd56, 8'd136, 8'd56, 8'd200, 8'd72, 8'd136, 8'd88, 8'd72, 8'd136, 8'd240, 8'd0, 8'd176, 8'd176, 8'd152, 8'd192, 8'd248,
  8'd224, 8'd240, 8'd72, 8'd8, 8'd112, 8'd232, 8'd200, 8'd120, 8'd16, 8'd0, 8'd40, 8'd48, 8'd64, 8'd72, 8'd32, 8'd136,
  8'd104, 8'd152, 8'd16, 8'd240, 8'd184, 8'd80, 8'd0, 8'd152, 8'd32, 8'd176, 8'd128, 8'd120, 8'd0, 8'd160, 8'd40, 8'd64, 8'd112,
  8'd40, 8'd80, 8'd48, 8'd144, 8'd96, 8'd168, 8'd0, 8'd152, 8'd72, 8'd184, 8'd136, 8'd88, 8'd152, 8'd184, 8'd48,
  8'd88, 8'd152, 8'd96, 8'd216, 8'd240, 8'd184, 8'd200, 8'd136, 8'd64, 8'd104, 8'd112, 8'd232, 8'd0, 8'd208, 8'd176, 8'd128,
  8'd112, 8'd248, 8'd144, 8'd248, 8'd120, 8'd112, 8'd0, 8'd120, 8'd240, 8'd88, 8'd88, 8'd88, 8'd8, 8'd248, 8'd80, 8'd8,
  8'd64, 8'd216, 8'd240, 8'd56, 8'd56, 8'd144, 8'd112, 8'd208, 8'd144, 8'd72, 8'd16, 8'd160, 8'd136, 8'd216, 8'd176, 8'd112,
  8'd56, 8'd8, 8'd168, 8'd104, 8'd72, 8'd40, 8'd176, 8'd88, 8'd40, 8'd120, 8'd24, 8'd40, 8'd56, 8'd104, 8'd40, 8'd160,
  8'd232, 8'd160, 8'd24, 8'd144, 8'd144, 8'd232, 8'd120, 8'd144, 8'd112, 8'd96, 8'd136, 8'd176, 8'd8, 8'd128, 8'd112, 8'd184,
  8'd96, 8'd120, 8'd64, 8'd112, 8'd0, 8'd184, 8'd80, 8'd72, 8'd184, 8'd80, 8'd144, 8'd72, 8'd120, 8'd200, 8'd168, 8'd32,
  8'd24, 8'd0, 8'd144, 8'd72, 8'd24, 8'd248, 8'd24, 8'd152, 8'd72, 8'd128, 8'd0, 8'd8, 8'd224, 8'd32, 8'd72, 8'd72, 8'd48, 8'd112,
  8'd232, 8'd16, 8'd240, 8'd24, 8'd64, 8'd32, 8'd232, 8'd120, 8'd168, 8'd200, 8'd152, 8'd112, 8'd8, 8'd144,
  8'd0, 8'd120, 8'd112, 8'd0, 8'd112, 8'd144, 8'd72, 8'd160, 8'd24, 8'd216, 8'd112, 8'd128, 8'd224, 8'd152, 8'd104, 8'd136,
  8'd40, 8'd0, 8'd16, 8'd144, 8'd48, 8'd248, 8'd136, 8'd48, 8'd64, 8'd88, 8'd152, 8'd208, 8'd248, 8'd16, 8'd112, 8'd224,
  8'd184, 8'd168, 8'd40, 8'd168, 8'd64, 8'd248, 8'd144, 8'd104, 8'd200, 8'd144, 8'd152, 8'd16, 8'd168, 8'd192, 8'd240, 8'd96,
  8'd72, 8'd136, 8'd216, 8'd136, 8'd0, 8'd32, 8'd192, 8'd112, 8'd240, 8'd160, 8'd248, 8'd184, 8'd16, 8'd48, 8'd232, 8'd88,
  8'd160, 8'd16, 8'd104, 8'd176, 8'd144, 8'd136, 8'd24, 8'd240, 8'd184, 8'd160, 8'd8, 8'd16, 8'd32, 8'd56, 8'd176, 8'd144,
  8'd168, 8'd168, 8'd56, 8'd88, 8'd88, 8'd104, 8'd248, 8'd184, 8'd96, 8'd32, 8'd128, 8'd88, 8'd224, 8'd240, 8'd32, 8'd120,
  8'd216, 8'd136, 8'd8, 8'd72, 8'd80, 8'd104, 8'd120, 8'd152, 8'd32, 8'd96, 8'd232, 8'd80, 8'd232, 8'd24, 8'd80, 8'd200, 8'd208,
  8'd216, 8'd184, 8'd16, 8'd56, 8'd40, 8'd216, 8'd208, 8'd128, 8'd120, 8'd16, 8'd16, 8'd80, 8'd200, 8'd144, 8'd104,
  8'd160, 8'd72, 8'd24, 8'd136, 8'd176, 8'd32, 8'd192, 8'd120, 8'd136, 8'd80, 8'd16, 8'd88, 8'd208, 8'd160, 8'd16, 8'd232, 8'd40,
  8'd24, 8'd144, 8'd208, 8'd32, 8'd16, 8'd88, 8'd192, 8'd48, 8'd176, 8'd152, 8'd24, 8'd160, 8'd32, 8'd80, 8'd24,
  8'd240, 8'd80, 8'd160, 8'd152, 8'd160, 8'd128, 8'd80, 8'd88, 8'd40, 8'd184, 8'd208, 8'd144, 8'd48, 8'd200, 8'd200, 8'd48,
  8'd112, 8'd144, 8'd104, 8'd224, 8'd144, 8'd224, 8'd200, 8'd8, 8'd224, 8'd240, 8'd32, 8'd152, 8'd232, 8'd16, 8'd8, 8'd80,
  8'd184, 8'd40, 8'd184, 8'd248, 8'd64, 8'd8, 8'd232, 8'd16, 8'd88, 8'd88, 8'd8, 8'd120, 8'd128, 8'd48, 8'd240, 8'd88, 8'd64,
  8'd104, 8'd104, 8'd248, 8'd96, 8'd240, 8'd192, 8'd152, 8'd208, 8'd56, 8'd152, 8'd240, 8'd136, 8'd8, 8'd216, 8'd24,
  8'd112, 8'd168, 8'd88, 8'd136, 8'd80, 8'd224, 8'd136, 8'd152, 8'd40, 8'd24, 8'd248, 8'd216, 8'd152, 8'd136, 8'd96, 8'd224,
  8'd64, 8'd80, 8'd56, 8'd56, 8'd72, 8'd8, 8'd24, 8'd64, 8'd144, 8'd24, 8'd208, 8'd216, 8'd128, 8'd120, 8'd96, 8'd168,
  8'd120, 8'd152, 8'd112, 8'd232, 8'd136, 8'd80, 8'd72, 8'd96, 8'd152, 8'd208, 8'd72, 8'd216, 8'd64, 8'd120, 8'd120, 8'd48,
  8'd232, 8'd72, 8'd184, 8'd176, 8'd48, 8'd232, 8'd200, 8'd184, 8'd120, 8'd72, 8'd112, 8'd128, 8'd248, 8'd160, 8'd168,
  8'd216,
  8'd152, 8'd80, 8'd176, 8'd112, 8'd48, 8'd152, 8'd112, 8'd64, 8'd40, 8'd200, 8'd232, 8'd80, 8'd160, 8'd56, 8'd216, 8'd192,
  8'd168, 8'd72, 8'd40, 8'd64, 8'd208, 8'd32, 8'd224, 8'd240, 8'd24, 8'd104, 8'd232, 8'd240, 8'd168, 8'd24, 8'd248, 8'd32,
  8'd80, 8'd152, 8'd144, 8'd160, 8'd112, 8'd120, 8'd96, 8'd240, 8'd64, 8'd160, 8'd248, 8'd248, 8'd152, 8'd48, 8'd112, 8'd88,
  8'd128, 8'd232, 8'd240, 8'd240, 8'd232, 8'd168, 8'd120, 8'd32, 8'd152, 8'd176, 8'd104, 8'd16, 8'd80, 8'd152, 8'd240,
  8'd224,
  8'd128, 8'd16, 8'd48, 8'd32, 8'd216, 8'd8, 8'd104, 8'd248, 8'd184, 8'd208, 8'd216, 8'd120, 8'd80, 8'd208, 8'd128, 8'd56,
  8'd112, 8'd40, 8'd184, 8'd16, 8'd224, 8'd168, 8'd152, 8'd248, 8'd56, 8'd144, 8'd168, 8'd224, 8'd8, 8'd168, 8'd80, 8'd136,
  8'd152, 8'd48, 8'd96, 8'd0, 8'd184, 8'd88, 8'd192, 8'd24, 8'd16, 8'd128, 8'd0, 8'd176, 8'd152, 8'd40, 8'd96, 8'd72, 8'd192, 8'd0,
  8'd32, 8'd128, 8'd24, 8'd240, 8'd48, 8'd248, 8'd176, 8'd120, 8'd16, 8'd168, 8'd224, 8'd72, 8'd8, 8'd200,
  8'd48, 8'd176, 8'd112, 8'd224, 8'd160, 8'd8, 8'd152, 8'd64, 8'd16, 8'd16, 8'd240, 8'd224, 8'd64, 8'd144, 8'd128, 8'd80, 8'd184,
  8'd40, 8'd232, 8'd200, 8'd112, 8'd248, 8'd24, 8'd112, 8'd176, 8'd128, 8'd128, 8'd56, 8'd40, 8'd152, 8'd24, 8'd184,
  8'd120, 8'd104, 8'd72, 8'd64, 8'd200, 8'd48, 8'd224, 8'd0, 8'd56, 8'd232, 8'd32, 8'd240, 8'd184, 8'd104, 8'd104, 8'd32, 8'd192,
  8'd200, 8'd200, 8'd64, 8'd152, 8'd72, 8'd216, 8'd216, 8'd80, 8'd0, 8'd80, 8'd0, 8'd0, 8'd160, 8'd120, 8'd40,
  8'd136, 8'd240, 8'd32, 8'd120, 8'd152, 8'd216, 8'd56, 8'd112, 8'd16, 8'd24, 8'd8, 8'd120, 8'd104, 8'd192, 8'd144, 8'd176, 8'd8,
  8'd16, 8'd96, 8'd104, 8'd168, 8'd80, 8'd192, 8'd232, 8'd112, 8'd112, 8'd56, 8'd88, 8'd176, 8'd240, 8'd32, 8'd176,
  8'd248, 8'd80, 8'd176, 8'd24, 8'd224, 8'd192, 8'd8, 8'd176, 8'd168, 8'd16, 8'd232, 8'd248, 8'd16, 8'd16, 8'd104, 8'd128,
  8'd232, 8'd0, 8'd32, 8'd240, 8'd112, 8'd32, 8'd184, 8'd184, 8'd56, 8'd232, 8'd80, 8'd144, 8'd16, 8'd72, 8'd240, 8'd208,
  8'd64, 8'd176, 8'd240, 8'd16, 8'd136, 8'd16, 8'd80, 8'd192, 8'd24, 8'd72, 8'd216, 8'd56, 8'd80, 8'd216, 8'd32, 8'd144, 8'd72,
  8'd24, 8'd64, 8'd248, 8'd0, 8'd224, 8'd72, 8'd32, 8'd136, 8'd232, 8'd240, 8'd72, 8'd32, 8'd88, 8'd128, 8'd104,
  8'd16, 8'd8, 8'd32, 8'd192, 8'd224, 8'd8, 8'd152, 8'd248, 8'd224, 8'd0, 8'd176, 8'd48, 8'd16, 8'd104, 8'd216, 8'd176, 8'd24,
  8'd240, 8'd200, 8'd80, 8'd248, 8'd208, 8'd128, 8'd200, 8'd72, 8'd8, 8'd152, 8'd128, 8'd80, 8'd120, 8'd80, 8'd152,
  8'd232, 8'd200, 8'd168, 8'd88, 8'd16, 8'd176, 8'd232, 8'd40, 8'd72, 8'd208, 8'd232, 8'd112, 8'd240, 8'd112, 8'd80, 8'd176,
  8'd176, 8'd16, 8'd72, 8'd120, 8'd32, 8'd184, 8'd224, 8'd80, 8'd24, 8'd176, 8'd0, 8'd208, 8'd16, 8'd56, 8'd112, 8'd16,
  8'd120, 8'd160, 8'd24, 8'd216, 8'd128, 8'd136, 8'd192, 8'd152, 8'd248, 8'd120, 8'd160, 8'd56, 8'd192, 8'd224, 8'd0, 8'd136,
  8'd112, 8'd112, 8'd8, 8'd8, 8'd184, 8'd168, 8'd88, 8'd160, 8'd120, 8'd160, 8'd240, 8'd168, 8'd32, 8'd40, 8'd168, 8'd88,
  8'd8, 8'd16, 8'd24, 8'd104, 8'd104, 8'd48, 8'd248, 8'd136, 8'd72, 8'd144, 8'd128, 8'd160, 8'd216, 8'd88, 8'd240, 8'd120,
  8'd232, 8'd72, 8'd192, 8'd200, 8'd248, 8'd192, 8'd48, 8'd240, 8'd104, 8'd208, 8'd40, 8'd104, 8'd16, 8'd128, 8'd80, 8'd224,
  8'd224, 8'd56, 8'd56, 8'd120, 8'd40, 8'd24, 8'd176, 8'd16, 8'd184, 8'd24, 8'd176, 8'd224, 8'd168, 8'd16, 8'd184, 8'd104,
  8'd136, 8'd200, 8'd168, 8'd208, 8'd120, 8'd200, 8'd224, 8'd40, 8'd208, 8'd16, 8'd112, 8'd160, 8'd192, 8'd224, 8'd64,
  8'd40,
  8'd232, 8'd120, 8'd24, 8'd232, 8'd168, 8'd80, 8'd88, 8'd144, 8'd104, 8'd72, 8'd192, 8'd112, 8'd0, 8'd112, 8'd104, 8'd224,
  8'd232, 8'd160, 8'd112, 8'd208, 8'd176, 8'd216, 8'd56, 8'd224, 8'd224, 8'd160, 8'd104, 8'd56, 8'd176, 8'd216, 8'd192,
  8'd24,
  8'd208, 8'd8, 8'd40, 8'd56, 8'd248, 8'd8, 8'd120, 8'd184, 8'd128, 8'd40, 8'd168, 8'd56, 8'd184, 8'd192, 8'd136, 8'd96, 8'd72,
  8'd216, 8'd8, 8'd64, 8'd72, 8'd56, 8'd16, 8'd176, 8'd144, 8'd16, 8'd128, 8'd176, 8'd136, 8'd208, 8'd120, 8'd16,
  8'd184, 8'd224, 8'd160, 8'd216, 8'd144, 8'd88, 8'd208, 8'd200, 8'd144, 8'd96, 8'd152, 8'd200, 8'd224, 8'd208, 8'd240,
  8'd120, 8'd8, 8'd104, 8'd184, 8'd112, 8'd168, 8'd200, 8'd112, 8'd72, 8'd0, 8'd192, 8'd0, 8'd40, 8'd120, 8'd136, 8'd112,
  8'd40,
  8'd152, 8'd56, 8'd144, 8'd32, 8'd224, 8'd240, 8'd32, 8'd192, 8'd56, 8'd200, 8'd16, 8'd136, 8'd104, 8'd192, 8'd192, 8'd0, 8'd0,
  8'd0, 8'd8, 8'd232, 8'd104, 8'd240, 8'd88, 8'd192, 8'd8, 8'd168, 8'd216, 8'd208, 8'd184, 8'd224, 8'd240, 8'd72,
  8'd152, 8'd72, 8'd168, 8'd184, 8'd176, 8'd216, 8'd48, 8'd144, 8'd80, 8'd32, 8'd184, 8'd208, 8'd112, 8'd160, 8'd88, 8'd88, 8'd8,
  8'd144, 8'd144, 8'd120, 8'd152, 8'd48, 8'd200, 8'd168, 8'd112, 8'd8, 8'd160, 8'd216, 8'd240, 8'd128, 8'd104, 8'd128,
  8'd144, 8'd248, 8'd64, 8'd168, 8'd136, 8'd240, 8'd160, 8'd56, 8'd136, 8'd216, 8'd80, 8'd56, 8'd192, 8'd32, 8'd64, 8'd128,
  8'd80, 8'd32, 8'd32, 8'd96, 8'd88, 8'd200, 8'd152, 8'd72, 8'd160, 8'd16, 8'd128, 8'd200, 8'd160, 8'd144, 8'd112, 8'd16,
  8'd112, 8'd152, 8'd56, 8'd136, 8'd56, 8'd216, 8'd8, 8'd24, 8'd192, 8'd144, 8'd176, 8'd200, 8'd48, 8'd72, 8'd40, 8'd72, 8'd240,
  8'd120, 8'd120, 8'd160, 8'd80, 8'd152, 8'd144, 8'd216, 8'd224, 8'd152, 8'd40, 8'd144, 8'd160, 8'd88, 8'd184, 8'd184,
  8'd192, 8'd128, 8'd0, 8'd200, 8'd72, 8'd112, 8'd208, 8'd248, 8'd152, 8'd0, 8'd152, 8'd8, 8'd40, 8'd16, 8'd168, 8'd152, 8'd64,
  8'd176, 8'd88, 8'd24, 8'd232, 8'd136, 8'd32, 8'd152, 8'd232, 8'd208, 8'd192, 8'd240, 8'd136, 8'd0, 8'd232, 8'd200,
  8'd8, 8'd216, 8'd104, 8'd184, 8'd64, 8'd192, 8'd8, 8'd96, 8'd184, 8'd120, 8'd208, 8'd80, 8'd16, 8'd64, 8'd136, 8'd136, 8'd72,
  8'd8, 8'd112, 8'd184, 8'd248, 8'd120, 8'd136, 8'd8, 8'd56, 8'd232, 8'd208, 8'd96, 8'd16, 8'd64, 8'd168, 8'd112,
  8'd48, 8'd32, 8'd184, 8'd224, 8'd72, 8'd88, 8'd128, 8'd184, 8'd72, 8'd168, 8'd224, 8'd216, 8'd160, 8'd232, 8'd64, 8'd168,
  8'd48, 8'd152, 8'd64, 8'd152, 8'd16, 8'd200, 8'd168, 8'd56, 8'd144, 8'd192, 8'd64, 8'd120, 8'd168, 8'd8, 8'd128, 8'd216,
  8'd16, 8'd8, 8'd104, 8'd32, 8'd128, 8'd96, 8'd160, 8'd88, 8'd136, 8'd96, 8'd56, 8'd16, 8'd128, 8'd56, 8'd88, 8'd16, 8'd208,
  8'd200, 8'd24, 8'd96, 8'd240, 8'd32, 8'd232, 8'd192, 8'd104, 8'd168, 8'd40, 8'd0, 8'd192, 8'd40, 8'd200, 8'd96,
  8'd184, 8'd8, 8'd72, 8'd216, 8'd104, 8'd232, 8'd112, 8'd248, 8'd8, 8'd8, 8'd248, 8'd192, 8'd152, 8'd32, 8'd0, 8'd168, 8'd232,
  8'd80, 8'd248, 8'd64, 8'd8, 8'd24, 8'd80, 8'd32, 8'd96, 8'd240, 8'd232, 8'd48, 8'd80, 8'd16, 8'd144, 8'd200,
  8'd16, 8'd48, 8'd88, 8'd40, 8'd112, 8'd232, 8'd88, 8'd168, 8'd56, 8'd160, 8'd232, 8'd16, 8'd128, 8'd248, 8'd48, 8'd80, 8'd200,
  8'd168, 8'd152, 8'd72, 8'd216, 8'd224, 8'd72, 8'd208, 8'd152, 8'd192, 8'd0, 8'd224, 8'd48, 8'd136, 8'd168, 8'd96,
  8'd16, 8'd152, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd224, 8'd227, 8'd227, 8'd227,
  8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0
};


  reg rst;
  reg [31:0] N;
  reg in_valid;
  wire in_bfr;
  reg [31:0] out_ld_bfr;
  reg [31:0] out_incnt;
  reg done;

  
endmodule; // test_flush_buf


test_flush_buf tfb(clock.val);
